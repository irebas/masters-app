<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Piotr Bujak" version="11.69132">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Lublin" name="2021 Główne Mistrzostwa Województwa Lubelskiego" course="LCM" deadline="2021-06-15" organizer="LOZP" reservecount="2" result.url="http://www.megatiming.pl/pkregowe" startmethod="1" timing="AUTOMATIC" nation="POL">
      <AGEDATE value="2021-06-19" type="YEAR" />
      <POOL name="Aqua Lublin" lanemax="9" />
      <FACILITY city="Lublin" name="Aqua Lublin" nation="POL" />
      <POINTTABLE pointtableid="3014" name="FINA Point Scoring" version="2021" />
      <CONTACT email="pioswim@wp.pl" name="Piotr Bujak" phone="510089179" />
      <QUALIFY from="2020-03-12" until="2021-06-17" />
      <SESSIONS>
        <SESSION date="2021-06-18" daytime="15:30" endtime="19:21" name="I BLOK" number="1" warmupfrom="15:00" warmupuntil="15:25">
          <EVENTS>
            <EVENT eventid="1059" daytime="15:30" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1061" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16909" />
                    <RANKING order="2" place="2" resultid="16915" />
                    <RANKING order="3" place="3" resultid="17090" />
                    <RANKING order="4" place="4" resultid="18483" />
                    <RANKING order="5" place="5" resultid="18400" />
                    <RANKING order="6" place="6" resultid="18141" />
                    <RANKING order="7" place="7" resultid="17607" />
                    <RANKING order="8" place="8" resultid="17096" />
                    <RANKING order="9" place="9" resultid="17601" />
                    <RANKING order="10" place="10" resultid="17324" />
                    <RANKING order="11" place="11" resultid="18620" />
                    <RANKING order="12" place="12" resultid="17318" />
                    <RANKING order="13" place="13" resultid="18348" />
                    <RANKING order="14" place="14" resultid="17158" />
                    <RANKING order="15" place="15" resultid="18101" />
                    <RANKING order="16" place="16" resultid="18144" />
                    <RANKING order="17" place="17" resultid="18341" />
                    <RANKING order="18" place="18" resultid="17613" />
                    <RANKING order="19" place="19" resultid="18108" />
                    <RANKING order="20" place="20" resultid="17930" />
                    <RANKING order="21" place="21" resultid="17976" />
                    <RANKING order="22" place="22" resultid="18128" />
                    <RANKING order="23" place="23" resultid="18584" />
                    <RANKING order="24" place="24" resultid="18587" />
                    <RANKING order="25" place="-1" resultid="18200" />
                    <RANKING order="26" place="-1" resultid="18476" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1062" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18057" />
                    <RANKING order="2" place="2" resultid="17083" />
                    <RANKING order="3" place="3" resultid="17766" />
                    <RANKING order="4" place="4" resultid="18051" />
                    <RANKING order="5" place="5" resultid="16921" />
                    <RANKING order="6" place="5" resultid="17587" />
                    <RANKING order="7" place="7" resultid="18545" />
                    <RANKING order="8" place="8" resultid="18366" />
                    <RANKING order="9" place="9" resultid="18395" />
                    <RANKING order="10" place="10" resultid="17593" />
                    <RANKING order="11" place="11" resultid="18121" />
                    <RANKING order="12" place="12" resultid="17979" />
                    <RANKING order="13" place="-1" resultid="17596" />
                    <RANKING order="14" place="-1" resultid="17923" />
                    <RANKING order="15" place="-1" resultid="18391" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1060" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17257" />
                    <RANKING order="2" place="2" resultid="18057" />
                    <RANKING order="3" place="3" resultid="17302" />
                    <RANKING order="4" place="4" resultid="18193" />
                    <RANKING order="5" place="5" resultid="18207" />
                    <RANKING order="6" place="6" resultid="17264" />
                    <RANKING order="7" place="7" resultid="18215" />
                    <RANKING order="8" place="8" resultid="17270" />
                    <RANKING order="9" place="9" resultid="17283" />
                    <RANKING order="10" place="10" resultid="17290" />
                    <RANKING order="11" place="11" resultid="17083" />
                    <RANKING order="12" place="12" resultid="17309" />
                    <RANKING order="13" place="13" resultid="16909" />
                    <RANKING order="14" place="14" resultid="17315" />
                    <RANKING order="15" place="15" resultid="16915" />
                    <RANKING order="16" place="16" resultid="17296" />
                    <RANKING order="17" place="17" resultid="17766" />
                    <RANKING order="18" place="18" resultid="17165" />
                    <RANKING order="19" place="19" resultid="17277" />
                    <RANKING order="20" place="20" resultid="16930" />
                    <RANKING order="21" place="21" resultid="18051" />
                    <RANKING order="22" place="22" resultid="16921" />
                    <RANKING order="23" place="22" resultid="17587" />
                    <RANKING order="24" place="24" resultid="17090" />
                    <RANKING order="25" place="25" resultid="18545" />
                    <RANKING order="26" place="26" resultid="18483" />
                    <RANKING order="27" place="27" resultid="16925" />
                    <RANKING order="28" place="28" resultid="18400" />
                    <RANKING order="29" place="29" resultid="17078" />
                    <RANKING order="30" place="30" resultid="18141" />
                    <RANKING order="31" place="31" resultid="18366" />
                    <RANKING order="32" place="32" resultid="17607" />
                    <RANKING order="33" place="33" resultid="17096" />
                    <RANKING order="34" place="34" resultid="17601" />
                    <RANKING order="35" place="35" resultid="17324" />
                    <RANKING order="36" place="36" resultid="18395" />
                    <RANKING order="37" place="37" resultid="17171" />
                    <RANKING order="38" place="38" resultid="18620" />
                    <RANKING order="39" place="39" resultid="17318" />
                    <RANKING order="40" place="40" resultid="18590" />
                    <RANKING order="41" place="41" resultid="18348" />
                    <RANKING order="42" place="42" resultid="18115" />
                    <RANKING order="43" place="43" resultid="17593" />
                    <RANKING order="44" place="44" resultid="17158" />
                    <RANKING order="45" place="45" resultid="18101" />
                    <RANKING order="46" place="46" resultid="17584" />
                    <RANKING order="47" place="47" resultid="18121" />
                    <RANKING order="48" place="48" resultid="18144" />
                    <RANKING order="49" place="49" resultid="18341" />
                    <RANKING order="50" place="50" resultid="17613" />
                    <RANKING order="51" place="51" resultid="18108" />
                    <RANKING order="52" place="52" resultid="17930" />
                    <RANKING order="53" place="53" resultid="17976" />
                    <RANKING order="54" place="54" resultid="18128" />
                    <RANKING order="55" place="55" resultid="18584" />
                    <RANKING order="56" place="56" resultid="18587" />
                    <RANKING order="57" place="57" resultid="17979" />
                    <RANKING order="58" place="-1" resultid="17596" />
                    <RANKING order="59" place="-1" resultid="17923" />
                    <RANKING order="60" place="-1" resultid="18200" />
                    <RANKING order="61" place="-1" resultid="18391" />
                    <RANKING order="62" place="-1" resultid="18476" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="18945" daytime="15:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="18946" daytime="15:31" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="18947" daytime="15:33" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="18948" daytime="15:34" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="18949" daytime="15:35" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="18950" daytime="15:37" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="18951" daytime="15:38" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1063" daytime="15:39" gender="M" number="2" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1064" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18222" />
                    <RANKING order="2" place="2" resultid="17235" />
                    <RANKING order="3" place="3" resultid="18564" />
                    <RANKING order="4" place="4" resultid="18150" />
                    <RANKING order="5" place="5" resultid="18147" />
                    <RANKING order="6" place="6" resultid="18153" />
                    <RANKING order="7" place="7" resultid="16959" />
                    <RANKING order="8" place="8" resultid="18605" />
                    <RANKING order="9" place="9" resultid="17355" />
                    <RANKING order="10" place="10" resultid="17801" />
                    <RANKING order="11" place="11" resultid="17202" />
                    <RANKING order="12" place="12" resultid="18162" />
                    <RANKING order="13" place="13" resultid="17242" />
                    <RANKING order="14" place="14" resultid="17794" />
                    <RANKING order="15" place="15" resultid="17361" />
                    <RANKING order="16" place="16" resultid="18159" />
                    <RANKING order="17" place="17" resultid="17374" />
                    <RANKING order="18" place="18" resultid="17177" />
                    <RANKING order="19" place="19" resultid="18498" />
                    <RANKING order="20" place="20" resultid="17102" />
                    <RANKING order="21" place="21" resultid="17660" />
                    <RANKING order="22" place="22" resultid="17998" />
                    <RANKING order="23" place="23" resultid="18489" />
                    <RANKING order="24" place="24" resultid="17667" />
                    <RANKING order="25" place="25" resultid="17368" />
                    <RANKING order="26" place="26" resultid="16964" />
                    <RANKING order="27" place="27" resultid="17808" />
                    <RANKING order="28" place="28" resultid="16945" />
                    <RANKING order="29" place="29" resultid="18494" />
                    <RANKING order="30" place="30" resultid="18595" />
                    <RANKING order="31" place="31" resultid="18269" />
                    <RANKING order="32" place="32" resultid="17656" />
                    <RANKING order="33" place="33" resultid="17512" />
                    <RANKING order="34" place="34" resultid="17348" />
                    <RANKING order="35" place="35" resultid="17815" />
                    <RANKING order="36" place="36" resultid="18290" />
                    <RANKING order="37" place="37" resultid="18251" />
                    <RANKING order="38" place="38" resultid="18602" />
                    <RANKING order="39" place="39" resultid="18237" />
                    <RANKING order="40" place="40" resultid="17648" />
                    <RANKING order="41" place="41" resultid="18011" />
                    <RANKING order="42" place="42" resultid="18283" />
                    <RANKING order="43" place="43" resultid="18516" />
                    <RANKING order="44" place="44" resultid="18276" />
                    <RANKING order="45" place="45" resultid="17993" />
                    <RANKING order="46" place="-1" resultid="17554" />
                    <RANKING order="47" place="-1" resultid="18511" />
                    <RANKING order="48" place="-1" resultid="17505" />
                    <RANKING order="49" place="-1" resultid="17988" />
                    <RANKING order="50" place="-1" resultid="18156" />
                    <RANKING order="51" place="-1" resultid="18165" />
                    <RANKING order="52" place="-1" resultid="18244" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17641" />
                    <RANKING order="2" place="2" resultid="17184" />
                    <RANKING order="3" place="3" resultid="17228" />
                    <RANKING order="4" place="4" resultid="18262" />
                    <RANKING order="5" place="5" resultid="16976" />
                    <RANKING order="6" place="6" resultid="17215" />
                    <RANKING order="7" place="7" resultid="17249" />
                    <RANKING order="8" place="8" resultid="16955" />
                    <RANKING order="9" place="9" resultid="17634" />
                    <RANKING order="10" place="10" resultid="18353" />
                    <RANKING order="11" place="11" resultid="17548" />
                    <RANKING order="12" place="12" resultid="16950" />
                    <RANKING order="13" place="13" resultid="18549" />
                    <RANKING order="14" place="14" resultid="17681" />
                    <RANKING order="15" place="15" resultid="18230" />
                    <RANKING order="16" place="16" resultid="17787" />
                    <RANKING order="17" place="17" resultid="18016" />
                    <RANKING order="18" place="18" resultid="17559" />
                    <RANKING order="19" place="19" resultid="17630" />
                    <RANKING order="20" place="20" resultid="18005" />
                    <RANKING order="21" place="21" resultid="17982" />
                    <RANKING order="22" place="22" resultid="18409" />
                    <RANKING order="23" place="23" resultid="18504" />
                    <RANKING order="24" place="24" resultid="18554" />
                    <RANKING order="25" place="25" resultid="18559" />
                    <RANKING order="26" place="26" resultid="18168" />
                    <RANKING order="27" place="27" resultid="18419" />
                    <RANKING order="28" place="28" resultid="18415" />
                    <RANKING order="29" place="29" resultid="17196" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17222" />
                    <RANKING order="2" place="2" resultid="17336" />
                    <RANKING order="3" place="3" resultid="17342" />
                    <RANKING order="4" place="4" resultid="17380" />
                    <RANKING order="5" place="5" resultid="17545" />
                    <RANKING order="6" place="6" resultid="17208" />
                    <RANKING order="7" place="7" resultid="17386" />
                    <RANKING order="8" place="8" resultid="17641" />
                    <RANKING order="9" place="9" resultid="17184" />
                    <RANKING order="10" place="10" resultid="18258" />
                    <RANKING order="11" place="11" resultid="16982" />
                    <RANKING order="12" place="12" resultid="17189" />
                    <RANKING order="13" place="13" resultid="17539" />
                    <RANKING order="14" place="14" resultid="17228" />
                    <RANKING order="15" place="15" resultid="18262" />
                    <RANKING order="16" place="16" resultid="16969" />
                    <RANKING order="17" place="17" resultid="16976" />
                    <RANKING order="18" place="18" resultid="18133" />
                    <RANKING order="19" place="19" resultid="17399" />
                    <RANKING order="20" place="20" resultid="17215" />
                    <RANKING order="21" place="21" resultid="18222" />
                    <RANKING order="22" place="22" resultid="17249" />
                    <RANKING order="23" place="23" resultid="16955" />
                    <RANKING order="24" place="24" resultid="17235" />
                    <RANKING order="25" place="25" resultid="17634" />
                    <RANKING order="26" place="26" resultid="17620" />
                    <RANKING order="27" place="27" resultid="17533" />
                    <RANKING order="28" place="28" resultid="18564" />
                    <RANKING order="29" place="29" resultid="18353" />
                    <RANKING order="30" place="30" resultid="18150" />
                    <RANKING order="31" place="31" resultid="17548" />
                    <RANKING order="32" place="32" resultid="16950" />
                    <RANKING order="33" place="33" resultid="18549" />
                    <RANKING order="34" place="34" resultid="17681" />
                    <RANKING order="35" place="35" resultid="18147" />
                    <RANKING order="36" place="36" resultid="17650" />
                    <RANKING order="37" place="37" resultid="18230" />
                    <RANKING order="38" place="38" resultid="17787" />
                    <RANKING order="39" place="39" resultid="18016" />
                    <RANKING order="40" place="40" resultid="17559" />
                    <RANKING order="41" place="41" resultid="17527" />
                    <RANKING order="42" place="42" resultid="17630" />
                    <RANKING order="43" place="43" resultid="18153" />
                    <RANKING order="44" place="44" resultid="18005" />
                    <RANKING order="45" place="45" resultid="16959" />
                    <RANKING order="46" place="46" resultid="18605" />
                    <RANKING order="47" place="47" resultid="17355" />
                    <RANKING order="48" place="48" resultid="17801" />
                    <RANKING order="49" place="49" resultid="17202" />
                    <RANKING order="50" place="50" resultid="17982" />
                    <RANKING order="51" place="51" resultid="18162" />
                    <RANKING order="52" place="52" resultid="18409" />
                    <RANKING order="53" place="53" resultid="17242" />
                    <RANKING order="54" place="54" resultid="18504" />
                    <RANKING order="55" place="55" resultid="17794" />
                    <RANKING order="56" place="56" resultid="17361" />
                    <RANKING order="57" place="57" resultid="18554" />
                    <RANKING order="58" place="58" resultid="18559" />
                    <RANKING order="59" place="59" resultid="18159" />
                    <RANKING order="60" place="60" resultid="17374" />
                    <RANKING order="61" place="61" resultid="17177" />
                    <RANKING order="62" place="62" resultid="17625" />
                    <RANKING order="63" place="63" resultid="18498" />
                    <RANKING order="64" place="64" resultid="18168" />
                    <RANKING order="65" place="65" resultid="17102" />
                    <RANKING order="66" place="66" resultid="17660" />
                    <RANKING order="67" place="67" resultid="18419" />
                    <RANKING order="68" place="68" resultid="17998" />
                    <RANKING order="69" place="69" resultid="18489" />
                    <RANKING order="70" place="70" resultid="17667" />
                    <RANKING order="71" place="71" resultid="17368" />
                    <RANKING order="72" place="72" resultid="16964" />
                    <RANKING order="73" place="73" resultid="18415" />
                    <RANKING order="74" place="74" resultid="17808" />
                    <RANKING order="75" place="75" resultid="16945" />
                    <RANKING order="76" place="76" resultid="18494" />
                    <RANKING order="77" place="77" resultid="17196" />
                    <RANKING order="78" place="78" resultid="18595" />
                    <RANKING order="79" place="79" resultid="18269" />
                    <RANKING order="80" place="80" resultid="17656" />
                    <RANKING order="81" place="81" resultid="17512" />
                    <RANKING order="82" place="82" resultid="17348" />
                    <RANKING order="83" place="83" resultid="17815" />
                    <RANKING order="84" place="84" resultid="18290" />
                    <RANKING order="85" place="85" resultid="18251" />
                    <RANKING order="86" place="86" resultid="18602" />
                    <RANKING order="87" place="87" resultid="18237" />
                    <RANKING order="88" place="88" resultid="17648" />
                    <RANKING order="89" place="89" resultid="18011" />
                    <RANKING order="90" place="90" resultid="18283" />
                    <RANKING order="91" place="91" resultid="18516" />
                    <RANKING order="92" place="92" resultid="18276" />
                    <RANKING order="93" place="93" resultid="17993" />
                    <RANKING order="94" place="-1" resultid="17554" />
                    <RANKING order="95" place="-1" resultid="18511" />
                    <RANKING order="96" place="-1" resultid="17505" />
                    <RANKING order="97" place="-1" resultid="17988" />
                    <RANKING order="98" place="-1" resultid="18156" />
                    <RANKING order="99" place="-1" resultid="18165" />
                    <RANKING order="100" place="-1" resultid="18244" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="18952" daytime="15:39" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="18953" daytime="15:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="18954" daytime="15:42" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="18955" daytime="15:43" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="18956" daytime="15:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="18957" daytime="15:46" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="18958" daytime="15:47" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="18959" daytime="15:48" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="18960" daytime="15:49" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="18961" daytime="15:51" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="18962" daytime="15:52" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1067" daytime="15:53" gender="F" number="3" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1068" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16990" />
                    <RANKING order="2" place="2" resultid="17688" />
                    <RANKING order="3" place="3" resultid="17709" />
                    <RANKING order="4" place="4" resultid="16995" />
                    <RANKING order="5" place="5" resultid="17319" />
                    <RANKING order="6" place="6" resultid="17608" />
                    <RANKING order="7" place="7" resultid="17716" />
                    <RANKING order="8" place="8" resultid="17159" />
                    <RANKING order="9" place="9" resultid="18102" />
                    <RANKING order="10" place="10" resultid="17931" />
                    <RANKING order="11" place="11" resultid="18145" />
                    <RANKING order="12" place="12" resultid="18349" />
                    <RANKING order="13" place="13" resultid="17944" />
                    <RANKING order="14" place="14" resultid="18588" />
                    <RANKING order="15" place="15" resultid="17614" />
                    <RANKING order="16" place="16" resultid="18585" />
                    <RANKING order="17" place="17" resultid="18129" />
                    <RANKING order="18" place="18" resultid="17977" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17109" />
                    <RANKING order="2" place="2" resultid="18058" />
                    <RANKING order="3" place="3" resultid="18566" />
                    <RANKING order="4" place="4" resultid="17702" />
                    <RANKING order="5" place="5" resultid="17822" />
                    <RANKING order="6" place="6" resultid="17123" />
                    <RANKING order="7" place="7" resultid="17695" />
                    <RANKING order="8" place="8" resultid="18297" />
                    <RANKING order="9" place="9" resultid="17002" />
                    <RANKING order="10" place="10" resultid="17588" />
                    <RANKING order="11" place="11" resultid="18304" />
                    <RANKING order="12" place="12" resultid="18122" />
                    <RANKING order="13" place="13" resultid="17597" />
                    <RANKING order="14" place="14" resultid="17980" />
                    <RANKING order="15" place="-1" resultid="17924" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17404" />
                    <RANKING order="2" place="2" resultid="17258" />
                    <RANKING order="3" place="3" resultid="17109" />
                    <RANKING order="4" place="4" resultid="18058" />
                    <RANKING order="5" place="5" resultid="17408" />
                    <RANKING order="6" place="6" resultid="17116" />
                    <RANKING order="7" place="7" resultid="18566" />
                    <RANKING order="8" place="8" resultid="17702" />
                    <RANKING order="9" place="9" resultid="17822" />
                    <RANKING order="10" place="10" resultid="16990" />
                    <RANKING order="11" place="10" resultid="17123" />
                    <RANKING order="12" place="12" resultid="17695" />
                    <RANKING order="13" place="13" resultid="18297" />
                    <RANKING order="14" place="14" resultid="17002" />
                    <RANKING order="15" place="15" resultid="17588" />
                    <RANKING order="16" place="16" resultid="18063" />
                    <RANKING order="17" place="17" resultid="17688" />
                    <RANKING order="18" place="18" resultid="17709" />
                    <RANKING order="19" place="19" resultid="16995" />
                    <RANKING order="20" place="20" resultid="17319" />
                    <RANKING order="21" place="21" resultid="18304" />
                    <RANKING order="22" place="22" resultid="17608" />
                    <RANKING order="23" place="23" resultid="17716" />
                    <RANKING order="24" place="24" resultid="18122" />
                    <RANKING order="25" place="25" resultid="17159" />
                    <RANKING order="26" place="26" resultid="18102" />
                    <RANKING order="27" place="27" resultid="18591" />
                    <RANKING order="28" place="28" resultid="17931" />
                    <RANKING order="29" place="29" resultid="18145" />
                    <RANKING order="30" place="30" resultid="18116" />
                    <RANKING order="31" place="31" resultid="18349" />
                    <RANKING order="32" place="32" resultid="17597" />
                    <RANKING order="33" place="33" resultid="17944" />
                    <RANKING order="34" place="34" resultid="18588" />
                    <RANKING order="35" place="35" resultid="17980" />
                    <RANKING order="36" place="36" resultid="17614" />
                    <RANKING order="37" place="37" resultid="18585" />
                    <RANKING order="38" place="38" resultid="18129" />
                    <RANKING order="39" place="39" resultid="17977" />
                    <RANKING order="40" place="-1" resultid="17924" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="18963" daytime="15:53" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="18964" daytime="15:54" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="18965" daytime="15:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="18966" daytime="15:58" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="18967" daytime="15:59" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1071" daytime="16:00" gender="M" number="4" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1072" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18148" />
                    <RANKING order="2" place="2" resultid="18175" />
                    <RANKING order="3" place="3" resultid="17130" />
                    <RANKING order="4" place="4" resultid="17843" />
                    <RANKING order="5" place="5" resultid="17722" />
                    <RANKING order="6" place="6" resultid="17950" />
                    <RANKING order="7" place="7" resultid="17414" />
                    <RANKING order="8" place="8" resultid="17375" />
                    <RANKING order="9" place="9" resultid="17795" />
                    <RANKING order="10" place="10" resultid="17203" />
                    <RANKING order="11" place="11" resultid="18614" />
                    <RANKING order="12" place="12" resultid="17519" />
                    <RANKING order="13" place="13" resultid="17243" />
                    <RANKING order="14" place="14" resultid="18318" />
                    <RANKING order="15" place="15" resultid="18610" />
                    <RANKING order="16" place="16" resultid="18163" />
                    <RANKING order="17" place="17" resultid="17362" />
                    <RANKING order="18" place="18" resultid="18372" />
                    <RANKING order="19" place="19" resultid="17136" />
                    <RANKING order="20" place="20" resultid="16965" />
                    <RANKING order="21" place="21" resultid="17007" />
                    <RANKING order="22" place="22" resultid="17999" />
                    <RANKING order="23" place="23" resultid="17816" />
                    <RANKING order="24" place="24" resultid="18532" />
                    <RANKING order="25" place="25" resultid="17349" />
                    <RANKING order="26" place="26" resultid="18596" />
                    <RANKING order="27" place="27" resultid="18277" />
                    <RANKING order="28" place="28" resultid="17513" />
                    <RANKING order="29" place="29" resultid="18603" />
                    <RANKING order="30" place="30" resultid="18012" />
                    <RANKING order="31" place="31" resultid="17994" />
                    <RANKING order="32" place="32" resultid="18284" />
                    <RANKING order="33" place="-1" resultid="18154" />
                    <RANKING order="34" place="-1" resultid="18527" />
                    <RANKING order="35" place="-1" resultid="17989" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1073" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17836" />
                    <RANKING order="2" place="2" resultid="17642" />
                    <RANKING order="3" place="3" resultid="16977" />
                    <RANKING order="4" place="4" resultid="18069" />
                    <RANKING order="5" place="5" resultid="17829" />
                    <RANKING order="6" place="6" resultid="18311" />
                    <RANKING order="7" place="7" resultid="17788" />
                    <RANKING order="8" place="8" resultid="18505" />
                    <RANKING order="9" place="9" resultid="17568" />
                    <RANKING order="10" place="10" resultid="16951" />
                    <RANKING order="11" place="11" resultid="17017" />
                    <RANKING order="12" place="12" resultid="18354" />
                    <RANKING order="13" place="13" resultid="18410" />
                    <RANKING order="14" place="14" resultid="18006" />
                    <RANKING order="15" place="15" resultid="18560" />
                    <RANKING order="16" place="-1" resultid="17631" />
                    <RANKING order="17" place="-1" resultid="17983" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1074" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17427" />
                    <RANKING order="2" place="2" resultid="17431" />
                    <RANKING order="3" place="3" resultid="17564" />
                    <RANKING order="4" place="4" resultid="17021" />
                    <RANKING order="5" place="5" resultid="17012" />
                    <RANKING order="6" place="6" resultid="17420" />
                    <RANKING order="7" place="7" resultid="17836" />
                    <RANKING order="8" place="8" resultid="17642" />
                    <RANKING order="9" place="9" resultid="18134" />
                    <RANKING order="10" place="10" resultid="16977" />
                    <RANKING order="11" place="11" resultid="18069" />
                    <RANKING order="12" place="12" resultid="17829" />
                    <RANKING order="13" place="13" resultid="18148" />
                    <RANKING order="14" place="14" resultid="18175" />
                    <RANKING order="15" place="15" resultid="17130" />
                    <RANKING order="16" place="16" resultid="18311" />
                    <RANKING order="17" place="17" resultid="17788" />
                    <RANKING order="18" place="18" resultid="18505" />
                    <RANKING order="19" place="19" resultid="17568" />
                    <RANKING order="20" place="20" resultid="16951" />
                    <RANKING order="21" place="21" resultid="17017" />
                    <RANKING order="22" place="22" resultid="17843" />
                    <RANKING order="23" place="23" resultid="18354" />
                    <RANKING order="24" place="24" resultid="18410" />
                    <RANKING order="25" place="25" resultid="17722" />
                    <RANKING order="26" place="26" resultid="18006" />
                    <RANKING order="27" place="27" resultid="17950" />
                    <RANKING order="28" place="28" resultid="17414" />
                    <RANKING order="29" place="29" resultid="17375" />
                    <RANKING order="30" place="30" resultid="17795" />
                    <RANKING order="31" place="31" resultid="17203" />
                    <RANKING order="32" place="32" resultid="18614" />
                    <RANKING order="33" place="33" resultid="17519" />
                    <RANKING order="34" place="34" resultid="18560" />
                    <RANKING order="35" place="35" resultid="17243" />
                    <RANKING order="36" place="36" resultid="17626" />
                    <RANKING order="37" place="37" resultid="18318" />
                    <RANKING order="38" place="38" resultid="18610" />
                    <RANKING order="39" place="39" resultid="18163" />
                    <RANKING order="40" place="40" resultid="17362" />
                    <RANKING order="41" place="41" resultid="18372" />
                    <RANKING order="42" place="42" resultid="17136" />
                    <RANKING order="43" place="43" resultid="16965" />
                    <RANKING order="44" place="44" resultid="17007" />
                    <RANKING order="45" place="45" resultid="17999" />
                    <RANKING order="46" place="46" resultid="17816" />
                    <RANKING order="47" place="47" resultid="18532" />
                    <RANKING order="48" place="48" resultid="17349" />
                    <RANKING order="49" place="49" resultid="18596" />
                    <RANKING order="50" place="50" resultid="18277" />
                    <RANKING order="51" place="51" resultid="17513" />
                    <RANKING order="52" place="52" resultid="18603" />
                    <RANKING order="53" place="53" resultid="18012" />
                    <RANKING order="54" place="54" resultid="17994" />
                    <RANKING order="55" place="55" resultid="18284" />
                    <RANKING order="56" place="-1" resultid="17631" />
                    <RANKING order="57" place="-1" resultid="17651" />
                    <RANKING order="58" place="-1" resultid="18154" />
                    <RANKING order="59" place="-1" resultid="18527" />
                    <RANKING order="60" place="-1" resultid="17983" />
                    <RANKING order="61" place="-1" resultid="17989" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="18968" daytime="16:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="18969" daytime="16:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="18970" daytime="16:03" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="18971" daytime="16:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="18972" daytime="16:06" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="18973" daytime="16:08" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="18974" daytime="16:09" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1075" daytime="16:16" gender="F" number="5" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1076" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18178" />
                    <RANKING order="2" place="2" resultid="16996" />
                    <RANKING order="3" place="3" resultid="17142" />
                    <RANKING order="4" place="4" resultid="17729" />
                    <RANKING order="5" place="5" resultid="18023" />
                    <RANKING order="6" place="6" resultid="18109" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1077" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17026" />
                    <RANKING order="2" place="2" resultid="18325" />
                    <RANKING order="3" place="3" resultid="17084" />
                    <RANKING order="4" place="4" resultid="17823" />
                    <RANKING order="5" place="5" resultid="18075" />
                    <RANKING order="6" place="6" resultid="18537" />
                    <RANKING order="7" place="7" resultid="17043" />
                    <RANKING order="8" place="8" resultid="17957" />
                    <RANKING order="9" place="9" resultid="17032" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1078" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17405" />
                    <RANKING order="2" place="2" resultid="17444" />
                    <RANKING order="3" place="3" resultid="17437" />
                    <RANKING order="4" place="4" resultid="17457" />
                    <RANKING order="5" place="5" resultid="17291" />
                    <RANKING order="6" place="6" resultid="17451" />
                    <RANKING order="7" place="7" resultid="17026" />
                    <RANKING order="8" place="8" resultid="18178" />
                    <RANKING order="9" place="9" resultid="18325" />
                    <RANKING order="10" place="10" resultid="17084" />
                    <RANKING order="11" place="11" resultid="17823" />
                    <RANKING order="12" place="12" resultid="18075" />
                    <RANKING order="13" place="13" resultid="17037" />
                    <RANKING order="14" place="14" resultid="18537" />
                    <RANKING order="15" place="15" resultid="18064" />
                    <RANKING order="16" place="16" resultid="17043" />
                    <RANKING order="17" place="17" resultid="17957" />
                    <RANKING order="18" place="18" resultid="17166" />
                    <RANKING order="19" place="19" resultid="16996" />
                    <RANKING order="20" place="20" resultid="17142" />
                    <RANKING order="21" place="21" resultid="17032" />
                    <RANKING order="22" place="22" resultid="17729" />
                    <RANKING order="23" place="23" resultid="18023" />
                    <RANKING order="24" place="24" resultid="18109" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="18975" daytime="16:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="18976" daytime="16:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="18977" daytime="16:20" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1079" daytime="16:22" gender="M" number="6" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1080" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17149" />
                    <RANKING order="2" place="2" resultid="17802" />
                    <RANKING order="3" place="3" resultid="18030" />
                    <RANKING order="4" place="4" resultid="18606" />
                    <RANKING order="5" place="5" resultid="17103" />
                    <RANKING order="6" place="6" resultid="18291" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1081" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18081" />
                    <RANKING order="2" place="2" resultid="17837" />
                    <RANKING order="3" place="3" resultid="17229" />
                    <RANKING order="4" place="4" resultid="17572" />
                    <RANKING order="5" place="5" resultid="17736" />
                    <RANKING order="6" place="6" resultid="17049" />
                    <RANKING order="7" place="7" resultid="17851" />
                    <RANKING order="8" place="8" resultid="18263" />
                    <RANKING order="9" place="9" resultid="17858" />
                    <RANKING order="10" place="10" resultid="18416" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1082" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17337" />
                    <RANKING order="2" place="2" resultid="17472" />
                    <RANKING order="3" place="3" resultid="17478" />
                    <RANKING order="4" place="4" resultid="17464" />
                    <RANKING order="5" place="5" resultid="16983" />
                    <RANKING order="6" place="6" resultid="18081" />
                    <RANKING order="7" place="7" resultid="17468" />
                    <RANKING order="8" place="8" resultid="17837" />
                    <RANKING order="9" place="9" resultid="17229" />
                    <RANKING order="10" place="10" resultid="17209" />
                    <RANKING order="11" place="11" resultid="17572" />
                    <RANKING order="12" place="12" resultid="17736" />
                    <RANKING order="13" place="13" resultid="17387" />
                    <RANKING order="14" place="14" resultid="17049" />
                    <RANKING order="15" place="15" resultid="17851" />
                    <RANKING order="16" place="16" resultid="18360" />
                    <RANKING order="17" place="17" resultid="18263" />
                    <RANKING order="18" place="18" resultid="17540" />
                    <RANKING order="19" place="19" resultid="17858" />
                    <RANKING order="20" place="20" resultid="17149" />
                    <RANKING order="21" place="21" resultid="17802" />
                    <RANKING order="22" place="22" resultid="18030" />
                    <RANKING order="23" place="23" resultid="18606" />
                    <RANKING order="24" place="24" resultid="18416" />
                    <RANKING order="25" place="25" resultid="17103" />
                    <RANKING order="26" place="26" resultid="18291" />
                    <RANKING order="27" place="-1" resultid="16841" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="18978" daytime="16:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="18979" daytime="16:24" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="18980" daytime="16:26" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="18981" daytime="16:28" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1083" daytime="16:36" gender="F" number="7" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1084" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16910" />
                    <RANKING order="2" place="2" resultid="18484" />
                    <RANKING order="3" place="3" resultid="16991" />
                    <RANKING order="4" place="4" resultid="16916" />
                    <RANKING order="5" place="5" resultid="18142" />
                    <RANKING order="6" place="6" resultid="18036" />
                    <RANKING order="7" place="7" resultid="17091" />
                    <RANKING order="8" place="8" resultid="17602" />
                    <RANKING order="9" place="9" resultid="17325" />
                    <RANKING order="10" place="10" resultid="17717" />
                    <RANKING order="11" place="-1" resultid="18201" />
                    <RANKING order="12" place="-1" resultid="18477" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1085" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17124" />
                    <RANKING order="2" place="2" resultid="17696" />
                    <RANKING order="3" place="3" resultid="18326" />
                    <RANKING order="4" place="4" resultid="17003" />
                    <RANKING order="5" place="5" resultid="18367" />
                    <RANKING order="6" place="6" resultid="18396" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1086" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17055" />
                    <RANKING order="2" place="2" resultid="18332" />
                    <RANKING order="3" place="3" resultid="18208" />
                    <RANKING order="4" place="4" resultid="17284" />
                    <RANKING order="5" place="5" resultid="17310" />
                    <RANKING order="6" place="6" resultid="17271" />
                    <RANKING order="7" place="7" resultid="17485" />
                    <RANKING order="8" place="8" resultid="17445" />
                    <RANKING order="9" place="9" resultid="18194" />
                    <RANKING order="10" place="10" resultid="17458" />
                    <RANKING order="11" place="11" resultid="17438" />
                    <RANKING order="12" place="12" resultid="17124" />
                    <RANKING order="13" place="13" resultid="17278" />
                    <RANKING order="14" place="14" resultid="17452" />
                    <RANKING order="15" place="15" resultid="17038" />
                    <RANKING order="16" place="16" resultid="17696" />
                    <RANKING order="17" place="17" resultid="16910" />
                    <RANKING order="18" place="18" resultid="17079" />
                    <RANKING order="19" place="19" resultid="16931" />
                    <RANKING order="20" place="20" resultid="17117" />
                    <RANKING order="21" place="21" resultid="18484" />
                    <RANKING order="22" place="22" resultid="16991" />
                    <RANKING order="23" place="23" resultid="16916" />
                    <RANKING order="24" place="24" resultid="18326" />
                    <RANKING order="25" place="25" resultid="18142" />
                    <RANKING order="26" place="26" resultid="18036" />
                    <RANKING order="27" place="27" resultid="17003" />
                    <RANKING order="28" place="28" resultid="17091" />
                    <RANKING order="29" place="29" resultid="18367" />
                    <RANKING order="30" place="30" resultid="18396" />
                    <RANKING order="31" place="31" resultid="17602" />
                    <RANKING order="32" place="32" resultid="17325" />
                    <RANKING order="33" place="33" resultid="17717" />
                    <RANKING order="34" place="34" resultid="17172" />
                    <RANKING order="35" place="-1" resultid="18201" />
                    <RANKING order="36" place="-1" resultid="18477" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="18982" daytime="16:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="18983" daytime="16:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="18984" daytime="16:43" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="18985" daytime="16:46" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1087" daytime="16:49" gender="M" number="8" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1088" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18223" />
                    <RANKING order="2" place="2" resultid="18151" />
                    <RANKING order="3" place="3" resultid="17236" />
                    <RANKING order="4" place="4" resultid="17415" />
                    <RANKING order="5" place="5" resultid="17879" />
                    <RANKING order="6" place="6" resultid="17555" />
                    <RANKING order="7" place="7" resultid="16960" />
                    <RANKING order="8" place="8" resultid="17506" />
                    <RANKING order="9" place="9" resultid="18031" />
                    <RANKING order="10" place="10" resultid="18499" />
                    <RANKING order="11" place="11" resultid="17008" />
                    <RANKING order="12" place="12" resultid="17520" />
                    <RANKING order="13" place="13" resultid="17668" />
                    <RANKING order="14" place="14" resultid="17951" />
                    <RANKING order="15" place="15" resultid="18533" />
                    <RANKING order="16" place="16" resultid="17661" />
                    <RANKING order="17" place="17" resultid="17176" />
                    <RANKING order="18" place="18" resultid="18495" />
                    <RANKING order="19" place="19" resultid="18270" />
                    <RANKING order="20" place="20" resultid="17872" />
                    <RANKING order="21" place="21" resultid="18252" />
                    <RANKING order="22" place="22" resultid="17809" />
                    <RANKING order="23" place="23" resultid="18512" />
                    <RANKING order="24" place="24" resultid="18517" />
                    <RANKING order="25" place="-1" resultid="17865" />
                    <RANKING order="26" place="-1" resultid="18157" />
                    <RANKING order="27" place="-1" resultid="18160" />
                    <RANKING order="28" place="-1" resultid="18166" />
                    <RANKING order="29" place="-1" resultid="18238" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1089" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17060" />
                    <RANKING order="2" place="2" resultid="18312" />
                    <RANKING order="3" place="3" resultid="17183" />
                    <RANKING order="4" place="4" resultid="18043" />
                    <RANKING order="5" place="5" resultid="17549" />
                    <RANKING order="6" place="6" resultid="18550" />
                    <RANKING order="7" place="7" resultid="18424" />
                    <RANKING order="8" place="8" resultid="17216" />
                    <RANKING order="9" place="9" resultid="17682" />
                    <RANKING order="10" place="10" resultid="18231" />
                    <RANKING order="11" place="11" resultid="18169" />
                    <RANKING order="12" place="12" resultid="18555" />
                    <RANKING order="13" place="13" resultid="18017" />
                    <RANKING order="14" place="14" resultid="17195" />
                    <RANKING order="15" place="-1" resultid="18522" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1090" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17223" />
                    <RANKING order="2" place="2" resultid="17343" />
                    <RANKING order="3" place="3" resultid="17492" />
                    <RANKING order="4" place="4" resultid="17381" />
                    <RANKING order="5" place="5" resultid="17388" />
                    <RANKING order="6" place="6" resultid="17421" />
                    <RANKING order="7" place="7" resultid="17400" />
                    <RANKING order="8" place="8" resultid="17060" />
                    <RANKING order="9" place="9" resultid="17394" />
                    <RANKING order="10" place="10" resultid="16984" />
                    <RANKING order="11" place="11" resultid="18223" />
                    <RANKING order="12" place="12" resultid="18312" />
                    <RANKING order="13" place="13" resultid="17188" />
                    <RANKING order="14" place="14" resultid="17183" />
                    <RANKING order="15" place="15" resultid="18043" />
                    <RANKING order="16" place="16" resultid="17549" />
                    <RANKING order="17" place="17" resultid="18151" />
                    <RANKING order="18" place="18" resultid="18550" />
                    <RANKING order="19" place="19" resultid="18424" />
                    <RANKING order="20" place="20" resultid="17236" />
                    <RANKING order="21" place="21" resultid="17216" />
                    <RANKING order="22" place="22" resultid="17415" />
                    <RANKING order="23" place="23" resultid="17682" />
                    <RANKING order="24" place="24" resultid="18231" />
                    <RANKING order="25" place="25" resultid="17879" />
                    <RANKING order="26" place="26" resultid="17528" />
                    <RANKING order="27" place="27" resultid="17555" />
                    <RANKING order="28" place="28" resultid="16960" />
                    <RANKING order="29" place="29" resultid="18169" />
                    <RANKING order="30" place="30" resultid="18555" />
                    <RANKING order="31" place="31" resultid="17506" />
                    <RANKING order="32" place="32" resultid="18031" />
                    <RANKING order="33" place="33" resultid="18017" />
                    <RANKING order="34" place="34" resultid="18499" />
                    <RANKING order="35" place="35" resultid="17008" />
                    <RANKING order="36" place="36" resultid="17520" />
                    <RANKING order="37" place="37" resultid="17668" />
                    <RANKING order="38" place="38" resultid="17951" />
                    <RANKING order="39" place="39" resultid="18533" />
                    <RANKING order="40" place="40" resultid="17661" />
                    <RANKING order="41" place="41" resultid="17176" />
                    <RANKING order="42" place="42" resultid="17195" />
                    <RANKING order="43" place="43" resultid="18495" />
                    <RANKING order="44" place="44" resultid="18270" />
                    <RANKING order="45" place="45" resultid="17872" />
                    <RANKING order="46" place="46" resultid="18252" />
                    <RANKING order="47" place="47" resultid="17809" />
                    <RANKING order="48" place="48" resultid="18512" />
                    <RANKING order="49" place="49" resultid="18517" />
                    <RANKING order="50" place="-1" resultid="17865" />
                    <RANKING order="51" place="-1" resultid="18157" />
                    <RANKING order="52" place="-1" resultid="18160" />
                    <RANKING order="53" place="-1" resultid="18166" />
                    <RANKING order="54" place="-1" resultid="18238" />
                    <RANKING order="55" place="-1" resultid="18522" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="18986" daytime="16:49" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="18987" daytime="16:54" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="18988" daytime="16:58" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="18989" daytime="17:02" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="18990" daytime="17:05" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="18991" daytime="17:08" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1091" daytime="17:17" gender="F" number="9" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1092" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17066" />
                    <RANKING order="2" place="2" resultid="18179" />
                    <RANKING order="3" place="3" resultid="18037" />
                    <RANKING order="4" place="4" resultid="18185" />
                    <RANKING order="5" place="5" resultid="17097" />
                    <RANKING order="6" place="6" resultid="17689" />
                    <RANKING order="7" place="7" resultid="17743" />
                    <RANKING order="8" place="8" resultid="18342" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1093" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18429" />
                    <RANKING order="2" place="2" resultid="17767" />
                    <RANKING order="3" place="3" resultid="17027" />
                    <RANKING order="4" place="4" resultid="18052" />
                    <RANKING order="5" place="5" resultid="18569" />
                    <RANKING order="6" place="6" resultid="17958" />
                    <RANKING order="7" place="7" resultid="18305" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17303" />
                    <RANKING order="2" place="2" resultid="17265" />
                    <RANKING order="3" place="3" resultid="18216" />
                    <RANKING order="4" place="4" resultid="17908" />
                    <RANKING order="5" place="5" resultid="17066" />
                    <RANKING order="6" place="6" resultid="17297" />
                    <RANKING order="7" place="7" resultid="18429" />
                    <RANKING order="8" place="8" resultid="17767" />
                    <RANKING order="9" place="9" resultid="17498" />
                    <RANKING order="10" place="10" resultid="17027" />
                    <RANKING order="11" place="11" resultid="18052" />
                    <RANKING order="12" place="12" resultid="18179" />
                    <RANKING order="13" place="13" resultid="18569" />
                    <RANKING order="14" place="14" resultid="18037" />
                    <RANKING order="15" place="15" resultid="17958" />
                    <RANKING order="16" place="16" resultid="18185" />
                    <RANKING order="17" place="17" resultid="17097" />
                    <RANKING order="18" place="18" resultid="17689" />
                    <RANKING order="19" place="19" resultid="17743" />
                    <RANKING order="20" place="20" resultid="18305" />
                    <RANKING order="21" place="21" resultid="18342" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="18992" daytime="17:17" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="18993" daytime="17:21" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="18994" daytime="17:25" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1095" daytime="17:28" gender="M" number="10" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1096" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17886" />
                    <RANKING order="2" place="2" resultid="17748" />
                    <RANKING order="3" place="3" resultid="17137" />
                    <RANKING order="4" place="4" resultid="18490" />
                    <RANKING order="5" place="5" resultid="17369" />
                    <RANKING order="6" place="6" resultid="18373" />
                    <RANKING order="7" place="7" resultid="17873" />
                    <RANKING order="8" place="8" resultid="18528" />
                    <RANKING order="9" place="-1" resultid="18245" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1097" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17901" />
                    <RANKING order="2" place="2" resultid="18088" />
                    <RANKING order="3" place="3" resultid="18440" />
                    <RANKING order="4" place="4" resultid="17250" />
                    <RANKING order="5" place="5" resultid="17859" />
                    <RANKING order="6" place="6" resultid="17560" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17901" />
                    <RANKING order="2" place="2" resultid="18435" />
                    <RANKING order="3" place="3" resultid="17894" />
                    <RANKING order="4" place="4" resultid="16970" />
                    <RANKING order="5" place="5" resultid="18088" />
                    <RANKING order="6" place="6" resultid="18440" />
                    <RANKING order="7" place="7" resultid="17250" />
                    <RANKING order="8" place="8" resultid="17886" />
                    <RANKING order="9" place="9" resultid="17859" />
                    <RANKING order="10" place="10" resultid="17748" />
                    <RANKING order="11" place="11" resultid="17534" />
                    <RANKING order="12" place="12" resultid="17560" />
                    <RANKING order="13" place="13" resultid="17137" />
                    <RANKING order="14" place="14" resultid="18490" />
                    <RANKING order="15" place="15" resultid="17369" />
                    <RANKING order="16" place="16" resultid="18373" />
                    <RANKING order="17" place="17" resultid="17873" />
                    <RANKING order="18" place="18" resultid="18528" />
                    <RANKING order="19" place="-1" resultid="17579" />
                    <RANKING order="20" place="-1" resultid="18245" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="18995" daytime="17:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="18996" daytime="17:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="18997" daytime="17:37" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1099" daytime="17:46" gender="F" number="11" order="23" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1100" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17143" />
                    <RANKING order="2" place="2" resultid="17710" />
                    <RANKING order="3" place="3" resultid="18024" />
                    <RANKING order="4" place="-1" resultid="18186" />
                    <RANKING order="5" place="-1" resultid="17730" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1101" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17110" />
                    <RANKING order="2" place="2" resultid="17072" />
                    <RANKING order="3" place="3" resultid="18538" />
                    <RANKING order="4" place="4" resultid="17703" />
                    <RANKING order="5" place="5" resultid="18076" />
                    <RANKING order="6" place="-1" resultid="18298" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17110" />
                    <RANKING order="2" place="2" resultid="18333" />
                    <RANKING order="3" place="3" resultid="17056" />
                    <RANKING order="4" place="4" resultid="17072" />
                    <RANKING order="5" place="5" resultid="17486" />
                    <RANKING order="6" place="6" resultid="18538" />
                    <RANKING order="7" place="7" resultid="17703" />
                    <RANKING order="8" place="8" resultid="18076" />
                    <RANKING order="9" place="9" resultid="17143" />
                    <RANKING order="10" place="10" resultid="17710" />
                    <RANKING order="11" place="11" resultid="18024" />
                    <RANKING order="12" place="-1" resultid="18186" />
                    <RANKING order="13" place="-1" resultid="17730" />
                    <RANKING order="14" place="-1" resultid="18298" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="18998" daytime="17:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="18999" daytime="17:54" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1103" daytime="18:01" gender="M" number="12" order="27" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1104" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18176" />
                    <RANKING order="2" place="2" resultid="17131" />
                    <RANKING order="3" place="3" resultid="17880" />
                    <RANKING order="4" place="4" resultid="17723" />
                    <RANKING order="5" place="5" resultid="18319" />
                    <RANKING order="6" place="-1" resultid="17150" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1105" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17830" />
                    <RANKING order="2" place="2" resultid="17737" />
                    <RANKING order="3" place="3" resultid="17573" />
                    <RANKING order="4" place="4" resultid="18070" />
                    <RANKING order="5" place="5" resultid="18044" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1106" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17473" />
                    <RANKING order="2" place="2" resultid="17013" />
                    <RANKING order="3" place="3" resultid="18176" />
                    <RANKING order="4" place="4" resultid="17830" />
                    <RANKING order="5" place="5" resultid="17737" />
                    <RANKING order="6" place="6" resultid="17573" />
                    <RANKING order="7" place="7" resultid="18070" />
                    <RANKING order="8" place="8" resultid="18044" />
                    <RANKING order="9" place="9" resultid="17131" />
                    <RANKING order="10" place="10" resultid="17880" />
                    <RANKING order="11" place="11" resultid="17723" />
                    <RANKING order="12" place="12" resultid="18319" />
                    <RANKING order="13" place="-1" resultid="17150" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19000" daytime="18:01" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19001" daytime="18:09" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6365" daytime="18:28" gender="M" number="13" order="33" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6366" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17866" />
                    <RANKING order="2" place="2" resultid="17887" />
                    <RANKING order="3" place="3" resultid="17356" />
                    <RANKING order="4" place="4" resultid="17749" />
                    <RANKING order="5" place="5" resultid="17844" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6367" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17902" />
                    <RANKING order="2" place="2" resultid="18082" />
                    <RANKING order="3" place="3" resultid="17061" />
                    <RANKING order="4" place="4" resultid="17852" />
                    <RANKING order="5" place="5" resultid="18089" />
                    <RANKING order="6" place="6" resultid="17635" />
                    <RANKING order="7" place="7" resultid="17050" />
                    <RANKING order="8" place="-1" resultid="18523" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6368" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17493" />
                    <RANKING order="2" place="2" resultid="17479" />
                    <RANKING order="3" place="3" resultid="17344" />
                    <RANKING order="4" place="4" resultid="17902" />
                    <RANKING order="5" place="5" resultid="17389" />
                    <RANKING order="6" place="6" resultid="18082" />
                    <RANKING order="7" place="7" resultid="17895" />
                    <RANKING order="8" place="8" resultid="17061" />
                    <RANKING order="9" place="9" resultid="17395" />
                    <RANKING order="10" place="10" resultid="17852" />
                    <RANKING order="11" place="11" resultid="18089" />
                    <RANKING order="12" place="12" resultid="17866" />
                    <RANKING order="13" place="13" resultid="17635" />
                    <RANKING order="14" place="14" resultid="17050" />
                    <RANKING order="15" place="15" resultid="17887" />
                    <RANKING order="16" place="16" resultid="17356" />
                    <RANKING order="17" place="17" resultid="17749" />
                    <RANKING order="18" place="18" resultid="17844" />
                    <RANKING order="19" place="-1" resultid="18523" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19002" daytime="18:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19003" daytime="18:41" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2021-06-19" daytime="09:15" endtime="12:45" name="II BLOK" number="2" warmupfrom="08:45" warmupuntil="09:10">
          <EVENTS>
            <EVENT eventid="1125" daytime="09:15" gender="F" number="14" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1126" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16997" />
                    <RANKING order="2" place="2" resultid="17731" />
                    <RANKING order="3" place="3" resultid="18485" />
                    <RANKING order="4" place="4" resultid="18038" />
                    <RANKING order="5" place="5" resultid="17092" />
                    <RANKING order="6" place="6" resultid="17098" />
                    <RANKING order="7" place="7" resultid="18025" />
                    <RANKING order="8" place="8" resultid="17326" />
                    <RANKING order="9" place="9" resultid="17609" />
                    <RANKING order="10" place="-1" resultid="18478" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1127" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17768" />
                    <RANKING order="2" place="2" resultid="17125" />
                    <RANKING order="3" place="3" resultid="17704" />
                    <RANKING order="4" place="4" resultid="17044" />
                    <RANKING order="5" place="5" resultid="18397" />
                    <RANKING order="6" place="-1" resultid="17697" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1128" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18334" />
                    <RANKING order="2" place="2" resultid="17266" />
                    <RANKING order="3" place="3" resultid="17311" />
                    <RANKING order="4" place="4" resultid="17487" />
                    <RANKING order="5" place="5" resultid="17272" />
                    <RANKING order="6" place="6" resultid="17446" />
                    <RANKING order="7" place="7" resultid="18195" />
                    <RANKING order="8" place="8" resultid="17768" />
                    <RANKING order="9" place="9" resultid="17125" />
                    <RANKING order="10" place="10" resultid="17459" />
                    <RANKING order="11" place="11" resultid="17279" />
                    <RANKING order="12" place="12" resultid="17439" />
                    <RANKING order="13" place="13" resultid="16997" />
                    <RANKING order="14" place="14" resultid="17704" />
                    <RANKING order="15" place="15" resultid="17044" />
                    <RANKING order="16" place="16" resultid="16932" />
                    <RANKING order="17" place="17" resultid="17731" />
                    <RANKING order="18" place="18" resultid="18485" />
                    <RANKING order="19" place="19" resultid="18038" />
                    <RANKING order="20" place="20" resultid="17092" />
                    <RANKING order="21" place="21" resultid="17098" />
                    <RANKING order="22" place="22" resultid="18025" />
                    <RANKING order="23" place="23" resultid="18397" />
                    <RANKING order="24" place="24" resultid="17326" />
                    <RANKING order="25" place="25" resultid="17609" />
                    <RANKING order="26" place="-1" resultid="17697" />
                    <RANKING order="27" place="-1" resultid="18478" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19004" daytime="09:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19005" daytime="09:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19006" daytime="09:29" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19007" daytime="09:35" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1129" daytime="09:40" gender="M" number="15" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1130" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18224" />
                    <RANKING order="2" place="2" resultid="17867" />
                    <RANKING order="3" place="3" resultid="17888" />
                    <RANKING order="4" place="4" resultid="17416" />
                    <RANKING order="5" place="5" resultid="17803" />
                    <RANKING order="6" place="6" resultid="17104" />
                    <RANKING order="7" place="7" resultid="17370" />
                    <RANKING order="8" place="8" resultid="17669" />
                    <RANKING order="9" place="9" resultid="18534" />
                    <RANKING order="10" place="10" resultid="18271" />
                    <RANKING order="11" place="11" resultid="18529" />
                    <RANKING order="12" place="12" resultid="18292" />
                    <RANKING order="13" place="13" resultid="18513" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1131" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17062" />
                    <RANKING order="2" place="2" resultid="18083" />
                    <RANKING order="3" place="3" resultid="17051" />
                    <RANKING order="4" place="4" resultid="18313" />
                    <RANKING order="5" place="5" resultid="17636" />
                    <RANKING order="6" place="6" resultid="18090" />
                    <RANKING order="7" place="7" resultid="17853" />
                    <RANKING order="8" place="8" resultid="18045" />
                    <RANKING order="9" place="9" resultid="18551" />
                    <RANKING order="10" place="10" resultid="18425" />
                    <RANKING order="11" place="11" resultid="17217" />
                    <RANKING order="12" place="-1" resultid="18524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1132" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17224" />
                    <RANKING order="2" place="2" resultid="17494" />
                    <RANKING order="3" place="3" resultid="17345" />
                    <RANKING order="4" place="4" resultid="17382" />
                    <RANKING order="5" place="5" resultid="17422" />
                    <RANKING order="6" place="6" resultid="17480" />
                    <RANKING order="7" place="7" resultid="18436" />
                    <RANKING order="8" place="8" resultid="17390" />
                    <RANKING order="9" place="9" resultid="17396" />
                    <RANKING order="10" place="10" resultid="17062" />
                    <RANKING order="11" place="11" resultid="16985" />
                    <RANKING order="12" place="12" resultid="18083" />
                    <RANKING order="13" place="13" resultid="17401" />
                    <RANKING order="14" place="14" resultid="17051" />
                    <RANKING order="15" place="15" resultid="18224" />
                    <RANKING order="16" place="16" resultid="18313" />
                    <RANKING order="17" place="17" resultid="17636" />
                    <RANKING order="18" place="18" resultid="18090" />
                    <RANKING order="19" place="19" resultid="17853" />
                    <RANKING order="20" place="20" resultid="17867" />
                    <RANKING order="21" place="21" resultid="18045" />
                    <RANKING order="22" place="22" resultid="17896" />
                    <RANKING order="23" place="23" resultid="18551" />
                    <RANKING order="24" place="24" resultid="17888" />
                    <RANKING order="25" place="25" resultid="18425" />
                    <RANKING order="26" place="26" resultid="17416" />
                    <RANKING order="27" place="27" resultid="18361" />
                    <RANKING order="28" place="28" resultid="17217" />
                    <RANKING order="29" place="29" resultid="17529" />
                    <RANKING order="30" place="30" resultid="17803" />
                    <RANKING order="31" place="31" resultid="17104" />
                    <RANKING order="32" place="32" resultid="17370" />
                    <RANKING order="33" place="33" resultid="17669" />
                    <RANKING order="34" place="34" resultid="18534" />
                    <RANKING order="35" place="35" resultid="18271" />
                    <RANKING order="36" place="36" resultid="18529" />
                    <RANKING order="37" place="37" resultid="18292" />
                    <RANKING order="38" place="38" resultid="18513" />
                    <RANKING order="39" place="-1" resultid="18524" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19008" daytime="09:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19009" daytime="09:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19010" daytime="09:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19011" daytime="10:02" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19012" daytime="10:08" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1108" daytime="10:13" gender="F" number="16" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1110" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18180" />
                    <RANKING order="2" place="2" resultid="17144" />
                    <RANKING order="3" place="3" resultid="16998" />
                    <RANKING order="4" place="4" resultid="17718" />
                    <RANKING order="5" place="5" resultid="17320" />
                    <RANKING order="6" place="6" resultid="17093" />
                    <RANKING order="7" place="7" resultid="18110" />
                    <RANKING order="8" place="8" resultid="17744" />
                    <RANKING order="9" place="9" resultid="18343" />
                    <RANKING order="10" place="10" resultid="17156" />
                    <RANKING order="11" place="11" resultid="17615" />
                    <RANKING order="12" place="-1" resultid="18202" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1111" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18059" />
                    <RANKING order="2" place="2" resultid="17085" />
                    <RANKING order="3" place="3" resultid="17028" />
                    <RANKING order="4" place="4" resultid="18077" />
                    <RANKING order="5" place="5" resultid="18327" />
                    <RANKING order="6" place="6" resultid="17959" />
                    <RANKING order="7" place="7" resultid="17824" />
                    <RANKING order="8" place="8" resultid="17045" />
                    <RANKING order="9" place="9" resultid="18539" />
                    <RANKING order="10" place="10" resultid="17033" />
                    <RANKING order="11" place="11" resultid="17589" />
                    <RANKING order="12" place="12" resultid="18368" />
                    <RANKING order="13" place="13" resultid="16922" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1112" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18059" />
                    <RANKING order="2" place="2" resultid="17292" />
                    <RANKING order="3" place="3" resultid="17259" />
                    <RANKING order="4" place="4" resultid="18180" />
                    <RANKING order="5" place="5" resultid="17085" />
                    <RANKING order="6" place="6" resultid="17028" />
                    <RANKING order="7" place="7" resultid="18209" />
                    <RANKING order="8" place="8" resultid="17453" />
                    <RANKING order="9" place="9" resultid="18077" />
                    <RANKING order="10" place="10" resultid="18327" />
                    <RANKING order="11" place="11" resultid="17959" />
                    <RANKING order="12" place="12" resultid="17440" />
                    <RANKING order="13" place="13" resultid="17824" />
                    <RANKING order="14" place="14" resultid="17039" />
                    <RANKING order="15" place="14" resultid="17045" />
                    <RANKING order="16" place="16" resultid="17163" />
                    <RANKING order="17" place="17" resultid="17118" />
                    <RANKING order="18" place="18" resultid="18539" />
                    <RANKING order="19" place="19" resultid="17033" />
                    <RANKING order="20" place="20" resultid="17144" />
                    <RANKING order="21" place="21" resultid="18065" />
                    <RANKING order="22" place="22" resultid="17589" />
                    <RANKING order="23" place="23" resultid="18368" />
                    <RANKING order="24" place="24" resultid="16998" />
                    <RANKING order="25" place="25" resultid="17080" />
                    <RANKING order="26" place="26" resultid="16922" />
                    <RANKING order="27" place="27" resultid="17718" />
                    <RANKING order="28" place="28" resultid="17320" />
                    <RANKING order="29" place="29" resultid="18117" />
                    <RANKING order="30" place="30" resultid="17093" />
                    <RANKING order="31" place="31" resultid="17169" />
                    <RANKING order="32" place="32" resultid="18592" />
                    <RANKING order="33" place="33" resultid="18110" />
                    <RANKING order="34" place="34" resultid="17744" />
                    <RANKING order="35" place="35" resultid="18343" />
                    <RANKING order="36" place="36" resultid="17156" />
                    <RANKING order="37" place="37" resultid="17615" />
                    <RANKING order="38" place="-1" resultid="18202" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19013" daytime="10:13" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19014" daytime="10:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19015" daytime="10:16" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19016" daytime="10:17" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19017" daytime="10:18" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1113" daytime="10:20" gender="M" number="17" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1114" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18225" />
                    <RANKING order="2" place="2" resultid="17881" />
                    <RANKING order="3" place="3" resultid="17804" />
                    <RANKING order="4" place="4" resultid="17132" />
                    <RANKING order="5" place="5" resultid="18032" />
                    <RANKING order="6" place="6" resultid="17237" />
                    <RANKING order="7" place="7" resultid="18607" />
                    <RANKING order="8" place="8" resultid="17724" />
                    <RANKING order="9" place="9" resultid="17556" />
                    <RANKING order="10" place="10" resultid="17357" />
                    <RANKING order="11" place="11" resultid="17676" />
                    <RANKING order="12" place="12" resultid="17952" />
                    <RANKING order="13" place="13" resultid="17521" />
                    <RANKING order="14" place="14" resultid="17204" />
                    <RANKING order="15" place="15" resultid="17662" />
                    <RANKING order="16" place="16" resultid="18500" />
                    <RANKING order="17" place="17" resultid="17810" />
                    <RANKING order="18" place="18" resultid="18374" />
                    <RANKING order="19" place="19" resultid="18253" />
                    <RANKING order="20" place="20" resultid="18496" />
                    <RANKING order="21" place="21" resultid="18285" />
                    <RANKING order="22" place="22" resultid="18239" />
                    <RANKING order="23" place="23" resultid="18518" />
                    <RANKING order="24" place="-1" resultid="17507" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1115" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17903" />
                    <RANKING order="2" place="2" resultid="17738" />
                    <RANKING order="3" place="3" resultid="17838" />
                    <RANKING order="4" place="4" resultid="18084" />
                    <RANKING order="5" place="5" resultid="18264" />
                    <RANKING order="6" place="6" resultid="17230" />
                    <RANKING order="7" place="7" resultid="17185" />
                    <RANKING order="8" place="8" resultid="16956" />
                    <RANKING order="9" place="9" resultid="17574" />
                    <RANKING order="10" place="10" resultid="17854" />
                    <RANKING order="11" place="11" resultid="17550" />
                    <RANKING order="12" place="12" resultid="17251" />
                    <RANKING order="13" place="13" resultid="17860" />
                    <RANKING order="14" place="14" resultid="18355" />
                    <RANKING order="15" place="15" resultid="18046" />
                    <RANKING order="16" place="16" resultid="17789" />
                    <RANKING order="17" place="17" resultid="17683" />
                    <RANKING order="18" place="18" resultid="18426" />
                    <RANKING order="19" place="19" resultid="18071" />
                    <RANKING order="20" place="20" resultid="18232" />
                    <RANKING order="21" place="21" resultid="18018" />
                    <RANKING order="22" place="22" resultid="16952" />
                    <RANKING order="23" place="23" resultid="18556" />
                    <RANKING order="24" place="24" resultid="18007" />
                    <RANKING order="25" place="25" resultid="17984" />
                    <RANKING order="26" place="26" resultid="18417" />
                    <RANKING order="27" place="27" resultid="18170" />
                    <RANKING order="28" place="-1" resultid="17197" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1116" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17338" />
                    <RANKING order="2" place="2" resultid="17225" />
                    <RANKING order="3" place="3" resultid="17474" />
                    <RANKING order="4" place="4" resultid="17546" />
                    <RANKING order="5" place="5" resultid="17432" />
                    <RANKING order="6" place="6" resultid="17565" />
                    <RANKING order="7" place="7" resultid="17210" />
                    <RANKING order="8" place="8" resultid="17903" />
                    <RANKING order="9" place="9" resultid="17022" />
                    <RANKING order="10" place="10" resultid="17465" />
                    <RANKING order="11" place="11" resultid="17738" />
                    <RANKING order="12" place="12" resultid="16971" />
                    <RANKING order="13" place="13" resultid="17838" />
                    <RANKING order="14" place="14" resultid="18084" />
                    <RANKING order="15" place="15" resultid="18135" />
                    <RANKING order="16" place="16" resultid="17541" />
                    <RANKING order="17" place="17" resultid="18264" />
                    <RANKING order="18" place="18" resultid="16986" />
                    <RANKING order="19" place="19" resultid="17230" />
                    <RANKING order="20" place="20" resultid="17185" />
                    <RANKING order="21" place="21" resultid="16956" />
                    <RANKING order="22" place="22" resultid="17469" />
                    <RANKING order="23" place="23" resultid="17190" />
                    <RANKING order="24" place="24" resultid="17574" />
                    <RANKING order="25" place="25" resultid="18225" />
                    <RANKING order="26" place="26" resultid="17854" />
                    <RANKING order="27" place="27" resultid="17550" />
                    <RANKING order="28" place="28" resultid="17251" />
                    <RANKING order="29" place="29" resultid="17860" />
                    <RANKING order="30" place="30" resultid="18355" />
                    <RANKING order="31" place="31" resultid="17881" />
                    <RANKING order="32" place="31" resultid="18046" />
                    <RANKING order="33" place="33" resultid="17804" />
                    <RANKING order="34" place="34" resultid="17132" />
                    <RANKING order="35" place="35" resultid="17789" />
                    <RANKING order="36" place="36" resultid="17683" />
                    <RANKING order="37" place="37" resultid="18426" />
                    <RANKING order="38" place="38" resultid="18071" />
                    <RANKING order="39" place="39" resultid="18232" />
                    <RANKING order="40" place="40" resultid="17530" />
                    <RANKING order="41" place="41" resultid="18018" />
                    <RANKING order="42" place="42" resultid="16952" />
                    <RANKING order="43" place="43" resultid="18032" />
                    <RANKING order="44" place="44" resultid="17237" />
                    <RANKING order="45" place="45" resultid="18607" />
                    <RANKING order="46" place="46" resultid="17724" />
                    <RANKING order="47" place="47" resultid="17556" />
                    <RANKING order="48" place="48" resultid="18556" />
                    <RANKING order="49" place="49" resultid="17357" />
                    <RANKING order="50" place="50" resultid="18007" />
                    <RANKING order="51" place="51" resultid="17676" />
                    <RANKING order="52" place="52" resultid="17952" />
                    <RANKING order="53" place="53" resultid="17521" />
                    <RANKING order="54" place="54" resultid="17984" />
                    <RANKING order="55" place="55" resultid="17204" />
                    <RANKING order="56" place="56" resultid="18417" />
                    <RANKING order="57" place="57" resultid="18170" />
                    <RANKING order="58" place="58" resultid="17662" />
                    <RANKING order="59" place="59" resultid="18500" />
                    <RANKING order="60" place="60" resultid="17810" />
                    <RANKING order="61" place="61" resultid="18374" />
                    <RANKING order="62" place="62" resultid="18253" />
                    <RANKING order="63" place="63" resultid="18496" />
                    <RANKING order="64" place="64" resultid="18285" />
                    <RANKING order="65" place="65" resultid="18239" />
                    <RANKING order="66" place="66" resultid="18518" />
                    <RANKING order="67" place="-1" resultid="17197" />
                    <RANKING order="68" place="-1" resultid="16883" />
                    <RANKING order="69" place="-1" resultid="17507" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19018" daytime="10:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19019" daytime="10:21" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19020" daytime="10:23" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19021" daytime="10:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19022" daytime="10:26" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19023" daytime="10:27" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19024" daytime="10:29" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19025" daytime="10:30" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1117" daytime="10:37" gender="F" number="18" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1118" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17067" />
                    <RANKING order="2" place="2" resultid="18039" />
                    <RANKING order="3" place="3" resultid="16911" />
                    <RANKING order="4" place="4" resultid="16917" />
                    <RANKING order="5" place="5" resultid="17711" />
                    <RANKING order="6" place="6" resultid="17099" />
                    <RANKING order="7" place="7" resultid="18401" />
                    <RANKING order="8" place="8" resultid="17690" />
                    <RANKING order="9" place="9" resultid="17745" />
                    <RANKING order="10" place="10" resultid="17603" />
                    <RANKING order="11" place="11" resultid="18350" />
                    <RANKING order="12" place="12" resultid="17932" />
                    <RANKING order="13" place="13" resultid="17945" />
                    <RANKING order="14" place="14" resultid="18103" />
                    <RANKING order="15" place="15" resultid="18344" />
                    <RANKING order="16" place="16" resultid="18130" />
                    <RANKING order="17" place="-1" resultid="18181" />
                    <RANKING order="18" place="-1" resultid="18203" />
                    <RANKING order="19" place="-1" resultid="18479" />
                    <RANKING order="20" place="-1" resultid="18618" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1119" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17111" />
                    <RANKING order="2" place="2" resultid="17029" />
                    <RANKING order="3" place="3" resultid="18053" />
                    <RANKING order="4" place="4" resultid="18430" />
                    <RANKING order="5" place="5" resultid="18570" />
                    <RANKING order="6" place="6" resultid="18546" />
                    <RANKING order="7" place="7" resultid="18369" />
                    <RANKING order="8" place="8" resultid="18306" />
                    <RANKING order="9" place="9" resultid="18123" />
                    <RANKING order="10" place="10" resultid="17925" />
                    <RANKING order="11" place="-1" resultid="18392" />
                    <RANKING order="12" place="-1" resultid="19101" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1120" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17111" />
                    <RANKING order="2" place="2" resultid="18217" />
                    <RANKING order="3" place="3" resultid="17293" />
                    <RANKING order="4" place="4" resultid="17285" />
                    <RANKING order="5" place="5" resultid="18210" />
                    <RANKING order="6" place="6" resultid="17273" />
                    <RANKING order="7" place="7" resultid="17029" />
                    <RANKING order="8" place="8" resultid="17298" />
                    <RANKING order="9" place="9" resultid="17909" />
                    <RANKING order="10" place="10" resultid="17067" />
                    <RANKING order="11" place="11" resultid="18053" />
                    <RANKING order="12" place="12" resultid="17499" />
                    <RANKING order="13" place="13" resultid="18430" />
                    <RANKING order="14" place="14" resultid="18039" />
                    <RANKING order="15" place="15" resultid="16926" />
                    <RANKING order="16" place="16" resultid="18570" />
                    <RANKING order="17" place="17" resultid="18546" />
                    <RANKING order="18" place="18" resultid="16911" />
                    <RANKING order="19" place="19" resultid="17167" />
                    <RANKING order="20" place="20" resultid="17040" />
                    <RANKING order="21" place="21" resultid="16917" />
                    <RANKING order="22" place="22" resultid="17711" />
                    <RANKING order="23" place="23" resultid="17099" />
                    <RANKING order="24" place="24" resultid="18401" />
                    <RANKING order="25" place="25" resultid="17690" />
                    <RANKING order="26" place="26" resultid="17745" />
                    <RANKING order="27" place="27" resultid="18369" />
                    <RANKING order="28" place="28" resultid="18306" />
                    <RANKING order="29" place="29" resultid="17603" />
                    <RANKING order="30" place="30" resultid="17173" />
                    <RANKING order="31" place="31" resultid="18350" />
                    <RANKING order="32" place="32" resultid="18123" />
                    <RANKING order="33" place="33" resultid="17932" />
                    <RANKING order="34" place="34" resultid="17945" />
                    <RANKING order="35" place="35" resultid="18118" />
                    <RANKING order="36" place="36" resultid="18103" />
                    <RANKING order="37" place="37" resultid="17925" />
                    <RANKING order="38" place="37" resultid="18344" />
                    <RANKING order="39" place="39" resultid="17585" />
                    <RANKING order="40" place="40" resultid="18130" />
                    <RANKING order="41" place="-1" resultid="18181" />
                    <RANKING order="42" place="-1" resultid="17454" />
                    <RANKING order="43" place="-1" resultid="18203" />
                    <RANKING order="44" place="-1" resultid="18392" />
                    <RANKING order="45" place="-1" resultid="18479" />
                    <RANKING order="46" place="-1" resultid="18618" />
                    <RANKING order="47" place="-1" resultid="19101" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19026" daytime="10:37" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19027" daytime="10:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19028" daytime="10:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19029" daytime="10:41" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19030" daytime="10:43" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1121" daytime="10:44" gender="M" number="19" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1122" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17868" />
                    <RANKING order="2" place="2" resultid="17151" />
                    <RANKING order="3" place="3" resultid="17889" />
                    <RANKING order="4" place="4" resultid="17882" />
                    <RANKING order="5" place="5" resultid="17750" />
                    <RANKING order="6" place="6" resultid="17238" />
                    <RANKING order="7" place="7" resultid="17417" />
                    <RANKING order="8" place="8" resultid="17138" />
                    <RANKING order="9" place="9" resultid="18491" />
                    <RANKING order="10" place="10" resultid="17371" />
                    <RANKING order="11" place="11" resultid="17179" />
                    <RANKING order="12" place="12" resultid="17244" />
                    <RANKING order="13" place="13" resultid="17376" />
                    <RANKING order="14" place="14" resultid="17009" />
                    <RANKING order="15" place="15" resultid="18597" />
                    <RANKING order="16" place="16" resultid="17514" />
                    <RANKING order="17" place="17" resultid="17663" />
                    <RANKING order="18" place="18" resultid="18535" />
                    <RANKING order="19" place="19" resultid="16946" />
                    <RANKING order="20" place="20" resultid="18000" />
                    <RANKING order="21" place="21" resultid="18254" />
                    <RANKING order="22" place="22" resultid="18272" />
                    <RANKING order="23" place="23" resultid="17874" />
                    <RANKING order="24" place="24" resultid="17670" />
                    <RANKING order="25" place="25" resultid="18293" />
                    <RANKING order="26" place="26" resultid="17817" />
                    <RANKING order="27" place="27" resultid="17350" />
                    <RANKING order="28" place="28" resultid="18530" />
                    <RANKING order="29" place="29" resultid="18013" />
                    <RANKING order="30" place="30" resultid="18514" />
                    <RANKING order="31" place="31" resultid="17995" />
                    <RANKING order="32" place="32" resultid="18240" />
                    <RANKING order="33" place="33" resultid="17763" />
                    <RANKING order="34" place="34" resultid="17759" />
                    <RANKING order="35" place="-1" resultid="17508" />
                    <RANKING order="36" place="-1" resultid="17657" />
                    <RANKING order="37" place="-1" resultid="17755" />
                    <RANKING order="38" place="-1" resultid="17761" />
                    <RANKING order="39" place="-1" resultid="18246" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1123" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17252" />
                    <RANKING order="2" place="2" resultid="17231" />
                    <RANKING order="3" place="3" resultid="18091" />
                    <RANKING order="4" place="4" resultid="16978" />
                    <RANKING order="5" place="5" resultid="17218" />
                    <RANKING order="6" place="6" resultid="17637" />
                    <RANKING order="7" place="7" resultid="18441" />
                    <RANKING order="8" place="8" resultid="17561" />
                    <RANKING order="9" place="9" resultid="17861" />
                    <RANKING order="10" place="10" resultid="18411" />
                    <RANKING order="11" place="11" resultid="18356" />
                    <RANKING order="12" place="12" resultid="18506" />
                    <RANKING order="13" place="13" resultid="16953" />
                    <RANKING order="14" place="14" resultid="18019" />
                    <RANKING order="15" place="15" resultid="18171" />
                    <RANKING order="16" place="16" resultid="17198" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1124" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17339" />
                    <RANKING order="2" place="2" resultid="17191" />
                    <RANKING order="3" place="3" resultid="17897" />
                    <RANKING order="4" place="4" resultid="17211" />
                    <RANKING order="5" place="5" resultid="17252" />
                    <RANKING order="6" place="6" resultid="17231" />
                    <RANKING order="7" place="7" resultid="16972" />
                    <RANKING order="8" place="8" resultid="18091" />
                    <RANKING order="9" place="9" resultid="16978" />
                    <RANKING order="10" place="10" resultid="17621" />
                    <RANKING order="11" place="11" resultid="17218" />
                    <RANKING order="12" place="12" resultid="17868" />
                    <RANKING order="13" place="13" resultid="17637" />
                    <RANKING order="14" place="14" resultid="18441" />
                    <RANKING order="15" place="15" resultid="17151" />
                    <RANKING order="16" place="16" resultid="17889" />
                    <RANKING order="17" place="17" resultid="17882" />
                    <RANKING order="18" place="18" resultid="17561" />
                    <RANKING order="19" place="19" resultid="17535" />
                    <RANKING order="20" place="20" resultid="17750" />
                    <RANKING order="21" place="21" resultid="17861" />
                    <RANKING order="22" place="22" resultid="17238" />
                    <RANKING order="23" place="23" resultid="18411" />
                    <RANKING order="24" place="24" resultid="18356" />
                    <RANKING order="25" place="25" resultid="17417" />
                    <RANKING order="26" place="26" resultid="18506" />
                    <RANKING order="27" place="27" resultid="16953" />
                    <RANKING order="28" place="28" resultid="18019" />
                    <RANKING order="29" place="29" resultid="17138" />
                    <RANKING order="30" place="30" resultid="18491" />
                    <RANKING order="31" place="31" resultid="17371" />
                    <RANKING order="32" place="32" resultid="17179" />
                    <RANKING order="33" place="33" resultid="18171" />
                    <RANKING order="34" place="34" resultid="17244" />
                    <RANKING order="35" place="35" resultid="17376" />
                    <RANKING order="36" place="36" resultid="17009" />
                    <RANKING order="37" place="37" resultid="18597" />
                    <RANKING order="38" place="38" resultid="17514" />
                    <RANKING order="39" place="39" resultid="17198" />
                    <RANKING order="40" place="40" resultid="17663" />
                    <RANKING order="41" place="41" resultid="18535" />
                    <RANKING order="42" place="42" resultid="16946" />
                    <RANKING order="43" place="43" resultid="18000" />
                    <RANKING order="44" place="44" resultid="18254" />
                    <RANKING order="45" place="45" resultid="18272" />
                    <RANKING order="46" place="46" resultid="17874" />
                    <RANKING order="47" place="47" resultid="17670" />
                    <RANKING order="48" place="48" resultid="18293" />
                    <RANKING order="49" place="49" resultid="17817" />
                    <RANKING order="50" place="50" resultid="17350" />
                    <RANKING order="51" place="51" resultid="18530" />
                    <RANKING order="52" place="52" resultid="18013" />
                    <RANKING order="53" place="53" resultid="18514" />
                    <RANKING order="54" place="54" resultid="17995" />
                    <RANKING order="55" place="55" resultid="18240" />
                    <RANKING order="56" place="56" resultid="17763" />
                    <RANKING order="57" place="57" resultid="17759" />
                    <RANKING order="58" place="-1" resultid="17652" />
                    <RANKING order="59" place="-1" resultid="17508" />
                    <RANKING order="60" place="-1" resultid="17580" />
                    <RANKING order="61" place="-1" resultid="17657" />
                    <RANKING order="62" place="-1" resultid="17755" />
                    <RANKING order="63" place="-1" resultid="17761" />
                    <RANKING order="64" place="-1" resultid="18246" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19031" daytime="10:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19032" daytime="10:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19033" daytime="10:47" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19034" daytime="10:48" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19035" daytime="10:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19036" daytime="10:51" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19037" daytime="10:53" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1133" daytime="11:00" gender="F" number="20" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1134" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16992" />
                    <RANKING order="2" place="2" resultid="17691" />
                    <RANKING order="3" place="3" resultid="18187" />
                    <RANKING order="4" place="4" resultid="17610" />
                    <RANKING order="5" place="5" resultid="17160" />
                    <RANKING order="6" place="6" resultid="17933" />
                    <RANKING order="7" place="7" resultid="17946" />
                    <RANKING order="8" place="-1" resultid="17321" />
                    <RANKING order="9" place="-1" resultid="18104" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1135" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17705" />
                    <RANKING order="2" place="2" resultid="17825" />
                    <RANKING order="3" place="3" resultid="17126" />
                    <RANKING order="4" place="4" resultid="18567" />
                    <RANKING order="5" place="5" resultid="17086" />
                    <RANKING order="6" place="6" resultid="18054" />
                    <RANKING order="7" place="7" resultid="18299" />
                    <RANKING order="8" place="8" resultid="17034" />
                    <RANKING order="9" place="9" resultid="17004" />
                    <RANKING order="10" place="10" resultid="18307" />
                    <RANKING order="11" place="11" resultid="18124" />
                    <RANKING order="12" place="12" resultid="17926" />
                    <RANKING order="13" place="-1" resultid="17590" />
                    <RANKING order="14" place="-1" resultid="17598" />
                    <RANKING order="15" place="-1" resultid="17698" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1136" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17406" />
                    <RANKING order="2" place="2" resultid="17409" />
                    <RANKING order="3" place="3" resultid="17705" />
                    <RANKING order="4" place="4" resultid="17825" />
                    <RANKING order="5" place="5" resultid="17126" />
                    <RANKING order="6" place="6" resultid="18567" />
                    <RANKING order="7" place="7" resultid="16992" />
                    <RANKING order="8" place="8" resultid="17086" />
                    <RANKING order="9" place="9" resultid="18054" />
                    <RANKING order="10" place="10" resultid="18066" />
                    <RANKING order="11" place="11" resultid="18299" />
                    <RANKING order="12" place="12" resultid="17119" />
                    <RANKING order="13" place="13" resultid="17034" />
                    <RANKING order="14" place="14" resultid="17004" />
                    <RANKING order="15" place="15" resultid="17691" />
                    <RANKING order="16" place="16" resultid="18187" />
                    <RANKING order="17" place="17" resultid="18307" />
                    <RANKING order="18" place="18" resultid="18124" />
                    <RANKING order="19" place="19" resultid="17610" />
                    <RANKING order="20" place="20" resultid="17160" />
                    <RANKING order="21" place="21" resultid="17926" />
                    <RANKING order="22" place="22" resultid="17933" />
                    <RANKING order="23" place="23" resultid="17946" />
                    <RANKING order="24" place="-1" resultid="17590" />
                    <RANKING order="25" place="-1" resultid="17321" />
                    <RANKING order="26" place="-1" resultid="18104" />
                    <RANKING order="27" place="-1" resultid="17598" />
                    <RANKING order="28" place="-1" resultid="17698" />
                    <RANKING order="29" place="-1" resultid="18335" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19038" daytime="11:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19039" daytime="11:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19040" daytime="11:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19041" daytime="11:07" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1137" daytime="11:09" gender="M" number="21" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1138" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17133" />
                    <RANKING order="2" place="2" resultid="17845" />
                    <RANKING order="3" place="3" resultid="17725" />
                    <RANKING order="4" place="4" resultid="17205" />
                    <RANKING order="5" place="5" resultid="16961" />
                    <RANKING order="6" place="6" resultid="18615" />
                    <RANKING order="7" place="7" resultid="17796" />
                    <RANKING order="8" place="8" resultid="17953" />
                    <RANKING order="9" place="9" resultid="17377" />
                    <RANKING order="10" place="10" resultid="17522" />
                    <RANKING order="11" place="11" resultid="17178" />
                    <RANKING order="12" place="12" resultid="18320" />
                    <RANKING order="13" place="13" resultid="18375" />
                    <RANKING order="14" place="14" resultid="17245" />
                    <RANKING order="15" place="15" resultid="17363" />
                    <RANKING order="16" place="16" resultid="18611" />
                    <RANKING order="17" place="17" resultid="17105" />
                    <RANKING order="18" place="18" resultid="18001" />
                    <RANKING order="19" place="19" resultid="17875" />
                    <RANKING order="20" place="20" resultid="17351" />
                    <RANKING order="21" place="21" resultid="17818" />
                    <RANKING order="22" place="22" resultid="17515" />
                    <RANKING order="23" place="23" resultid="17811" />
                    <RANKING order="24" place="24" resultid="18278" />
                    <RANKING order="25" place="25" resultid="18519" />
                    <RANKING order="26" place="-1" resultid="17677" />
                    <RANKING order="27" place="-1" resultid="16966" />
                    <RANKING order="28" place="-1" resultid="17010" />
                    <RANKING order="29" place="-1" resultid="17990" />
                    <RANKING order="30" place="-1" resultid="18247" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1139" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17643" />
                    <RANKING order="2" place="2" resultid="17839" />
                    <RANKING order="3" place="3" resultid="17831" />
                    <RANKING order="4" place="4" resultid="18072" />
                    <RANKING order="5" place="5" resultid="16957" />
                    <RANKING order="6" place="6" resultid="17569" />
                    <RANKING order="7" place="7" resultid="16979" />
                    <RANKING order="8" place="8" resultid="18507" />
                    <RANKING order="9" place="9" resultid="17018" />
                    <RANKING order="10" place="10" resultid="17790" />
                    <RANKING order="11" place="11" resultid="18314" />
                    <RANKING order="12" place="12" resultid="18412" />
                    <RANKING order="13" place="13" resultid="17632" />
                    <RANKING order="14" place="14" resultid="18008" />
                    <RANKING order="15" place="15" resultid="18233" />
                    <RANKING order="16" place="16" resultid="18561" />
                    <RANKING order="17" place="-1" resultid="17985" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1140" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17433" />
                    <RANKING order="2" place="2" resultid="17428" />
                    <RANKING order="3" place="3" resultid="17023" />
                    <RANKING order="4" place="4" resultid="17423" />
                    <RANKING order="5" place="5" resultid="17643" />
                    <RANKING order="6" place="6" resultid="17839" />
                    <RANKING order="7" place="7" resultid="18136" />
                    <RANKING order="8" place="8" resultid="17831" />
                    <RANKING order="9" place="9" resultid="18072" />
                    <RANKING order="10" place="10" resultid="16957" />
                    <RANKING order="11" place="11" resultid="17133" />
                    <RANKING order="12" place="12" resultid="17569" />
                    <RANKING order="13" place="13" resultid="17845" />
                    <RANKING order="14" place="14" resultid="16979" />
                    <RANKING order="15" place="15" resultid="18507" />
                    <RANKING order="16" place="16" resultid="17018" />
                    <RANKING order="17" place="17" resultid="17790" />
                    <RANKING order="18" place="18" resultid="18314" />
                    <RANKING order="19" place="19" resultid="18412" />
                    <RANKING order="20" place="20" resultid="17632" />
                    <RANKING order="21" place="21" resultid="17725" />
                    <RANKING order="22" place="22" resultid="17205" />
                    <RANKING order="23" place="23" resultid="16961" />
                    <RANKING order="24" place="24" resultid="18615" />
                    <RANKING order="25" place="25" resultid="18008" />
                    <RANKING order="26" place="26" resultid="17796" />
                    <RANKING order="27" place="27" resultid="17953" />
                    <RANKING order="28" place="28" resultid="17377" />
                    <RANKING order="29" place="29" resultid="18233" />
                    <RANKING order="30" place="30" resultid="18561" />
                    <RANKING order="31" place="31" resultid="17522" />
                    <RANKING order="32" place="32" resultid="17178" />
                    <RANKING order="33" place="33" resultid="18320" />
                    <RANKING order="34" place="34" resultid="18375" />
                    <RANKING order="35" place="35" resultid="17245" />
                    <RANKING order="36" place="36" resultid="17363" />
                    <RANKING order="37" place="37" resultid="18611" />
                    <RANKING order="38" place="38" resultid="17105" />
                    <RANKING order="39" place="39" resultid="18001" />
                    <RANKING order="40" place="40" resultid="17875" />
                    <RANKING order="41" place="41" resultid="17351" />
                    <RANKING order="42" place="42" resultid="17818" />
                    <RANKING order="43" place="43" resultid="17515" />
                    <RANKING order="44" place="44" resultid="17811" />
                    <RANKING order="45" place="45" resultid="18278" />
                    <RANKING order="46" place="46" resultid="18519" />
                    <RANKING order="47" place="-1" resultid="17677" />
                    <RANKING order="48" place="-1" resultid="17985" />
                    <RANKING order="49" place="-1" resultid="16966" />
                    <RANKING order="50" place="-1" resultid="17010" />
                    <RANKING order="51" place="-1" resultid="17627" />
                    <RANKING order="52" place="-1" resultid="17990" />
                    <RANKING order="53" place="-1" resultid="18247" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19042" daytime="11:09" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19043" daytime="11:12" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19044" daytime="11:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19045" daytime="11:18" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19046" daytime="11:21" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19047" daytime="11:23" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1141" daytime="11:31" gender="F" number="22" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1142" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17068" />
                    <RANKING order="2" place="2" resultid="18188" />
                    <RANKING order="3" place="3" resultid="17145" />
                    <RANKING order="4" place="4" resultid="17712" />
                    <RANKING order="5" place="5" resultid="17732" />
                    <RANKING order="6" place="6" resultid="18026" />
                    <RANKING order="7" place="7" resultid="17719" />
                    <RANKING order="8" place="8" resultid="17327" />
                    <RANKING order="9" place="9" resultid="18111" />
                    <RANKING order="10" place="10" resultid="17616" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1143" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17112" />
                    <RANKING order="2" place="2" resultid="17073" />
                    <RANKING order="3" place="3" resultid="18540" />
                    <RANKING order="4" place="4" resultid="18431" />
                    <RANKING order="5" place="5" resultid="18328" />
                    <RANKING order="6" place="6" resultid="18300" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1144" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17112" />
                    <RANKING order="2" place="2" resultid="17260" />
                    <RANKING order="3" place="3" resultid="18336" />
                    <RANKING order="4" place="4" resultid="17057" />
                    <RANKING order="5" place="5" resultid="18218" />
                    <RANKING order="6" place="6" resultid="17073" />
                    <RANKING order="7" place="7" resultid="17447" />
                    <RANKING order="8" place="8" resultid="17286" />
                    <RANKING order="9" place="9" resultid="17488" />
                    <RANKING order="10" place="10" resultid="17910" />
                    <RANKING order="11" place="11" resultid="17500" />
                    <RANKING order="12" place="12" resultid="17410" />
                    <RANKING order="13" place="13" resultid="18540" />
                    <RANKING order="14" place="14" resultid="17068" />
                    <RANKING order="15" place="15" resultid="17299" />
                    <RANKING order="16" place="16" resultid="18431" />
                    <RANKING order="17" place="17" resultid="18328" />
                    <RANKING order="18" place="18" resultid="18188" />
                    <RANKING order="19" place="19" resultid="18300" />
                    <RANKING order="20" place="20" resultid="17145" />
                    <RANKING order="21" place="21" resultid="17712" />
                    <RANKING order="22" place="22" resultid="17732" />
                    <RANKING order="23" place="23" resultid="18026" />
                    <RANKING order="24" place="24" resultid="17719" />
                    <RANKING order="25" place="25" resultid="17327" />
                    <RANKING order="26" place="26" resultid="18111" />
                    <RANKING order="27" place="27" resultid="17616" />
                    <RANKING order="28" place="-1" resultid="18211" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19048" daytime="11:31" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19049" daytime="11:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19050" daytime="11:38" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1145" daytime="11:42" gender="M" number="23" order="24" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1146" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17152" />
                    <RANKING order="2" place="2" resultid="17846" />
                    <RANKING order="3" place="3" resultid="17751" />
                    <RANKING order="4" place="4" resultid="17358" />
                    <RANKING order="5" place="5" resultid="18492" />
                    <RANKING order="6" place="6" resultid="18033" />
                    <RANKING order="7" place="7" resultid="18321" />
                    <RANKING order="8" place="8" resultid="18501" />
                    <RANKING order="9" place="9" resultid="17797" />
                    <RANKING order="10" place="10" resultid="17364" />
                    <RANKING order="11" place="11" resultid="18598" />
                    <RANKING order="12" place="12" resultid="18279" />
                    <RANKING order="13" place="13" resultid="18286" />
                    <RANKING order="14" place="-1" resultid="17139" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1147" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17905" />
                    <RANKING order="2" place="2" resultid="17832" />
                    <RANKING order="3" place="3" resultid="17644" />
                    <RANKING order="4" place="4" resultid="17739" />
                    <RANKING order="5" place="5" resultid="17575" />
                    <RANKING order="6" place="6" resultid="18265" />
                    <RANKING order="7" place="7" resultid="17684" />
                    <RANKING order="8" place="-1" resultid="17551" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1148" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17434" />
                    <RANKING order="2" place="2" resultid="17383" />
                    <RANKING order="3" place="3" resultid="17475" />
                    <RANKING order="4" place="4" resultid="17481" />
                    <RANKING order="5" place="5" resultid="17905" />
                    <RANKING order="6" place="6" resultid="17014" />
                    <RANKING order="7" place="7" resultid="17832" />
                    <RANKING order="8" place="8" resultid="17644" />
                    <RANKING order="9" place="9" resultid="17739" />
                    <RANKING order="10" place="10" resultid="17152" />
                    <RANKING order="11" place="11" resultid="17575" />
                    <RANKING order="12" place="12" resultid="18265" />
                    <RANKING order="13" place="13" resultid="18362" />
                    <RANKING order="14" place="14" resultid="17684" />
                    <RANKING order="15" place="15" resultid="17846" />
                    <RANKING order="16" place="16" resultid="17751" />
                    <RANKING order="17" place="17" resultid="17358" />
                    <RANKING order="18" place="18" resultid="17536" />
                    <RANKING order="19" place="19" resultid="18492" />
                    <RANKING order="20" place="20" resultid="18033" />
                    <RANKING order="21" place="21" resultid="18321" />
                    <RANKING order="22" place="22" resultid="18501" />
                    <RANKING order="23" place="23" resultid="17797" />
                    <RANKING order="24" place="24" resultid="17364" />
                    <RANKING order="25" place="25" resultid="18598" />
                    <RANKING order="26" place="26" resultid="18279" />
                    <RANKING order="27" place="27" resultid="18286" />
                    <RANKING order="28" place="-1" resultid="17551" />
                    <RANKING order="29" place="-1" resultid="17139" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19051" daytime="11:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19052" daytime="11:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19053" daytime="11:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19054" daytime="11:53" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6361" daytime="12:09" gender="F" number="24" order="29" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6363" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17769" />
                    <RANKING order="2" place="-1" resultid="18574" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6364" agemax="-1" agemin="14" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18196" />
                    <RANKING order="2" place="2" resultid="17769" />
                    <RANKING order="3" place="-1" resultid="18574" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19055" daytime="12:09" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2021-06-19" daytime="15:30" endtime="19:14" name="III BLOK" number="3" warmupfrom="15:00" warmupuntil="15:25">
          <EVENTS>
            <EVENT eventid="1150" daytime="15:30" gender="F" number="25" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1152" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17069" />
                    <RANKING order="2" place="2" resultid="18027" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1153" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17074" />
                    <RANKING order="2" place="2" resultid="18078" />
                    <RANKING order="3" place="3" resultid="18329" />
                    <RANKING order="4" place="4" resultid="17960" />
                    <RANKING order="5" place="-1" resultid="17035" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1154" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17441" />
                    <RANKING order="2" place="2" resultid="17455" />
                    <RANKING order="3" place="3" resultid="17074" />
                    <RANKING order="4" place="4" resultid="17448" />
                    <RANKING order="5" place="5" resultid="18067" />
                    <RANKING order="6" place="6" resultid="17069" />
                    <RANKING order="7" place="7" resultid="18078" />
                    <RANKING order="8" place="8" resultid="18329" />
                    <RANKING order="9" place="9" resultid="17960" />
                    <RANKING order="10" place="10" resultid="18027" />
                    <RANKING order="11" place="-1" resultid="17035" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19056" daytime="15:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19057" daytime="15:34" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1155" daytime="15:38" gender="M" number="26" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1156" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17805" />
                    <RANKING order="2" place="2" resultid="17106" />
                    <RANKING order="3" place="3" resultid="17359" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1157" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18085" />
                    <RANKING order="2" place="2" resultid="17576" />
                    <RANKING order="3" place="3" resultid="17052" />
                    <RANKING order="4" place="4" resultid="17862" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1158" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17482" />
                    <RANKING order="2" place="2" resultid="17470" />
                    <RANKING order="3" place="3" resultid="18437" />
                    <RANKING order="4" place="4" resultid="16987" />
                    <RANKING order="5" place="5" resultid="18085" />
                    <RANKING order="6" place="6" resultid="17576" />
                    <RANKING order="7" place="7" resultid="17052" />
                    <RANKING order="8" place="8" resultid="17805" />
                    <RANKING order="9" place="9" resultid="17862" />
                    <RANKING order="10" place="10" resultid="17106" />
                    <RANKING order="11" place="11" resultid="17359" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19058" daytime="15:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19059" daytime="15:42" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1159" daytime="15:45" gender="F" number="27" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1160" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16912" />
                    <RANKING order="2" place="2" resultid="18182" />
                    <RANKING order="3" place="3" resultid="16918" />
                    <RANKING order="4" place="4" resultid="18486" />
                    <RANKING order="5" place="5" resultid="17094" />
                    <RANKING order="6" place="6" resultid="18402" />
                    <RANKING order="7" place="7" resultid="17322" />
                    <RANKING order="8" place="8" resultid="17604" />
                    <RANKING order="9" place="9" resultid="17146" />
                    <RANKING order="10" place="10" resultid="17611" />
                    <RANKING order="11" place="11" resultid="17328" />
                    <RANKING order="12" place="12" resultid="18345" />
                    <RANKING order="13" place="13" resultid="18351" />
                    <RANKING order="14" place="14" resultid="18105" />
                    <RANKING order="15" place="15" resultid="17157" />
                    <RANKING order="16" place="16" resultid="17947" />
                    <RANKING order="17" place="17" resultid="18112" />
                    <RANKING order="18" place="18" resultid="17617" />
                    <RANKING order="19" place="19" resultid="17934" />
                    <RANKING order="20" place="20" resultid="18131" />
                    <RANKING order="21" place="-1" resultid="18204" />
                    <RANKING order="22" place="-1" resultid="18480" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1161" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18060" />
                    <RANKING order="2" place="2" resultid="17113" />
                    <RANKING order="3" place="3" resultid="17826" />
                    <RANKING order="4" place="4" resultid="17087" />
                    <RANKING order="5" place="5" resultid="18432" />
                    <RANKING order="6" place="6" resultid="17127" />
                    <RANKING order="7" place="7" resultid="16923" />
                    <RANKING order="8" place="8" resultid="17706" />
                    <RANKING order="9" place="9" resultid="17961" />
                    <RANKING order="10" place="10" resultid="17005" />
                    <RANKING order="11" place="11" resultid="18330" />
                    <RANKING order="12" place="12" resultid="18547" />
                    <RANKING order="13" place="13" resultid="18370" />
                    <RANKING order="14" place="14" resultid="18398" />
                    <RANKING order="15" place="15" resultid="17594" />
                    <RANKING order="16" place="16" resultid="17599" />
                    <RANKING order="17" place="17" resultid="18125" />
                    <RANKING order="18" place="18" resultid="17927" />
                    <RANKING order="19" place="-1" resultid="18393" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1162" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18060" />
                    <RANKING order="2" place="2" resultid="17113" />
                    <RANKING order="3" place="3" resultid="17261" />
                    <RANKING order="4" place="4" resultid="17058" />
                    <RANKING order="5" place="5" resultid="18212" />
                    <RANKING order="6" place="6" resultid="17274" />
                    <RANKING order="7" place="7" resultid="18197" />
                    <RANKING order="8" place="8" resultid="17489" />
                    <RANKING order="9" place="9" resultid="17312" />
                    <RANKING order="10" place="10" resultid="17826" />
                    <RANKING order="11" place="11" resultid="17087" />
                    <RANKING order="12" place="12" resultid="17316" />
                    <RANKING order="13" place="13" resultid="17442" />
                    <RANKING order="14" place="14" resultid="18432" />
                    <RANKING order="15" place="15" resultid="17280" />
                    <RANKING order="16" place="16" resultid="16912" />
                    <RANKING order="17" place="17" resultid="18182" />
                    <RANKING order="18" place="18" resultid="17127" />
                    <RANKING order="19" place="19" resultid="16918" />
                    <RANKING order="20" place="20" resultid="16923" />
                    <RANKING order="21" place="21" resultid="17041" />
                    <RANKING order="22" place="22" resultid="17706" />
                    <RANKING order="23" place="23" resultid="16933" />
                    <RANKING order="24" place="24" resultid="17961" />
                    <RANKING order="25" place="25" resultid="17164" />
                    <RANKING order="26" place="26" resultid="17005" />
                    <RANKING order="27" place="27" resultid="18330" />
                    <RANKING order="28" place="28" resultid="18486" />
                    <RANKING order="29" place="29" resultid="17120" />
                    <RANKING order="30" place="30" resultid="18547" />
                    <RANKING order="31" place="31" resultid="16927" />
                    <RANKING order="32" place="32" resultid="18370" />
                    <RANKING order="33" place="33" resultid="17094" />
                    <RANKING order="34" place="34" resultid="18402" />
                    <RANKING order="35" place="35" resultid="17081" />
                    <RANKING order="36" place="36" resultid="17322" />
                    <RANKING order="37" place="37" resultid="17604" />
                    <RANKING order="38" place="38" resultid="17146" />
                    <RANKING order="39" place="39" resultid="18398" />
                    <RANKING order="40" place="40" resultid="17611" />
                    <RANKING order="41" place="41" resultid="17170" />
                    <RANKING order="42" place="42" resultid="17328" />
                    <RANKING order="43" place="43" resultid="18119" />
                    <RANKING order="44" place="44" resultid="18593" />
                    <RANKING order="45" place="45" resultid="17594" />
                    <RANKING order="46" place="46" resultid="17599" />
                    <RANKING order="47" place="47" resultid="18345" />
                    <RANKING order="48" place="48" resultid="18351" />
                    <RANKING order="49" place="49" resultid="18105" />
                    <RANKING order="50" place="50" resultid="18125" />
                    <RANKING order="51" place="51" resultid="17157" />
                    <RANKING order="52" place="52" resultid="17947" />
                    <RANKING order="53" place="53" resultid="18112" />
                    <RANKING order="54" place="54" resultid="17617" />
                    <RANKING order="55" place="55" resultid="17927" />
                    <RANKING order="56" place="56" resultid="17934" />
                    <RANKING order="57" place="57" resultid="18131" />
                    <RANKING order="58" place="-1" resultid="18204" />
                    <RANKING order="59" place="-1" resultid="18393" />
                    <RANKING order="60" place="-1" resultid="18480" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19060" daytime="15:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19061" daytime="15:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19062" daytime="15:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19063" daytime="15:52" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19064" daytime="15:54" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19065" daytime="15:56" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19066" daytime="15:58" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1163" daytime="15:59" gender="M" number="28" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1164" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18227" />
                    <RANKING order="2" place="2" resultid="17869" />
                    <RANKING order="3" place="3" resultid="17239" />
                    <RANKING order="4" place="4" resultid="17890" />
                    <RANKING order="5" place="5" resultid="17883" />
                    <RANKING order="6" place="6" resultid="17418" />
                    <RANKING order="7" place="7" resultid="16962" />
                    <RANKING order="8" place="8" resultid="17557" />
                    <RANKING order="9" place="9" resultid="17806" />
                    <RANKING order="10" place="10" resultid="18608" />
                    <RANKING order="11" place="11" resultid="18034" />
                    <RANKING order="12" place="12" resultid="17206" />
                    <RANKING order="13" place="13" resultid="17246" />
                    <RANKING order="14" place="14" resultid="17365" />
                    <RANKING order="15" place="15" resultid="17678" />
                    <RANKING order="16" place="16" resultid="17847" />
                    <RANKING order="17" place="17" resultid="18322" />
                    <RANKING order="18" place="18" resultid="17509" />
                    <RANKING order="19" place="19" resultid="17671" />
                    <RANKING order="20" place="20" resultid="17107" />
                    <RANKING order="21" place="21" resultid="17378" />
                    <RANKING order="22" place="22" resultid="18502" />
                    <RANKING order="23" place="23" resultid="17180" />
                    <RANKING order="24" place="24" resultid="16947" />
                    <RANKING order="25" place="25" resultid="17523" />
                    <RANKING order="26" place="26" resultid="17664" />
                    <RANKING order="27" place="27" resultid="17372" />
                    <RANKING order="28" place="28" resultid="17954" />
                    <RANKING order="29" place="29" resultid="18002" />
                    <RANKING order="30" place="30" resultid="18599" />
                    <RANKING order="31" place="31" resultid="17812" />
                    <RANKING order="32" place="32" resultid="18273" />
                    <RANKING order="33" place="33" resultid="17876" />
                    <RANKING order="34" place="34" resultid="17352" />
                    <RANKING order="35" place="35" resultid="18255" />
                    <RANKING order="36" place="36" resultid="18294" />
                    <RANKING order="37" place="37" resultid="17516" />
                    <RANKING order="38" place="38" resultid="18241" />
                    <RANKING order="39" place="39" resultid="17819" />
                    <RANKING order="40" place="40" resultid="18287" />
                    <RANKING order="41" place="41" resultid="18014" />
                    <RANKING order="42" place="42" resultid="17996" />
                    <RANKING order="43" place="43" resultid="18280" />
                    <RANKING order="44" place="-1" resultid="16967" />
                    <RANKING order="45" place="-1" resultid="17658" />
                    <RANKING order="46" place="-1" resultid="17798" />
                    <RANKING order="47" place="-1" resultid="17991" />
                    <RANKING order="48" place="-1" resultid="18248" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1165" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17645" />
                    <RANKING order="2" place="2" resultid="17232" />
                    <RANKING order="3" place="3" resultid="17186" />
                    <RANKING order="4" place="4" resultid="17840" />
                    <RANKING order="5" place="5" resultid="17740" />
                    <RANKING order="6" place="6" resultid="17638" />
                    <RANKING order="7" place="7" resultid="18266" />
                    <RANKING order="8" place="8" resultid="18315" />
                    <RANKING order="9" place="9" resultid="17219" />
                    <RANKING order="10" place="10" resultid="16980" />
                    <RANKING order="11" place="11" resultid="17552" />
                    <RANKING order="12" place="12" resultid="17855" />
                    <RANKING order="13" place="13" resultid="18047" />
                    <RANKING order="14" place="14" resultid="18092" />
                    <RANKING order="15" place="15" resultid="18427" />
                    <RANKING order="16" place="16" resultid="18552" />
                    <RANKING order="17" place="17" resultid="17063" />
                    <RANKING order="18" place="18" resultid="17685" />
                    <RANKING order="19" place="19" resultid="17019" />
                    <RANKING order="20" place="20" resultid="18234" />
                    <RANKING order="21" place="21" resultid="17791" />
                    <RANKING order="22" place="22" resultid="18009" />
                    <RANKING order="23" place="23" resultid="18020" />
                    <RANKING order="24" place="24" resultid="18557" />
                    <RANKING order="25" place="25" resultid="18508" />
                    <RANKING order="26" place="26" resultid="18172" />
                    <RANKING order="27" place="27" resultid="18562" />
                    <RANKING order="28" place="28" resultid="17986" />
                    <RANKING order="29" place="29" resultid="17199" />
                    <RANKING order="30" place="-1" resultid="17253" />
                    <RANKING order="31" place="-1" resultid="18357" />
                    <RANKING order="32" place="-1" resultid="18525" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1166" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17226" />
                    <RANKING order="2" place="2" resultid="17384" />
                    <RANKING order="3" place="3" resultid="17346" />
                    <RANKING order="4" place="4" resultid="17495" />
                    <RANKING order="5" place="5" resultid="17212" />
                    <RANKING order="6" place="6" resultid="17340" />
                    <RANKING order="7" place="7" resultid="17391" />
                    <RANKING order="8" place="8" resultid="17424" />
                    <RANKING order="9" place="9" resultid="17402" />
                    <RANKING order="10" place="10" resultid="17645" />
                    <RANKING order="11" place="11" resultid="18259" />
                    <RANKING order="12" place="12" resultid="18137" />
                    <RANKING order="13" place="13" resultid="16973" />
                    <RANKING order="14" place="14" resultid="17232" />
                    <RANKING order="15" place="15" resultid="17192" />
                    <RANKING order="16" place="16" resultid="17542" />
                    <RANKING order="17" place="17" resultid="17186" />
                    <RANKING order="18" place="18" resultid="17466" />
                    <RANKING order="19" place="19" resultid="17015" />
                    <RANKING order="20" place="20" resultid="17840" />
                    <RANKING order="21" place="21" resultid="17397" />
                    <RANKING order="22" place="22" resultid="17740" />
                    <RANKING order="23" place="23" resultid="16988" />
                    <RANKING order="24" place="24" resultid="17638" />
                    <RANKING order="25" place="25" resultid="18266" />
                    <RANKING order="26" place="26" resultid="18227" />
                    <RANKING order="27" place="27" resultid="18315" />
                    <RANKING order="28" place="28" resultid="17219" />
                    <RANKING order="29" place="29" resultid="16980" />
                    <RANKING order="30" place="30" resultid="17552" />
                    <RANKING order="31" place="31" resultid="17869" />
                    <RANKING order="32" place="32" resultid="17239" />
                    <RANKING order="33" place="33" resultid="17855" />
                    <RANKING order="34" place="34" resultid="18047" />
                    <RANKING order="35" place="35" resultid="18092" />
                    <RANKING order="36" place="36" resultid="18427" />
                    <RANKING order="37" place="37" resultid="18552" />
                    <RANKING order="38" place="38" resultid="17890" />
                    <RANKING order="39" place="39" resultid="17063" />
                    <RANKING order="40" place="40" resultid="17685" />
                    <RANKING order="41" place="41" resultid="17883" />
                    <RANKING order="42" place="42" resultid="17019" />
                    <RANKING order="43" place="43" resultid="18234" />
                    <RANKING order="44" place="44" resultid="17791" />
                    <RANKING order="45" place="45" resultid="17418" />
                    <RANKING order="46" place="46" resultid="16962" />
                    <RANKING order="47" place="47" resultid="17531" />
                    <RANKING order="48" place="48" resultid="17557" />
                    <RANKING order="49" place="49" resultid="18009" />
                    <RANKING order="50" place="50" resultid="17806" />
                    <RANKING order="51" place="51" resultid="18020" />
                    <RANKING order="52" place="52" resultid="18608" />
                    <RANKING order="53" place="53" resultid="18557" />
                    <RANKING order="54" place="54" resultid="18508" />
                    <RANKING order="55" place="55" resultid="18034" />
                    <RANKING order="56" place="56" resultid="17206" />
                    <RANKING order="57" place="57" resultid="18172" />
                    <RANKING order="58" place="58" resultid="17246" />
                    <RANKING order="59" place="59" resultid="18562" />
                    <RANKING order="60" place="60" resultid="17365" />
                    <RANKING order="61" place="61" resultid="17678" />
                    <RANKING order="62" place="62" resultid="17847" />
                    <RANKING order="63" place="63" resultid="18322" />
                    <RANKING order="64" place="64" resultid="17509" />
                    <RANKING order="65" place="65" resultid="17671" />
                    <RANKING order="66" place="66" resultid="17107" />
                    <RANKING order="67" place="67" resultid="17378" />
                    <RANKING order="68" place="68" resultid="18502" />
                    <RANKING order="69" place="69" resultid="17180" />
                    <RANKING order="70" place="70" resultid="16947" />
                    <RANKING order="71" place="71" resultid="17523" />
                    <RANKING order="72" place="72" resultid="17664" />
                    <RANKING order="73" place="73" resultid="17372" />
                    <RANKING order="74" place="74" resultid="17954" />
                    <RANKING order="75" place="75" resultid="17986" />
                    <RANKING order="76" place="76" resultid="18002" />
                    <RANKING order="77" place="77" resultid="17199" />
                    <RANKING order="78" place="78" resultid="18599" />
                    <RANKING order="79" place="79" resultid="17812" />
                    <RANKING order="80" place="80" resultid="18273" />
                    <RANKING order="81" place="81" resultid="17876" />
                    <RANKING order="82" place="82" resultid="17352" />
                    <RANKING order="83" place="83" resultid="18255" />
                    <RANKING order="84" place="84" resultid="18294" />
                    <RANKING order="85" place="85" resultid="17516" />
                    <RANKING order="86" place="86" resultid="18241" />
                    <RANKING order="87" place="87" resultid="17819" />
                    <RANKING order="88" place="88" resultid="18287" />
                    <RANKING order="89" place="89" resultid="18014" />
                    <RANKING order="90" place="90" resultid="17996" />
                    <RANKING order="91" place="91" resultid="18280" />
                    <RANKING order="92" place="-1" resultid="16967" />
                    <RANKING order="93" place="-1" resultid="16887" />
                    <RANKING order="94" place="-1" resultid="17253" />
                    <RANKING order="95" place="-1" resultid="17628" />
                    <RANKING order="96" place="-1" resultid="17658" />
                    <RANKING order="97" place="-1" resultid="17798" />
                    <RANKING order="98" place="-1" resultid="17991" />
                    <RANKING order="99" place="-1" resultid="18248" />
                    <RANKING order="100" place="-1" resultid="18357" />
                    <RANKING order="101" place="-1" resultid="18525" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19067" daytime="15:59" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19068" daytime="16:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19069" daytime="16:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19070" daytime="16:07" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19071" daytime="16:09" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19072" daytime="16:11" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19073" daytime="16:13" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19074" daytime="16:14" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="19075" daytime="16:16" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="19076" daytime="16:18" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="19077" daytime="16:19" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1167" daytime="16:27" gender="F" number="29" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1168" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17070" />
                    <RANKING order="2" place="2" resultid="18183" />
                    <RANKING order="3" place="3" resultid="16913" />
                    <RANKING order="4" place="4" resultid="18040" />
                    <RANKING order="5" place="5" resultid="16919" />
                    <RANKING order="6" place="6" resultid="18189" />
                    <RANKING order="7" place="7" resultid="17100" />
                    <RANKING order="8" place="8" resultid="17746" />
                    <RANKING order="9" place="9" resultid="17713" />
                    <RANKING order="10" place="10" resultid="18028" />
                    <RANKING order="11" place="11" resultid="17733" />
                    <RANKING order="12" place="12" resultid="18403" />
                    <RANKING order="13" place="13" resultid="17147" />
                    <RANKING order="14" place="14" resultid="17605" />
                    <RANKING order="15" place="15" resultid="18106" />
                    <RANKING order="16" place="16" resultid="18113" />
                    <RANKING order="17" place="17" resultid="18346" />
                    <RANKING order="18" place="18" resultid="17948" />
                    <RANKING order="19" place="19" resultid="17618" />
                    <RANKING order="20" place="20" resultid="17935" />
                    <RANKING order="21" place="-1" resultid="17692" />
                    <RANKING order="22" place="-1" resultid="18205" />
                    <RANKING order="23" place="-1" resultid="18481" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1169" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17030" />
                    <RANKING order="2" place="2" resultid="18433" />
                    <RANKING order="3" place="3" resultid="17770" />
                    <RANKING order="4" place="4" resultid="18055" />
                    <RANKING order="5" place="5" resultid="17046" />
                    <RANKING order="6" place="6" resultid="18571" />
                    <RANKING order="7" place="7" resultid="18541" />
                    <RANKING order="8" place="8" resultid="18308" />
                    <RANKING order="9" place="9" resultid="17928" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1170" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17287" />
                    <RANKING order="2" place="2" resultid="18219" />
                    <RANKING order="3" place="3" resultid="17267" />
                    <RANKING order="4" place="4" resultid="17294" />
                    <RANKING order="5" place="5" resultid="17030" />
                    <RANKING order="6" place="6" resultid="17911" />
                    <RANKING order="7" place="7" resultid="17070" />
                    <RANKING order="8" place="8" resultid="18183" />
                    <RANKING order="9" place="9" resultid="18433" />
                    <RANKING order="10" place="10" resultid="17300" />
                    <RANKING order="11" place="11" resultid="18213" />
                    <RANKING order="12" place="12" resultid="17770" />
                    <RANKING order="13" place="13" resultid="18055" />
                    <RANKING order="14" place="14" resultid="17501" />
                    <RANKING order="15" place="15" resultid="17046" />
                    <RANKING order="16" place="16" resultid="18571" />
                    <RANKING order="17" place="17" resultid="16928" />
                    <RANKING order="18" place="18" resultid="16913" />
                    <RANKING order="19" place="19" resultid="18040" />
                    <RANKING order="20" place="20" resultid="18541" />
                    <RANKING order="21" place="21" resultid="16919" />
                    <RANKING order="22" place="22" resultid="18189" />
                    <RANKING order="23" place="23" resultid="17100" />
                    <RANKING order="24" place="24" resultid="17746" />
                    <RANKING order="25" place="25" resultid="17713" />
                    <RANKING order="26" place="26" resultid="18028" />
                    <RANKING order="27" place="27" resultid="17733" />
                    <RANKING order="28" place="28" resultid="18403" />
                    <RANKING order="29" place="29" resultid="18308" />
                    <RANKING order="30" place="30" resultid="17147" />
                    <RANKING order="31" place="31" resultid="17174" />
                    <RANKING order="32" place="32" resultid="17605" />
                    <RANKING order="33" place="33" resultid="18106" />
                    <RANKING order="34" place="34" resultid="18113" />
                    <RANKING order="35" place="35" resultid="18346" />
                    <RANKING order="36" place="36" resultid="17948" />
                    <RANKING order="37" place="37" resultid="17618" />
                    <RANKING order="38" place="38" resultid="17935" />
                    <RANKING order="39" place="39" resultid="17928" />
                    <RANKING order="40" place="-1" resultid="17692" />
                    <RANKING order="41" place="-1" resultid="18205" />
                    <RANKING order="42" place="-1" resultid="18481" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19078" daytime="16:27" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19079" daytime="16:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19080" daytime="16:32" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19081" daytime="16:34" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19082" daytime="16:36" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1171" daytime="16:38" gender="M" number="30" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1172" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18228" />
                    <RANKING order="2" place="2" resultid="17870" />
                    <RANKING order="3" place="3" resultid="17891" />
                    <RANKING order="4" place="4" resultid="17752" />
                    <RANKING order="5" place="5" resultid="17884" />
                    <RANKING order="6" place="6" resultid="17240" />
                    <RANKING order="7" place="7" resultid="17140" />
                    <RANKING order="8" place="8" resultid="17726" />
                    <RANKING order="9" place="9" resultid="17181" />
                    <RANKING order="10" place="10" resultid="17679" />
                    <RANKING order="11" place="11" resultid="16948" />
                    <RANKING order="12" place="12" resultid="17247" />
                    <RANKING order="13" place="13" resultid="18600" />
                    <RANKING order="14" place="14" resultid="18256" />
                    <RANKING order="15" place="15" resultid="17665" />
                    <RANKING order="16" place="16" resultid="18003" />
                    <RANKING order="17" place="17" resultid="17877" />
                    <RANKING order="18" place="18" resultid="18274" />
                    <RANKING order="19" place="19" resultid="18295" />
                    <RANKING order="20" place="20" resultid="17517" />
                    <RANKING order="21" place="21" resultid="17672" />
                    <RANKING order="22" place="22" resultid="17820" />
                    <RANKING order="23" place="23" resultid="17813" />
                    <RANKING order="24" place="24" resultid="18242" />
                    <RANKING order="25" place="25" resultid="18288" />
                    <RANKING order="26" place="-1" resultid="17153" />
                    <RANKING order="27" place="-1" resultid="17510" />
                    <RANKING order="28" place="-1" resultid="17848" />
                    <RANKING order="29" place="-1" resultid="18249" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1173" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17906" />
                    <RANKING order="2" place="2" resultid="17254" />
                    <RANKING order="3" place="3" resultid="17833" />
                    <RANKING order="4" place="4" resultid="18442" />
                    <RANKING order="5" place="5" resultid="17233" />
                    <RANKING order="6" place="6" resultid="17863" />
                    <RANKING order="7" place="7" resultid="17562" />
                    <RANKING order="8" place="8" resultid="17220" />
                    <RANKING order="9" place="9" resultid="18509" />
                    <RANKING order="10" place="10" resultid="18021" />
                    <RANKING order="11" place="11" resultid="17686" />
                    <RANKING order="12" place="12" resultid="18173" />
                    <RANKING order="13" place="-1" resultid="17200" />
                    <RANKING order="14" place="-1" resultid="17639" />
                    <RANKING order="15" place="-1" resultid="18358" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1174" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17476" />
                    <RANKING order="2" place="2" resultid="17906" />
                    <RANKING order="3" place="3" resultid="17429" />
                    <RANKING order="4" place="4" resultid="18438" />
                    <RANKING order="5" place="5" resultid="17898" />
                    <RANKING order="6" place="6" resultid="17193" />
                    <RANKING order="7" place="7" resultid="17254" />
                    <RANKING order="8" place="8" resultid="16974" />
                    <RANKING order="9" place="9" resultid="17833" />
                    <RANKING order="10" place="10" resultid="18442" />
                    <RANKING order="11" place="11" resultid="17233" />
                    <RANKING order="12" place="12" resultid="18260" />
                    <RANKING order="13" place="13" resultid="18228" />
                    <RANKING order="14" place="14" resultid="17870" />
                    <RANKING order="15" place="15" resultid="17623" />
                    <RANKING order="16" place="16" resultid="17863" />
                    <RANKING order="17" place="17" resultid="17891" />
                    <RANKING order="18" place="18" resultid="17537" />
                    <RANKING order="19" place="19" resultid="17752" />
                    <RANKING order="20" place="20" resultid="17562" />
                    <RANKING order="21" place="21" resultid="17654" />
                    <RANKING order="22" place="22" resultid="17884" />
                    <RANKING order="23" place="23" resultid="17220" />
                    <RANKING order="24" place="24" resultid="18509" />
                    <RANKING order="25" place="25" resultid="17240" />
                    <RANKING order="26" place="26" resultid="18021" />
                    <RANKING order="27" place="27" resultid="17140" />
                    <RANKING order="28" place="28" resultid="17686" />
                    <RANKING order="29" place="29" resultid="17726" />
                    <RANKING order="30" place="30" resultid="17181" />
                    <RANKING order="31" place="31" resultid="17679" />
                    <RANKING order="32" place="32" resultid="18173" />
                    <RANKING order="33" place="33" resultid="16948" />
                    <RANKING order="34" place="34" resultid="17247" />
                    <RANKING order="35" place="35" resultid="18600" />
                    <RANKING order="36" place="36" resultid="18256" />
                    <RANKING order="37" place="37" resultid="17665" />
                    <RANKING order="38" place="38" resultid="18003" />
                    <RANKING order="39" place="39" resultid="17877" />
                    <RANKING order="40" place="40" resultid="18274" />
                    <RANKING order="41" place="41" resultid="18295" />
                    <RANKING order="42" place="42" resultid="17517" />
                    <RANKING order="43" place="43" resultid="17672" />
                    <RANKING order="44" place="44" resultid="17820" />
                    <RANKING order="45" place="45" resultid="17813" />
                    <RANKING order="46" place="46" resultid="18242" />
                    <RANKING order="47" place="47" resultid="18288" />
                    <RANKING order="48" place="-1" resultid="17153" />
                    <RANKING order="49" place="-1" resultid="17200" />
                    <RANKING order="50" place="-1" resultid="17510" />
                    <RANKING order="51" place="-1" resultid="17581" />
                    <RANKING order="52" place="-1" resultid="17639" />
                    <RANKING order="53" place="-1" resultid="17848" />
                    <RANKING order="54" place="-1" resultid="18249" />
                    <RANKING order="55" place="-1" resultid="18358" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19083" daytime="16:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19084" daytime="16:41" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19085" daytime="16:44" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19086" daytime="16:46" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19087" daytime="16:48" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19088" daytime="16:50" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1175" daytime="16:58" gender="F" number="31" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1176" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16993" />
                    <RANKING order="2" place="2" resultid="16999" />
                    <RANKING order="3" place="3" resultid="18190" />
                    <RANKING order="4" place="4" resultid="17693" />
                    <RANKING order="5" place="5" resultid="17714" />
                    <RANKING order="6" place="6" resultid="19110" />
                    <RANKING order="7" place="7" resultid="17161" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1177" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17114" />
                    <RANKING order="2" place="2" resultid="17827" />
                    <RANKING order="3" place="3" resultid="17707" />
                    <RANKING order="4" place="4" resultid="17075" />
                    <RANKING order="5" place="5" resultid="17128" />
                    <RANKING order="6" place="6" resultid="18301" />
                    <RANKING order="7" place="7" resultid="18309" />
                    <RANKING order="8" place="8" resultid="18126" />
                    <RANKING order="9" place="-1" resultid="17088" />
                    <RANKING order="10" place="-1" resultid="17699" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1178" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17411" />
                    <RANKING order="2" place="2" resultid="18337" />
                    <RANKING order="3" place="3" resultid="17114" />
                    <RANKING order="4" place="4" resultid="17827" />
                    <RANKING order="5" place="5" resultid="17707" />
                    <RANKING order="6" place="6" resultid="17075" />
                    <RANKING order="7" place="7" resultid="17128" />
                    <RANKING order="8" place="8" resultid="16993" />
                    <RANKING order="9" place="9" resultid="18301" />
                    <RANKING order="10" place="10" resultid="16999" />
                    <RANKING order="11" place="11" resultid="17121" />
                    <RANKING order="12" place="12" resultid="18190" />
                    <RANKING order="13" place="13" resultid="17693" />
                    <RANKING order="14" place="14" resultid="17714" />
                    <RANKING order="15" place="15" resultid="18309" />
                    <RANKING order="16" place="16" resultid="19110" />
                    <RANKING order="17" place="17" resultid="18126" />
                    <RANKING order="18" place="18" resultid="17161" />
                    <RANKING order="19" place="-1" resultid="17088" />
                    <RANKING order="20" place="-1" resultid="17699" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19089" daytime="16:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19090" daytime="17:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19091" daytime="17:06" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1179" daytime="17:10" gender="M" number="32" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1180" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17849" />
                    <RANKING order="2" place="2" resultid="17134" />
                    <RANKING order="3" place="3" resultid="17753" />
                    <RANKING order="4" place="4" resultid="17727" />
                    <RANKING order="5" place="5" resultid="18616" />
                    <RANKING order="6" place="6" resultid="17955" />
                    <RANKING order="7" place="7" resultid="17799" />
                    <RANKING order="8" place="8" resultid="17366" />
                    <RANKING order="9" place="9" resultid="18376" />
                    <RANKING order="10" place="10" resultid="17524" />
                    <RANKING order="11" place="11" resultid="18323" />
                    <RANKING order="12" place="12" resultid="18612" />
                    <RANKING order="13" place="13" resultid="17353" />
                    <RANKING order="14" place="14" resultid="18281" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1181" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17834" />
                    <RANKING order="2" place="2" resultid="17646" />
                    <RANKING order="3" place="3" resultid="18073" />
                    <RANKING order="4" place="4" resultid="17570" />
                    <RANKING order="5" place="5" resultid="17792" />
                    <RANKING order="6" place="6" resultid="18413" />
                    <RANKING order="7" place="7" resultid="18235" />
                    <RANKING order="8" place="-1" resultid="17841" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1182" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17435" />
                    <RANKING order="2" place="2" resultid="17425" />
                    <RANKING order="3" place="3" resultid="17024" />
                    <RANKING order="4" place="4" resultid="17834" />
                    <RANKING order="5" place="5" resultid="17646" />
                    <RANKING order="6" place="6" resultid="18138" />
                    <RANKING order="7" place="7" resultid="18073" />
                    <RANKING order="8" place="8" resultid="17570" />
                    <RANKING order="9" place="9" resultid="17849" />
                    <RANKING order="10" place="10" resultid="17792" />
                    <RANKING order="11" place="11" resultid="17134" />
                    <RANKING order="12" place="12" resultid="18413" />
                    <RANKING order="13" place="13" resultid="17753" />
                    <RANKING order="14" place="14" resultid="17727" />
                    <RANKING order="15" place="15" resultid="18616" />
                    <RANKING order="16" place="16" resultid="17955" />
                    <RANKING order="17" place="17" resultid="18235" />
                    <RANKING order="18" place="18" resultid="17799" />
                    <RANKING order="19" place="19" resultid="17366" />
                    <RANKING order="20" place="20" resultid="18376" />
                    <RANKING order="21" place="21" resultid="17524" />
                    <RANKING order="22" place="22" resultid="18323" />
                    <RANKING order="23" place="23" resultid="18612" />
                    <RANKING order="24" place="24" resultid="17353" />
                    <RANKING order="25" place="25" resultid="18281" />
                    <RANKING order="26" place="-1" resultid="17841" />
                    <RANKING order="27" place="-1" resultid="18944" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19092" daytime="17:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19093" daytime="17:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19094" daytime="17:19" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1183" daytime="17:23" gender="F" number="33" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1184" agemax="13" agemin="12" name="MŁODZIK">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17000" />
                    <RANKING order="2" place="2" resultid="18487" />
                    <RANKING order="3" place="3" resultid="17734" />
                    <RANKING order="4" place="4" resultid="18041" />
                    <RANKING order="5" place="5" resultid="17720" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1185" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18061" />
                    <RANKING order="2" place="2" resultid="17771" />
                    <RANKING order="3" place="3" resultid="18542" />
                    <RANKING order="4" place="4" resultid="18079" />
                    <RANKING order="5" place="5" resultid="17047" />
                    <RANKING order="6" place="6" resultid="18302" />
                    <RANKING order="7" place="-1" resultid="17700" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1186" agemax="-1" agemin="12" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18338" />
                    <RANKING order="2" place="2" resultid="17262" />
                    <RANKING order="3" place="3" resultid="17490" />
                    <RANKING order="4" place="4" resultid="17313" />
                    <RANKING order="5" place="5" resultid="17268" />
                    <RANKING order="6" place="6" resultid="18198" />
                    <RANKING order="7" place="7" resultid="17275" />
                    <RANKING order="8" place="8" resultid="17449" />
                    <RANKING order="9" place="9" resultid="18061" />
                    <RANKING order="10" place="10" resultid="17912" />
                    <RANKING order="11" place="11" resultid="18220" />
                    <RANKING order="12" place="12" resultid="17771" />
                    <RANKING order="13" place="13" resultid="17288" />
                    <RANKING order="14" place="14" resultid="17281" />
                    <RANKING order="15" place="15" resultid="18542" />
                    <RANKING order="16" place="16" resultid="17412" />
                    <RANKING order="17" place="17" resultid="17000" />
                    <RANKING order="18" place="18" resultid="18079" />
                    <RANKING order="19" place="19" resultid="18487" />
                    <RANKING order="20" place="20" resultid="17734" />
                    <RANKING order="21" place="21" resultid="18041" />
                    <RANKING order="22" place="22" resultid="17047" />
                    <RANKING order="23" place="23" resultid="18302" />
                    <RANKING order="24" place="24" resultid="17720" />
                    <RANKING order="25" place="-1" resultid="17700" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19095" daytime="17:23" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19096" daytime="17:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19097" daytime="17:47" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1191" daytime="17:58" gender="M" number="34" order="23" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1194" agemax="15" agemin="14" name="JUNIOR MŁODSZY">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17064" />
                    <RANKING order="2" place="2" resultid="18086" />
                    <RANKING order="3" place="3" resultid="17856" />
                    <RANKING order="4" place="4" resultid="18316" />
                    <RANKING order="5" place="5" resultid="18267" />
                    <RANKING order="6" place="6" resultid="18093" />
                    <RANKING order="7" place="7" resultid="17053" />
                    <RANKING order="8" place="8" resultid="18048" />
                    <RANKING order="9" place="-1" resultid="17741" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6371" agemax="-1" agemin="14" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17496" />
                    <RANKING order="2" place="2" resultid="17064" />
                    <RANKING order="3" place="3" resultid="18086" />
                    <RANKING order="4" place="4" resultid="17856" />
                    <RANKING order="5" place="5" resultid="18316" />
                    <RANKING order="6" place="6" resultid="18267" />
                    <RANKING order="7" place="7" resultid="18093" />
                    <RANKING order="8" place="8" resultid="17053" />
                    <RANKING order="9" place="9" resultid="18048" />
                    <RANKING order="10" place="-1" resultid="17741" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19099" daytime="17:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19100" daytime="18:19" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="01603" nation="POL" region="03" clubid="18139" name="UKS &quot;Piątka&quot;">
          <ATHLETES>
            <ATHLETE firstname="Igor" lastname="Kozak" birthdate="2008-02-29" gender="M" nation="POL" license="101603700010" swrid="5109152" athleteid="18158">
              <RESULTS>
                <RESULT eventid="1063" points="246" reactiontime="+77" swimtime="00:00:33.37" resultid="18159" heatid="18957" lane="8" entrytime="00:00:34.10" entrycourse="LCM" />
                <RESULT eventid="1087" status="DNS" swimtime="00:00:00.00" resultid="18160" heatid="18988" lane="4" entrytime="00:02:49.08" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Tworkowski" birthdate="2008-03-17" gender="M" nation="POL" license="101603700003" swrid="5109148" athleteid="18146">
              <RESULTS>
                <RESULT eventid="1063" points="345" reactiontime="+70" swimtime="00:00:29.80" resultid="18147" heatid="18959" lane="6" entrytime="00:00:30.44" entrycourse="LCM" />
                <RESULT eventid="1071" points="393" reactiontime="+54" swimtime="00:00:35.40" resultid="18148" heatid="18974" lane="9" entrytime="00:00:34.92" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonina" lastname="Szabała" birthdate="2009-06-04" gender="F" nation="POL" license="101603600002" swrid="5112631" athleteid="18177">
              <RESULTS>
                <RESULT eventid="1075" points="498" reactiontime="+70" swimtime="00:01:09.96" resultid="18178" heatid="18977" lane="1" entrytime="00:01:08.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1091" points="496" reactiontime="+75" swimtime="00:02:35.82" resultid="18179" heatid="18992" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.14" />
                    <SPLIT distance="100" swimtime="00:01:17.73" />
                    <SPLIT distance="150" swimtime="00:01:57.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="533" reactiontime="+54" swimtime="00:00:30.13" resultid="18180" heatid="19017" lane="2" entrytime="00:00:29.79" entrycourse="LCM" />
                <RESULT comment="G2 - Pływak zanurzył się całkowicie w trakcie wyścigu (z wyjątkiem 15 m po starcie lub nawrocie)" eventid="1117" reactiontime="+72" status="DSQ" swimtime="00:00:33.32" resultid="18181" heatid="19026" lane="7" />
                <RESULT eventid="1159" points="503" reactiontime="+73" swimtime="00:01:05.00" resultid="18182" heatid="19065" lane="0" entrytime="00:01:06.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="544" reactiontime="+76" swimtime="00:01:10.50" resultid="18183" heatid="19081" lane="2" entrytime="00:01:12.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Miazio" birthdate="2008-04-20" gender="M" nation="POL" license="101603700012" swrid="5331607" athleteid="18152">
              <RESULTS>
                <RESULT eventid="1063" points="307" reactiontime="+52" swimtime="00:00:30.97" resultid="18153" heatid="18959" lane="2" entrytime="00:00:30.47" entrycourse="LCM" />
                <RESULT comment="K14 - Pływak wykonał kopnięcie nóg w płaszczyźnie pionowej w dół (z wyjątkiem jednego ruchu po starcie lub nawrocie)" eventid="1071" reactiontime="+75" status="DSQ" swimtime="00:00:43.03" resultid="18154" heatid="18972" lane="7" entrytime="00:00:40.84" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maksymilian" lastname="Woliński" birthdate="2007-04-19" gender="M" nation="POL" license="101603700029" swrid="5455438" athleteid="18167">
              <RESULTS>
                <RESULT eventid="1063" points="233" reactiontime="+88" swimtime="00:00:33.98" resultid="18168" heatid="18957" lane="9" entrytime="00:00:34.26" entrycourse="LCM" />
                <RESULT eventid="1087" points="264" reactiontime="+85" swimtime="00:02:38.84" resultid="18169" heatid="18987" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="159" reactiontime="+91" swimtime="00:00:41.05" resultid="18170" heatid="19019" lane="3" />
                <RESULT eventid="1121" points="197" reactiontime="+77" swimtime="00:00:41.24" resultid="18171" heatid="19035" lane="8" entrytime="00:00:41.16" entrycourse="LCM" />
                <RESULT eventid="1163" points="263" reactiontime="+88" swimtime="00:01:13.15" resultid="18172" heatid="19071" lane="1" entrytime="00:01:15.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="192" reactiontime="+66" swimtime="00:01:29.73" resultid="18173" heatid="19085" lane="3" entrytime="00:01:30.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrian" lastname="Sternik" birthdate="2008-06-04" gender="M" nation="POL" license="101603700008" swrid="5164074" athleteid="18164">
              <RESULTS>
                <RESULT eventid="1063" status="DNS" swimtime="00:00:00.00" resultid="18165" heatid="18958" lane="4" entrytime="00:00:31.24" entrycourse="LCM" />
                <RESULT eventid="1087" status="DNS" swimtime="00:00:00.00" resultid="18166" heatid="18989" lane="2" entrytime="00:02:37.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Łachowski" birthdate="2008-12-02" gender="M" nation="POL" license="101603700005" swrid="5173029" athleteid="18155">
              <RESULTS>
                <RESULT eventid="1063" status="DNS" swimtime="00:00:00.00" resultid="18156" heatid="18952" lane="6" />
                <RESULT eventid="1087" status="DNS" swimtime="00:00:00.00" resultid="18157" heatid="18989" lane="6" entrytime="00:02:35.69" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kaja" lastname="Kostyła" birthdate="2009-11-28" gender="F" nation="POL" license="101603600006" swrid="5173249" athleteid="18184">
              <RESULTS>
                <RESULT eventid="1091" points="366" reactiontime="+58" swimtime="00:02:52.36" resultid="18185" heatid="18993" lane="7" entrytime="00:02:56.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.36" />
                    <SPLIT distance="100" swimtime="00:01:26.65" />
                    <SPLIT distance="150" swimtime="00:02:11.24" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G8 - Pływak ukończył wyścig w położeniu na piersiach" eventid="1099" status="DSQ" swimtime="00:06:02.54" resultid="18186" heatid="18998" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.06" />
                    <SPLIT distance="100" swimtime="00:01:26.31" />
                    <SPLIT distance="150" swimtime="00:02:13.21" />
                    <SPLIT distance="200" swimtime="00:02:58.13" />
                    <SPLIT distance="250" swimtime="00:03:50.99" />
                    <SPLIT distance="300" swimtime="00:04:41.29" />
                    <SPLIT distance="350" swimtime="00:05:22.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="325" swimtime="00:01:33.26" resultid="18187" heatid="19039" lane="5" entrytime="00:01:44.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="376" reactiontime="+67" swimtime="00:02:54.67" resultid="18188" heatid="19048" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.27" />
                    <SPLIT distance="100" swimtime="00:01:22.97" />
                    <SPLIT distance="150" swimtime="00:02:15.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="375" reactiontime="+63" swimtime="00:01:19.79" resultid="18189" heatid="19081" lane="9" entrytime="00:01:21.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="353" swimtime="00:03:16.80" resultid="18190" heatid="19090" lane="7" entrytime="00:03:30.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.98" />
                    <SPLIT distance="100" swimtime="00:01:38.11" />
                    <SPLIT distance="150" swimtime="00:02:28.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Złomańczuk" birthdate="2008-06-08" gender="M" nation="POL" license="101603700004" swrid="5173036" athleteid="18149">
              <RESULTS>
                <RESULT eventid="1063" points="369" reactiontime="+73" swimtime="00:00:29.13" resultid="18150" heatid="18960" lane="9" entrytime="00:00:29.46" entrycourse="LCM" />
                <RESULT eventid="1087" points="374" reactiontime="+80" swimtime="00:02:21.50" resultid="18151" heatid="18990" lane="0" entrytime="00:02:23.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                    <SPLIT distance="100" swimtime="00:01:09.73" />
                    <SPLIT distance="150" swimtime="00:01:46.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Kostyła" birthdate="2008-04-24" gender="M" nation="POL" license="101603700009" swrid="5173254" athleteid="18161">
              <RESULTS>
                <RESULT eventid="1063" points="274" reactiontime="+62" swimtime="00:00:32.18" resultid="18162" heatid="18957" lane="4" entrytime="00:00:32.68" entrycourse="LCM" />
                <RESULT eventid="1071" points="175" reactiontime="+50" swimtime="00:00:46.34" resultid="18163" heatid="18971" lane="8" entrytime="00:00:44.91" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patryk" lastname="Joachimowicz" birthdate="2008-06-07" gender="M" nation="POL" license="101603700011" swrid="5109163" athleteid="18174">
              <RESULTS>
                <RESULT eventid="1071" points="391" reactiontime="+63" swimtime="00:00:35.48" resultid="18175" heatid="18973" lane="9" entrytime="00:00:38.24" entrycourse="LCM" />
                <RESULT eventid="1103" points="482" reactiontime="+75" swimtime="00:05:10.92" resultid="18176" heatid="19000" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                    <SPLIT distance="100" swimtime="00:01:08.49" />
                    <SPLIT distance="150" swimtime="00:01:49.46" />
                    <SPLIT distance="200" swimtime="00:02:30.08" />
                    <SPLIT distance="250" swimtime="00:03:14.22" />
                    <SPLIT distance="300" swimtime="00:03:59.27" />
                    <SPLIT distance="350" swimtime="00:04:35.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Szpak" birthdate="2008-07-26" gender="F" nation="POL" license="101603600026" swrid="5455437" athleteid="18143">
              <RESULTS>
                <RESULT eventid="1059" points="248" reactiontime="+88" swimtime="00:00:37.67" resultid="18144" heatid="18947" lane="7" entrytime="00:00:37.62" entrycourse="LCM" />
                <RESULT eventid="1067" points="210" swimtime="00:00:49.45" resultid="18145" heatid="18965" lane="2" entrytime="00:00:48.83" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michalina" lastname="Szkoda" birthdate="2008-02-16" gender="F" nation="POL" license="101603600032" swrid="5331606" athleteid="18140">
              <RESULTS>
                <RESULT eventid="1059" points="394" reactiontime="+65" swimtime="00:00:32.28" resultid="18141" heatid="18948" lane="4" entrytime="00:00:31.85" entrycourse="LCM" />
                <RESULT eventid="1083" points="398" reactiontime="+75" swimtime="00:02:33.58" resultid="18142" heatid="18983" lane="1" entrytime="00:02:34.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                    <SPLIT distance="100" swimtime="00:01:16.30" />
                    <SPLIT distance="150" swimtime="00:01:57.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00309" nation="POL" region="09" clubid="17577" name="MKS Juvenia Białystok">
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Danilewski" birthdate="1998-10-19" gender="M" nation="POL" license="100309700396" swrid="4406045" athleteid="17578">
              <RESULTS>
                <RESULT eventid="1095" status="DNS" swimtime="00:00:00.00" resultid="17579" heatid="18995" lane="5" />
                <RESULT eventid="1121" status="DNS" swimtime="00:00:00.00" resultid="17580" heatid="19032" lane="3" />
                <RESULT eventid="1171" reactiontime="+97" status="DNS" swimtime="00:00:00.00" resultid="17581" heatid="19084" lane="7" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00203" nation="POL" region="03" clubid="18191" name="UKS ,,ORKA&apos;&apos; Zamość">
          <ATHLETES>
            <ATHLETE firstname="Julia" lastname="Malinoś" birthdate="2004-03-09" gender="F" nation="POL" license="100203600118" swrid="4936860" athleteid="18192">
              <RESULTS>
                <RESULT eventid="1059" points="621" reactiontime="+62" swimtime="00:00:27.73" resultid="18193" heatid="18951" lane="7" entrytime="00:00:27.51" entrycourse="LCM" />
                <RESULT eventid="1083" points="564" reactiontime="+66" swimtime="00:02:16.74" resultid="18194" heatid="18984" lane="4" entrytime="00:02:14.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                    <SPLIT distance="100" swimtime="00:01:06.78" />
                    <SPLIT distance="150" swimtime="00:01:42.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="537" reactiontime="+63" swimtime="00:04:50.83" resultid="18195" heatid="19007" lane="8" entrytime="00:04:42.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                    <SPLIT distance="100" swimtime="00:01:07.84" />
                    <SPLIT distance="150" swimtime="00:01:45.22" />
                    <SPLIT distance="200" swimtime="00:02:22.19" />
                    <SPLIT distance="250" swimtime="00:02:59.81" />
                    <SPLIT distance="300" swimtime="00:03:37.16" />
                    <SPLIT distance="350" swimtime="00:04:14.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6361" points="565" reactiontime="+64" swimtime="00:18:32.95" resultid="18196" heatid="19055" lane="4" entrytime="00:18:48.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                    <SPLIT distance="100" swimtime="00:01:08.24" />
                    <SPLIT distance="150" swimtime="00:01:44.88" />
                    <SPLIT distance="200" swimtime="00:02:21.41" />
                    <SPLIT distance="250" swimtime="00:02:58.20" />
                    <SPLIT distance="300" swimtime="00:03:35.07" />
                    <SPLIT distance="350" swimtime="00:04:12.52" />
                    <SPLIT distance="400" swimtime="00:04:49.54" />
                    <SPLIT distance="450" swimtime="00:05:26.93" />
                    <SPLIT distance="500" swimtime="00:06:04.25" />
                    <SPLIT distance="550" swimtime="00:06:41.95" />
                    <SPLIT distance="600" swimtime="00:07:19.34" />
                    <SPLIT distance="650" swimtime="00:07:57.20" />
                    <SPLIT distance="700" swimtime="00:08:34.53" />
                    <SPLIT distance="750" swimtime="00:09:11.95" />
                    <SPLIT distance="800" swimtime="00:09:49.21" />
                    <SPLIT distance="850" swimtime="00:10:26.97" />
                    <SPLIT distance="900" swimtime="00:11:04.27" />
                    <SPLIT distance="950" swimtime="00:11:41.81" />
                    <SPLIT distance="1000" swimtime="00:12:19.18" />
                    <SPLIT distance="1050" swimtime="00:12:56.79" />
                    <SPLIT distance="1100" swimtime="00:13:34.19" />
                    <SPLIT distance="1150" swimtime="00:14:12.06" />
                    <SPLIT distance="1200" swimtime="00:14:49.73" />
                    <SPLIT distance="1250" swimtime="00:15:27.49" />
                    <SPLIT distance="1300" swimtime="00:16:04.71" />
                    <SPLIT distance="1350" swimtime="00:16:42.45" />
                    <SPLIT distance="1400" swimtime="00:17:19.83" />
                    <SPLIT distance="1450" swimtime="00:17:57.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="554" reactiontime="+66" swimtime="00:01:02.95" resultid="18197" heatid="19066" lane="1" entrytime="00:01:01.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="564" reactiontime="+68" swimtime="00:09:46.45" resultid="18198" heatid="19097" lane="6" entrytime="00:09:42.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                    <SPLIT distance="100" swimtime="00:01:08.41" />
                    <SPLIT distance="150" swimtime="00:01:44.81" />
                    <SPLIT distance="200" swimtime="00:02:21.52" />
                    <SPLIT distance="250" swimtime="00:02:58.12" />
                    <SPLIT distance="300" swimtime="00:03:35.04" />
                    <SPLIT distance="350" swimtime="00:04:12.16" />
                    <SPLIT distance="400" swimtime="00:04:49.57" />
                    <SPLIT distance="450" swimtime="00:05:26.99" />
                    <SPLIT distance="500" swimtime="00:06:04.41" />
                    <SPLIT distance="550" swimtime="00:06:41.72" />
                    <SPLIT distance="600" swimtime="00:07:19.12" />
                    <SPLIT distance="650" swimtime="00:07:56.06" />
                    <SPLIT distance="700" swimtime="00:08:33.40" />
                    <SPLIT distance="750" swimtime="00:09:10.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Sioma" birthdate="2004-10-04" gender="F" nation="POL" license="100203600144" swrid="5032671" athleteid="18214">
              <RESULTS>
                <RESULT eventid="1059" points="579" reactiontime="+73" swimtime="00:00:28.39" resultid="18215" heatid="18946" lane="7" />
                <RESULT eventid="1091" points="590" reactiontime="+64" swimtime="00:02:27.03" resultid="18216" heatid="18994" lane="3" entrytime="00:02:26.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                    <SPLIT distance="100" swimtime="00:01:11.69" />
                    <SPLIT distance="150" swimtime="00:01:50.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="647" reactiontime="+67" swimtime="00:00:31.18" resultid="18217" heatid="19030" lane="5" entrytime="00:00:31.21" entrycourse="LCM" />
                <RESULT eventid="1141" points="569" reactiontime="+74" swimtime="00:02:32.15" resultid="18218" heatid="19050" lane="6" entrytime="00:02:28.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                    <SPLIT distance="100" swimtime="00:01:10.48" />
                    <SPLIT distance="150" swimtime="00:01:55.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="606" reactiontime="+71" swimtime="00:01:08.02" resultid="18219" heatid="19082" lane="5" entrytime="00:01:06.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="514" reactiontime="+75" swimtime="00:10:04.88" resultid="18220" heatid="19097" lane="7" entrytime="00:10:03.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                    <SPLIT distance="100" swimtime="00:01:08.99" />
                    <SPLIT distance="150" swimtime="00:01:45.76" />
                    <SPLIT distance="200" swimtime="00:02:23.38" />
                    <SPLIT distance="250" swimtime="00:03:01.64" />
                    <SPLIT distance="300" swimtime="00:03:39.77" />
                    <SPLIT distance="350" swimtime="00:04:19.06" />
                    <SPLIT distance="400" swimtime="00:04:57.48" />
                    <SPLIT distance="450" swimtime="00:05:36.17" />
                    <SPLIT distance="500" swimtime="00:06:14.75" />
                    <SPLIT distance="550" swimtime="00:06:53.22" />
                    <SPLIT distance="600" swimtime="00:07:32.55" />
                    <SPLIT distance="650" swimtime="00:08:11.18" />
                    <SPLIT distance="700" swimtime="00:08:49.86" />
                    <SPLIT distance="750" swimtime="00:09:28.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Bondyra" birthdate="2009-07-31" gender="M" nation="POL" license="100203700253" swrid="4889159" athleteid="18317">
              <RESULTS>
                <RESULT eventid="1071" points="194" reactiontime="+79" swimtime="00:00:44.81" resultid="18318" heatid="18971" lane="2" entrytime="00:00:44.07" entrycourse="LCM" />
                <RESULT eventid="1103" points="214" reactiontime="+58" swimtime="00:06:47.12" resultid="18319" heatid="19001" lane="9" entrytime="00:07:09.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.02" />
                    <SPLIT distance="100" swimtime="00:01:41.18" />
                    <SPLIT distance="150" swimtime="00:02:34.13" />
                    <SPLIT distance="200" swimtime="00:03:22.96" />
                    <SPLIT distance="250" swimtime="00:04:19.50" />
                    <SPLIT distance="300" swimtime="00:05:14.85" />
                    <SPLIT distance="350" swimtime="00:06:02.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1137" points="191" swimtime="00:01:38.68" resultid="18320" heatid="19044" lane="5" entrytime="00:01:39.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="198" swimtime="00:03:15.56" resultid="18321" heatid="19053" lane="9" entrytime="00:03:10.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.00" />
                    <SPLIT distance="100" swimtime="00:01:36.30" />
                    <SPLIT distance="150" swimtime="00:02:33.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="241" swimtime="00:01:15.30" resultid="18322" heatid="19069" lane="5" entrytime="00:01:23.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="185" swimtime="00:03:41.06" resultid="18323" heatid="19093" lane="9" entrytime="00:03:29.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.76" />
                    <SPLIT distance="100" swimtime="00:01:47.14" />
                    <SPLIT distance="150" swimtime="00:02:44.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Kowalczuk" birthdate="2008-07-25" gender="M" nation="POL" license="100203700271" swrid="5455433" athleteid="18243">
              <RESULTS>
                <RESULT eventid="1063" status="DNS" swimtime="00:00:00.00" resultid="18244" heatid="18954" lane="3" entrytime="00:00:42.56" entrycourse="LCM" />
                <RESULT eventid="1095" status="DNS" swimtime="00:00:00.00" resultid="18245" heatid="18996" lane="2" entrytime="00:03:51.06" entrycourse="LCM" />
                <RESULT eventid="1121" status="DNS" swimtime="00:00:00.00" resultid="18246" heatid="19034" lane="8" entrytime="00:00:48.45" entrycourse="LCM" />
                <RESULT eventid="1137" status="DNS" swimtime="00:00:00.00" resultid="18247" heatid="19043" lane="7" />
                <RESULT eventid="1163" status="DNS" swimtime="00:00:00.00" resultid="18248" heatid="19068" lane="1" entrytime="00:01:52.82" entrycourse="LCM" />
                <RESULT eventid="1171" status="DNS" swimtime="00:00:00.00" resultid="18249" heatid="19084" lane="4" entrytime="00:01:46.49" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patrycja" lastname="Stadnik" birthdate="2009-07-05" gender="F" nation="POL" license="100203600289" swrid="5455133" athleteid="18199">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="18200" heatid="18946" lane="4" entrytime="00:00:41.28" entrycourse="LCM" />
                <RESULT eventid="1083" status="DNS" swimtime="00:00:00.00" resultid="18201" heatid="18982" lane="3" entrytime="00:03:14.98" entrycourse="LCM" />
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="18202" heatid="19015" lane="9" entrytime="00:00:45.25" entrycourse="LCM" />
                <RESULT eventid="1117" status="DNS" swimtime="00:00:00.00" resultid="18203" heatid="19027" lane="0" entrytime="00:00:51.12" entrycourse="LCM" />
                <RESULT eventid="1159" status="DNS" swimtime="00:00:00.00" resultid="18204" heatid="19061" lane="4" entrytime="00:01:27.66" entrycourse="LCM" />
                <RESULT eventid="1167" status="DNS" swimtime="00:00:00.00" resultid="18205" heatid="19079" lane="2" entrytime="00:01:58.23" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Bigos" birthdate="2008-11-27" gender="M" nation="POL" license="100203700254" swrid="5393765" athleteid="18268">
              <RESULTS>
                <RESULT eventid="1063" points="169" reactiontime="+91" swimtime="00:00:37.77" resultid="18269" heatid="18956" lane="0" entrytime="00:00:37.39" entrycourse="LCM" />
                <RESULT eventid="1087" points="150" reactiontime="+94" swimtime="00:03:11.81" resultid="18270" heatid="18988" lane="0" entrytime="00:03:13.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.81" />
                    <SPLIT distance="150" swimtime="00:02:24.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="154" reactiontime="+92" swimtime="00:06:50.28" resultid="18271" heatid="19009" lane="4" entrytime="00:06:45.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.91" />
                    <SPLIT distance="100" swimtime="00:01:32.75" />
                    <SPLIT distance="150" swimtime="00:02:27.10" />
                    <SPLIT distance="200" swimtime="00:03:19.55" />
                    <SPLIT distance="250" swimtime="00:04:13.38" />
                    <SPLIT distance="300" swimtime="00:05:06.90" />
                    <SPLIT distance="350" swimtime="00:06:00.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="142" reactiontime="+78" swimtime="00:00:45.95" resultid="18272" heatid="19034" lane="2" entrytime="00:00:45.56" entrycourse="LCM" />
                <RESULT eventid="1163" points="146" reactiontime="+85" swimtime="00:01:28.97" resultid="18273" heatid="19069" lane="6" entrytime="00:01:24.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="128" reactiontime="+83" swimtime="00:01:42.79" resultid="18274" heatid="19085" lane="1" entrytime="00:01:41.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nina" lastname="Leszkowicz" birthdate="2007-05-24" gender="F" nation="POL" license="100203600200" swrid="5219473" athleteid="18303">
              <RESULTS>
                <RESULT eventid="1067" points="310" reactiontime="+68" swimtime="00:00:43.44" resultid="18304" heatid="18966" lane="1" entrytime="00:00:40.91" entrycourse="LCM" />
                <RESULT eventid="1091" points="267" reactiontime="+68" swimtime="00:03:11.50" resultid="18305" heatid="18993" lane="1" entrytime="00:03:03.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.85" />
                    <SPLIT distance="100" swimtime="00:01:32.07" />
                    <SPLIT distance="150" swimtime="00:02:22.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="310" reactiontime="+58" swimtime="00:00:39.84" resultid="18306" heatid="19028" lane="8" entrytime="00:00:39.94" entrycourse="LCM" />
                <RESULT eventid="1133" points="319" reactiontime="+66" swimtime="00:01:33.81" resultid="18307" heatid="19040" lane="7" entrytime="00:01:31.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="292" reactiontime="+66" swimtime="00:01:26.71" resultid="18308" heatid="19080" lane="8" entrytime="00:01:27.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="311" reactiontime="+73" swimtime="00:03:25.11" resultid="18309" heatid="19090" lane="6" entrytime="00:03:20.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.08" />
                    <SPLIT distance="100" swimtime="00:01:37.11" />
                    <SPLIT distance="150" swimtime="00:02:31.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Kropornicki" birthdate="2006-01-10" gender="M" nation="POL" license="100203700204" swrid="5244408" athleteid="18261">
              <RESULTS>
                <RESULT eventid="1063" points="492" reactiontime="+55" swimtime="00:00:26.48" resultid="18262" heatid="18961" lane="2" entrytime="00:00:26.72" entrycourse="LCM" />
                <RESULT eventid="1079" points="379" reactiontime="+64" swimtime="00:01:08.37" resultid="18263" heatid="18980" lane="7" entrytime="00:01:08.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="450" reactiontime="+65" swimtime="00:00:29.05" resultid="18264" heatid="19023" lane="4" entrytime="00:00:29.59" entrycourse="LCM" />
                <RESULT eventid="1145" points="372" reactiontime="+67" swimtime="00:02:38.38" resultid="18265" heatid="19052" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                    <SPLIT distance="100" swimtime="00:01:14.36" />
                    <SPLIT distance="150" swimtime="00:02:02.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="475" reactiontime="+60" swimtime="00:01:00.11" resultid="18266" heatid="19075" lane="9" entrytime="00:01:00.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="461" reactiontime="+64" swimtime="00:18:47.40" resultid="18267" heatid="19099" lane="4" entrytime="00:19:22.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                    <SPLIT distance="100" swimtime="00:01:08.21" />
                    <SPLIT distance="150" swimtime="00:01:45.40" />
                    <SPLIT distance="200" swimtime="00:02:22.88" />
                    <SPLIT distance="250" swimtime="00:03:00.64" />
                    <SPLIT distance="300" swimtime="00:03:37.83" />
                    <SPLIT distance="350" swimtime="00:04:15.42" />
                    <SPLIT distance="400" swimtime="00:04:53.21" />
                    <SPLIT distance="450" swimtime="00:05:29.95" />
                    <SPLIT distance="500" swimtime="00:06:06.78" />
                    <SPLIT distance="550" swimtime="00:06:43.50" />
                    <SPLIT distance="600" swimtime="00:07:20.06" />
                    <SPLIT distance="650" swimtime="00:07:57.53" />
                    <SPLIT distance="700" swimtime="00:08:34.49" />
                    <SPLIT distance="750" swimtime="00:09:12.21" />
                    <SPLIT distance="800" swimtime="00:09:49.59" />
                    <SPLIT distance="850" swimtime="00:10:26.62" />
                    <SPLIT distance="900" swimtime="00:11:04.03" />
                    <SPLIT distance="950" swimtime="00:11:41.68" />
                    <SPLIT distance="1000" swimtime="00:12:20.13" />
                    <SPLIT distance="1050" swimtime="00:12:58.54" />
                    <SPLIT distance="1100" swimtime="00:13:37.52" />
                    <SPLIT distance="1150" swimtime="00:14:16.76" />
                    <SPLIT distance="1200" swimtime="00:14:56.02" />
                    <SPLIT distance="1250" swimtime="00:15:35.65" />
                    <SPLIT distance="1300" swimtime="00:16:15.05" />
                    <SPLIT distance="1350" swimtime="00:16:55.01" />
                    <SPLIT distance="1400" swimtime="00:17:34.00" />
                    <SPLIT distance="1450" swimtime="00:18:12.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alan" lastname="Mazur" birthdate="2009-11-22" gender="M" nation="POL" license="100203700247" swrid="5141018" athleteid="18282">
              <RESULTS>
                <RESULT eventid="1063" points="110" reactiontime="+96" swimtime="00:00:43.62" resultid="18283" heatid="18954" lane="5" entrytime="00:00:41.86" entrycourse="LCM" />
                <RESULT eventid="1071" points="79" reactiontime="+94" swimtime="00:01:00.47" resultid="18284" heatid="18969" lane="3" />
                <RESULT eventid="1113" points="77" swimtime="00:00:52.33" resultid="18285" heatid="19020" lane="8" />
                <RESULT eventid="1145" points="100" reactiontime="+99" swimtime="00:04:05.21" resultid="18286" heatid="19051" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.63" />
                    <SPLIT distance="100" swimtime="00:01:55.82" />
                    <SPLIT distance="150" swimtime="00:03:11.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="104" reactiontime="+93" swimtime="00:01:39.72" resultid="18287" heatid="19068" lane="6" entrytime="00:01:37.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="88" reactiontime="+98" swimtime="00:01:56.50" resultid="18288" heatid="19083" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Szuper" birthdate="2004-08-17" gender="F" nation="POL" license="100203600150" swrid="4892174" athleteid="18206">
              <RESULTS>
                <RESULT eventid="1059" points="603" reactiontime="+64" swimtime="00:00:28.01" resultid="18207" heatid="18951" lane="1" entrytime="00:00:28.09" entrycourse="LCM" />
                <RESULT eventid="1083" points="617" reactiontime="+65" swimtime="00:02:12.66" resultid="18208" heatid="18985" lane="8" entrytime="00:02:13.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                    <SPLIT distance="100" swimtime="00:01:04.62" />
                    <SPLIT distance="150" swimtime="00:01:38.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="514" reactiontime="+64" swimtime="00:00:30.48" resultid="18209" heatid="19017" lane="6" entrytime="00:00:29.75" entrycourse="LCM" />
                <RESULT eventid="1117" points="604" reactiontime="+71" swimtime="00:00:31.90" resultid="18210" heatid="19030" lane="2" entrytime="00:00:31.57" entrycourse="LCM" />
                <RESULT eventid="1141" status="DNS" swimtime="00:00:00.00" resultid="18211" heatid="19048" lane="8" />
                <RESULT eventid="1159" points="579" reactiontime="+67" swimtime="00:01:02.04" resultid="18212" heatid="19066" lane="7" entrytime="00:01:01.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="504" reactiontime="+73" swimtime="00:01:12.32" resultid="18213" heatid="19082" lane="7" entrytime="00:01:08.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Wołoszyn" birthdate="2009-12-26" gender="M" nation="POL" license="100203700240" swrid="5140943" athleteid="18289">
              <RESULTS>
                <RESULT eventid="1063" points="144" reactiontime="+77" swimtime="00:00:39.86" resultid="18290" heatid="18955" lane="1" entrytime="00:00:39.78" entrycourse="LCM" />
                <RESULT eventid="1079" points="55" reactiontime="+79" swimtime="00:02:09.61" resultid="18291" heatid="18979" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="134" reactiontime="+60" swimtime="00:07:09.38" resultid="18292" heatid="19009" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.16" />
                    <SPLIT distance="100" swimtime="00:01:35.29" />
                    <SPLIT distance="150" swimtime="00:02:30.44" />
                    <SPLIT distance="200" swimtime="00:03:25.96" />
                    <SPLIT distance="250" swimtime="00:04:23.78" />
                    <SPLIT distance="300" swimtime="00:05:21.00" />
                    <SPLIT distance="350" swimtime="00:06:15.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="129" reactiontime="+72" swimtime="00:00:47.40" resultid="18293" heatid="19033" lane="4" entrytime="00:00:49.05" entrycourse="LCM" />
                <RESULT eventid="1163" points="130" reactiontime="+68" swimtime="00:01:32.37" resultid="18294" heatid="19068" lane="5" entrytime="00:01:32.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="124" reactiontime="+71" swimtime="00:01:43.88" resultid="18295" heatid="19084" lane="6" entrytime="00:01:52.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Franczuk" birthdate="2009-09-12" gender="M" nation="POL" license="100203700264" swrid="5448196" athleteid="18275">
              <RESULTS>
                <RESULT eventid="1063" points="99" reactiontime="+51" swimtime="00:00:45.19" resultid="18276" heatid="18952" lane="8" />
                <RESULT eventid="1071" points="119" swimtime="00:00:52.67" resultid="18277" heatid="18970" lane="8" entrytime="00:00:52.09" entrycourse="LCM" />
                <RESULT eventid="1137" points="107" swimtime="00:01:59.75" resultid="18278" heatid="19044" lane="0" entrytime="00:01:57.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="106" swimtime="00:04:00.52" resultid="18279" heatid="19052" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.30" />
                    <SPLIT distance="100" swimtime="00:02:01.69" />
                    <SPLIT distance="150" swimtime="00:03:03.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="85" swimtime="00:01:46.32" resultid="18280" heatid="19068" lane="7" entrytime="00:01:47.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="122" reactiontime="+77" swimtime="00:04:14.20" resultid="18281" heatid="19092" lane="6" entrytime="00:04:05.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.85" />
                    <SPLIT distance="100" swimtime="00:02:04.29" />
                    <SPLIT distance="150" swimtime="00:03:08.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Bednarz" birthdate="2004-08-02" gender="F" nation="POL" license="100203600115" swrid="5032660" athleteid="18331">
              <RESULTS>
                <RESULT eventid="1083" points="634" reactiontime="+77" swimtime="00:02:11.51" resultid="18332" heatid="18985" lane="3" entrytime="00:02:11.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.10" />
                    <SPLIT distance="100" swimtime="00:01:04.50" />
                    <SPLIT distance="150" swimtime="00:01:38.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="651" reactiontime="+81" swimtime="00:05:07.29" resultid="18333" heatid="18999" lane="4" entrytime="00:05:06.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                    <SPLIT distance="100" swimtime="00:01:10.53" />
                    <SPLIT distance="150" swimtime="00:01:51.40" />
                    <SPLIT distance="200" swimtime="00:02:31.08" />
                    <SPLIT distance="250" swimtime="00:03:12.67" />
                    <SPLIT distance="300" swimtime="00:03:55.33" />
                    <SPLIT distance="350" swimtime="00:04:32.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="634" reactiontime="+81" swimtime="00:04:35.19" resultid="18334" heatid="19007" lane="3" entrytime="00:04:35.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                    <SPLIT distance="100" swimtime="00:01:06.38" />
                    <SPLIT distance="150" swimtime="00:01:41.28" />
                    <SPLIT distance="200" swimtime="00:02:16.14" />
                    <SPLIT distance="250" swimtime="00:02:51.03" />
                    <SPLIT distance="300" swimtime="00:03:26.15" />
                    <SPLIT distance="350" swimtime="00:04:00.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" status="DNS" swimtime="00:00:00.00" resultid="18335" heatid="19041" lane="3" entrytime="00:01:17.59" entrycourse="LCM" />
                <RESULT eventid="1141" points="649" reactiontime="+81" swimtime="00:02:25.61" resultid="18336" heatid="19050" lane="3" entrytime="00:02:25.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.16" />
                    <SPLIT distance="100" swimtime="00:01:10.79" />
                    <SPLIT distance="150" swimtime="00:01:52.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="621" reactiontime="+82" swimtime="00:02:42.98" resultid="18337" heatid="19091" lane="4" entrytime="00:02:40.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                    <SPLIT distance="100" swimtime="00:01:19.50" />
                    <SPLIT distance="150" swimtime="00:02:01.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="605" reactiontime="+86" swimtime="00:09:33.18" resultid="18338" heatid="19097" lane="3" entrytime="00:09:36.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.14" />
                    <SPLIT distance="100" swimtime="00:01:08.52" />
                    <SPLIT distance="150" swimtime="00:01:44.63" />
                    <SPLIT distance="200" swimtime="00:02:20.93" />
                    <SPLIT distance="250" swimtime="00:02:57.11" />
                    <SPLIT distance="300" swimtime="00:03:33.29" />
                    <SPLIT distance="350" swimtime="00:04:09.54" />
                    <SPLIT distance="400" swimtime="00:04:45.93" />
                    <SPLIT distance="450" swimtime="00:05:22.31" />
                    <SPLIT distance="500" swimtime="00:05:58.45" />
                    <SPLIT distance="550" swimtime="00:06:35.03" />
                    <SPLIT distance="600" swimtime="00:07:11.05" />
                    <SPLIT distance="650" swimtime="00:07:46.65" />
                    <SPLIT distance="700" swimtime="00:08:22.66" />
                    <SPLIT distance="750" swimtime="00:08:58.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Duda" birthdate="2008-09-01" gender="M" nation="POL" license="100203700276" swrid="5455431" athleteid="18236">
              <RESULTS>
                <RESULT eventid="1063" points="131" swimtime="00:00:41.07" resultid="18237" heatid="18955" lane="2" entrytime="00:00:39.41" entrycourse="LCM" />
                <RESULT eventid="1087" status="DNS" swimtime="00:00:00.00" resultid="18238" heatid="18987" lane="5" entrytime="00:03:29.87" entrycourse="LCM" />
                <RESULT eventid="1113" points="62" reactiontime="+80" swimtime="00:00:55.98" resultid="18239" heatid="19020" lane="4" entrytime="00:00:58.35" entrycourse="LCM" />
                <RESULT eventid="1121" points="99" reactiontime="+77" swimtime="00:00:51.81" resultid="18240" heatid="19033" lane="2" entrytime="00:00:53.07" entrycourse="LCM" />
                <RESULT eventid="1163" points="120" reactiontime="+86" swimtime="00:01:35.00" resultid="18241" heatid="19068" lane="3" entrytime="00:01:36.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="99" reactiontime="+76" swimtime="00:01:52.03" resultid="18242" heatid="19084" lane="2" entrytime="00:02:00.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabela" lastname="Naklicka" birthdate="2006-11-14" gender="F" nation="POL" license="100203600188" swrid="4901073" athleteid="18324">
              <RESULTS>
                <RESULT eventid="1075" points="490" reactiontime="+70" swimtime="00:01:10.34" resultid="18325" heatid="18977" lane="9" entrytime="00:01:11.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="403" reactiontime="+76" swimtime="00:02:32.94" resultid="18326" heatid="18984" lane="1" entrytime="00:02:25.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.17" />
                    <SPLIT distance="100" swimtime="00:01:14.53" />
                    <SPLIT distance="150" swimtime="00:01:54.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="457" swimtime="00:00:31.70" resultid="18327" heatid="19017" lane="9" entrytime="00:00:31.60" entrycourse="LCM" />
                <RESULT eventid="1141" points="412" reactiontime="+74" swimtime="00:02:49.39" resultid="18328" heatid="19048" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.49" />
                    <SPLIT distance="100" swimtime="00:01:18.36" />
                    <SPLIT distance="150" swimtime="00:02:09.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1150" points="364" reactiontime="+73" swimtime="00:02:50.59" resultid="18329" heatid="19057" lane="8" entrytime="00:02:50.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.56" />
                    <SPLIT distance="100" swimtime="00:01:23.60" />
                    <SPLIT distance="150" swimtime="00:02:09.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="428" reactiontime="+71" swimtime="00:01:08.57" resultid="18330" heatid="19065" lane="9" entrytime="00:01:06.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Charkot" birthdate="2008-01-07" gender="M" nation="POL" license="100203700206" swrid="5219465" athleteid="18221">
              <RESULTS>
                <RESULT eventid="1063" points="456" reactiontime="+69" swimtime="00:00:27.15" resultid="18222" heatid="18961" lane="8" entrytime="00:00:26.96" entrycourse="LCM" />
                <RESULT eventid="1087" points="489" reactiontime="+74" swimtime="00:02:09.43" resultid="18223" heatid="18990" lane="3" entrytime="00:02:14.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.54" />
                    <SPLIT distance="100" swimtime="00:01:04.22" />
                    <SPLIT distance="150" swimtime="00:01:38.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="486" reactiontime="+74" swimtime="00:04:39.75" resultid="18224" heatid="19009" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.77" />
                    <SPLIT distance="100" swimtime="00:01:07.31" />
                    <SPLIT distance="150" swimtime="00:01:43.35" />
                    <SPLIT distance="200" swimtime="00:02:18.95" />
                    <SPLIT distance="250" swimtime="00:02:56.68" />
                    <SPLIT distance="300" swimtime="00:03:32.14" />
                    <SPLIT distance="350" swimtime="00:04:07.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="404" reactiontime="+78" swimtime="00:00:30.12" resultid="18225" heatid="19023" lane="6" entrytime="00:00:30.11" entrycourse="LCM" />
                <RESULT eventid="1163" points="470" reactiontime="+77" swimtime="00:01:00.30" resultid="18227" heatid="19075" lane="0" entrytime="00:01:00.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="393" reactiontime="+91" swimtime="00:01:10.78" resultid="18228" heatid="19087" lane="2" entrytime="00:01:12.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kasjana" lastname="Wyłupek" birthdate="2007-03-27" gender="F" nation="POL" license="100203600225" swrid="4968998" athleteid="18296">
              <RESULTS>
                <RESULT eventid="1067" points="408" reactiontime="+65" swimtime="00:00:39.62" resultid="18297" heatid="18966" lane="6" entrytime="00:00:38.67" entrycourse="LCM" />
                <RESULT eventid="1099" reactiontime="+48" status="DNF" swimtime="00:00:00.00" resultid="18298" heatid="18999" lane="8" entrytime="00:06:02.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.06" />
                    <SPLIT distance="100" swimtime="00:01:31.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="392" reactiontime="+68" swimtime="00:01:27.62" resultid="18299" heatid="19040" lane="3" entrytime="00:01:24.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="370" reactiontime="+71" swimtime="00:02:55.58" resultid="18300" heatid="19049" lane="6" entrytime="00:02:52.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.40" />
                    <SPLIT distance="100" swimtime="00:01:24.53" />
                    <SPLIT distance="150" swimtime="00:02:12.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="409" reactiontime="+69" swimtime="00:03:07.38" resultid="18301" heatid="19091" lane="1" entrytime="00:02:56.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.33" />
                    <SPLIT distance="100" swimtime="00:01:30.29" />
                    <SPLIT distance="150" swimtime="00:02:19.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="338" reactiontime="+72" swimtime="00:11:35.54" resultid="18302" heatid="19096" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.71" />
                    <SPLIT distance="100" swimtime="00:01:20.66" />
                    <SPLIT distance="150" swimtime="00:02:04.49" />
                    <SPLIT distance="200" swimtime="00:02:48.94" />
                    <SPLIT distance="250" swimtime="00:03:32.56" />
                    <SPLIT distance="300" swimtime="00:04:16.52" />
                    <SPLIT distance="350" swimtime="00:05:00.96" />
                    <SPLIT distance="400" swimtime="00:05:44.74" />
                    <SPLIT distance="450" swimtime="00:06:30.03" />
                    <SPLIT distance="500" swimtime="00:07:13.74" />
                    <SPLIT distance="550" swimtime="00:07:58.21" />
                    <SPLIT distance="600" swimtime="00:08:42.12" />
                    <SPLIT distance="650" swimtime="00:09:26.66" />
                    <SPLIT distance="700" swimtime="00:10:09.94" />
                    <SPLIT distance="750" swimtime="00:10:53.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Chyrchała" birthdate="2002-11-19" gender="M" nation="POL" license="100203700147" swrid="4751340" athleteid="18257">
              <RESULTS>
                <RESULT eventid="1063" points="509" reactiontime="+70" swimtime="00:00:26.18" resultid="18258" heatid="18954" lane="9" />
                <RESULT eventid="1163" points="549" reactiontime="+74" swimtime="00:00:57.27" resultid="18259" heatid="19067" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="394" reactiontime="+67" swimtime="00:01:10.67" resultid="18260" heatid="19084" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="450" reactiontime="+75" status="EXH" swimtime="00:00:29.04" resultid="19111" heatid="19018" lane="6" late="yes" />
                <RESULT eventid="1121" points="436" reactiontime="+66" status="EXH" swimtime="00:00:31.65" resultid="19112" heatid="19031" lane="7" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olaf" lastname="Lupa" birthdate="2006-02-15" gender="M" nation="POL" license="100203700135" swrid="5165791" athleteid="18310">
              <RESULTS>
                <RESULT eventid="1071" points="361" reactiontime="+87" swimtime="00:00:36.44" resultid="18311" heatid="18973" lane="6" entrytime="00:00:36.14" entrycourse="LCM" />
                <RESULT eventid="1087" points="468" reactiontime="+86" swimtime="00:02:11.35" resultid="18312" heatid="18990" lane="5" entrytime="00:02:13.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                    <SPLIT distance="100" swimtime="00:01:03.74" />
                    <SPLIT distance="150" swimtime="00:01:38.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="470" reactiontime="+90" swimtime="00:04:42.98" resultid="18313" heatid="19010" lane="4" entrytime="00:04:43.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                    <SPLIT distance="100" swimtime="00:01:06.73" />
                    <SPLIT distance="150" swimtime="00:01:43.16" />
                    <SPLIT distance="200" swimtime="00:02:20.07" />
                    <SPLIT distance="250" swimtime="00:02:56.63" />
                    <SPLIT distance="300" swimtime="00:03:32.97" />
                    <SPLIT distance="350" swimtime="00:04:09.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1137" points="295" reactiontime="+91" swimtime="00:01:25.39" resultid="18314" heatid="19046" lane="4" entrytime="00:01:19.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="469" reactiontime="+92" swimtime="00:01:00.37" resultid="18315" heatid="19074" lane="5" entrytime="00:01:00.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="482" reactiontime="+90" swimtime="00:18:30.60" resultid="18316" heatid="19100" lane="9" entrytime="00:18:39.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                    <SPLIT distance="100" swimtime="00:01:09.94" />
                    <SPLIT distance="150" swimtime="00:01:47.49" />
                    <SPLIT distance="200" swimtime="00:02:24.45" />
                    <SPLIT distance="250" swimtime="00:03:01.17" />
                    <SPLIT distance="300" swimtime="00:03:39.01" />
                    <SPLIT distance="350" swimtime="00:04:16.87" />
                    <SPLIT distance="400" swimtime="00:04:54.17" />
                    <SPLIT distance="450" swimtime="00:05:32.20" />
                    <SPLIT distance="500" swimtime="00:06:10.14" />
                    <SPLIT distance="550" swimtime="00:06:48.04" />
                    <SPLIT distance="600" swimtime="00:07:25.38" />
                    <SPLIT distance="650" swimtime="00:08:03.24" />
                    <SPLIT distance="700" swimtime="00:08:40.40" />
                    <SPLIT distance="750" swimtime="00:09:18.31" />
                    <SPLIT distance="800" swimtime="00:09:56.33" />
                    <SPLIT distance="850" swimtime="00:10:33.46" />
                    <SPLIT distance="900" swimtime="00:11:10.97" />
                    <SPLIT distance="950" swimtime="00:11:49.12" />
                    <SPLIT distance="1000" swimtime="00:12:26.30" />
                    <SPLIT distance="1050" swimtime="00:13:04.18" />
                    <SPLIT distance="1100" swimtime="00:13:41.62" />
                    <SPLIT distance="1150" swimtime="00:14:19.42" />
                    <SPLIT distance="1200" swimtime="00:14:56.22" />
                    <SPLIT distance="1250" swimtime="00:15:33.53" />
                    <SPLIT distance="1300" swimtime="00:16:10.36" />
                    <SPLIT distance="1350" swimtime="00:16:46.40" />
                    <SPLIT distance="1400" swimtime="00:17:22.32" />
                    <SPLIT distance="1450" swimtime="00:17:56.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Baniak" birthdate="2007-02-02" gender="M" nation="POL" license="100203700210" swrid="5280822" athleteid="18229">
              <RESULTS>
                <RESULT eventid="1063" points="329" reactiontime="+73" swimtime="00:00:30.26" resultid="18230" heatid="18958" lane="5" entrytime="00:00:31.28" entrycourse="LCM" />
                <RESULT eventid="1087" points="310" reactiontime="+80" swimtime="00:02:30.58" resultid="18231" heatid="18989" lane="9" entrytime="00:02:44.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                    <SPLIT distance="100" swimtime="00:01:14.61" />
                    <SPLIT distance="150" swimtime="00:01:54.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="287" reactiontime="+79" swimtime="00:00:33.76" resultid="18232" heatid="19021" lane="5" entrytime="00:00:37.82" entrycourse="LCM" />
                <RESULT eventid="1137" points="226" reactiontime="+83" swimtime="00:01:33.25" resultid="18233" heatid="19044" lane="4" entrytime="00:01:39.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="340" reactiontime="+81" swimtime="00:01:07.18" resultid="18234" heatid="19071" lane="4" entrytime="00:01:13.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="229" reactiontime="+87" swimtime="00:03:25.87" resultid="18235" heatid="19092" lane="4" entrytime="00:03:38.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.67" />
                    <SPLIT distance="100" swimtime="00:01:37.30" />
                    <SPLIT distance="150" swimtime="00:02:32.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Kahan" birthdate="2009-11-05" gender="M" nation="POL" license="100203700273" swrid="5455124" athleteid="18250">
              <RESULTS>
                <RESULT eventid="1063" points="141" reactiontime="+80" swimtime="00:00:40.08" resultid="18251" heatid="18955" lane="8" entrytime="00:00:40.08" entrycourse="LCM" />
                <RESULT eventid="1087" points="129" reactiontime="+77" swimtime="00:03:21.45" resultid="18252" heatid="18988" lane="9" entrytime="00:03:18.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.60" />
                    <SPLIT distance="100" swimtime="00:01:38.47" />
                    <SPLIT distance="150" swimtime="00:02:32.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="86" swimtime="00:00:50.43" resultid="18253" heatid="19021" lane="9" entrytime="00:00:53.98" entrycourse="LCM" />
                <RESULT eventid="1121" points="150" reactiontime="+64" swimtime="00:00:45.09" resultid="18254" heatid="19034" lane="0" entrytime="00:00:48.55" entrycourse="LCM" />
                <RESULT eventid="1163" points="132" reactiontime="+79" swimtime="00:01:32.07" resultid="18255" heatid="19068" lane="4" entrytime="00:01:32.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="144" reactiontime="+73" swimtime="00:01:38.74" resultid="18256" heatid="19084" lane="3" entrytime="00:01:51.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02503" nation="POL" region="03" clubid="18474" name="UKS Olimpijczyk 23">
          <ATHLETES>
            <ATHLETE firstname="Aleksandra" lastname="Tkaczyk" birthdate="2009-04-06" gender="F" nation="POL" license="102503600140" swrid="5173034" athleteid="18475">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="18476" heatid="18948" lane="7" entrytime="00:00:34.64" entrycourse="LCM" />
                <RESULT eventid="1083" status="DNS" swimtime="00:00:00.00" resultid="18477" heatid="18982" lane="7" />
                <RESULT eventid="1125" status="DNS" swimtime="00:00:00.00" resultid="18478" heatid="19005" lane="9" />
                <RESULT eventid="1117" status="DNS" swimtime="00:00:00.00" resultid="18479" heatid="19028" lane="0" entrytime="00:00:40.28" entrycourse="LCM" />
                <RESULT eventid="1159" status="DNS" swimtime="00:00:00.00" resultid="18480" heatid="19062" lane="3" entrytime="00:01:18.18" entrycourse="LCM" />
                <RESULT eventid="1167" status="DNS" swimtime="00:00:00.00" resultid="18481" heatid="19080" lane="1" entrytime="00:01:26.46" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mikołaj" lastname="Jaskowiak" birthdate="2009-12-11" gender="M" nation="POL" license="102503700173" swrid="5440315" athleteid="18515">
              <RESULTS>
                <RESULT eventid="1063" points="107" swimtime="00:00:43.97" resultid="18516" heatid="18954" lane="2" entrytime="00:00:44.62" entrycourse="LCM" />
                <RESULT eventid="1087" points="108" reactiontime="+66" swimtime="00:03:33.98" resultid="18517" heatid="18986" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.29" />
                    <SPLIT distance="100" swimtime="00:01:44.91" />
                    <SPLIT distance="150" swimtime="00:02:40.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="52" reactiontime="+79" swimtime="00:00:59.38" resultid="18518" heatid="19020" lane="5" entrytime="00:00:59.03" entrycourse="LCM" />
                <RESULT eventid="1137" points="85" reactiontime="+59" swimtime="00:02:09.10" resultid="18519" heatid="19043" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Grabowski" birthdate="2009-08-09" gender="M" nation="POL" license="102503700139" swrid="5322105" athleteid="18531">
              <RESULTS>
                <RESULT eventid="1071" points="128" reactiontime="+72" swimtime="00:00:51.45" resultid="18532" heatid="18968" lane="3" />
                <RESULT eventid="1087" points="195" reactiontime="+63" swimtime="00:02:55.74" resultid="18533" heatid="18987" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                    <SPLIT distance="100" swimtime="00:01:26.36" />
                    <SPLIT distance="150" swimtime="00:02:14.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="220" reactiontime="+68" swimtime="00:06:04.31" resultid="18534" heatid="19010" lane="0" entrytime="00:05:56.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.73" />
                    <SPLIT distance="100" swimtime="00:01:24.99" />
                    <SPLIT distance="150" swimtime="00:02:11.07" />
                    <SPLIT distance="200" swimtime="00:02:58.60" />
                    <SPLIT distance="250" swimtime="00:03:46.82" />
                    <SPLIT distance="300" swimtime="00:04:34.53" />
                    <SPLIT distance="350" swimtime="00:05:21.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="158" reactiontime="+84" swimtime="00:00:44.39" resultid="18535" heatid="19034" lane="3" entrytime="00:00:44.86" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Pietroń" birthdate="2007-01-24" gender="M" nation="POL" license="102503700046" swrid="5019869" athleteid="18520">
              <RESULTS>
                <RESULT eventid="1087" status="DNS" swimtime="00:00:00.00" resultid="18522" heatid="18991" lane="1" entrytime="00:02:02.65" entrycourse="LCM" />
                <RESULT eventid="6365" status="DNS" swimtime="00:00:00.00" resultid="18523" heatid="19003" lane="7" entrytime="00:09:12.13" entrycourse="LCM" />
                <RESULT eventid="1129" status="DNS" swimtime="00:00:00.00" resultid="18524" heatid="19012" lane="0" entrytime="00:04:24.00" entrycourse="LCM" />
                <RESULT eventid="1163" status="DNS" swimtime="00:00:00.00" resultid="18525" heatid="19076" lane="3" entrytime="00:00:56.93" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Jasieczek" birthdate="2009-05-12" gender="M" nation="POL" license="102503700168" swrid="5440314" athleteid="18497">
              <RESULTS>
                <RESULT eventid="1063" points="234" reactiontime="+69" swimtime="00:00:33.91" resultid="18498" heatid="18956" lane="5" entrytime="00:00:34.56" entrycourse="LCM" />
                <RESULT eventid="1087" points="211" reactiontime="+70" swimtime="00:02:51.09" resultid="18499" heatid="18988" lane="2" entrytime="00:02:53.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.85" />
                    <SPLIT distance="100" swimtime="00:01:23.65" />
                    <SPLIT distance="150" swimtime="00:02:10.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="146" reactiontime="+56" swimtime="00:00:42.23" resultid="18500" heatid="19021" lane="8" entrytime="00:00:43.49" entrycourse="LCM" />
                <RESULT eventid="1145" points="197" reactiontime="+60" swimtime="00:03:15.81" resultid="18501" heatid="19052" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.32" />
                    <SPLIT distance="100" swimtime="00:01:34.21" />
                    <SPLIT distance="150" swimtime="00:02:32.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="218" reactiontime="+78" swimtime="00:01:17.85" resultid="18502" heatid="19070" lane="7" entrytime="00:01:17.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otylia" lastname="Kościołek" birthdate="2006-09-28" gender="F" nation="POL" license="102503600039" swrid="5109159" athleteid="18536">
              <RESULTS>
                <RESULT eventid="1075" points="426" reactiontime="+77" swimtime="00:01:13.73" resultid="18537" heatid="18976" lane="2" entrytime="00:01:14.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="478" reactiontime="+76" swimtime="00:05:40.47" resultid="18538" heatid="18999" lane="7" entrytime="00:05:44.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.99" />
                    <SPLIT distance="100" swimtime="00:01:15.75" />
                    <SPLIT distance="150" swimtime="00:01:58.72" />
                    <SPLIT distance="200" swimtime="00:02:41.93" />
                    <SPLIT distance="250" swimtime="00:03:31.36" />
                    <SPLIT distance="300" swimtime="00:04:20.82" />
                    <SPLIT distance="350" swimtime="00:05:01.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="393" swimtime="00:00:33.34" resultid="18539" heatid="19016" lane="2" entrytime="00:00:32.70" entrycourse="LCM" />
                <RESULT eventid="1141" points="488" reactiontime="+77" swimtime="00:02:40.09" resultid="18540" heatid="19049" lane="3" entrytime="00:02:45.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                    <SPLIT distance="100" swimtime="00:01:14.08" />
                    <SPLIT distance="150" swimtime="00:02:03.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="417" reactiontime="+80" swimtime="00:01:17.01" resultid="18541" heatid="19081" lane="8" entrytime="00:01:16.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="460" reactiontime="+74" swimtime="00:10:27.83" resultid="18542" heatid="19097" lane="9" entrytime="00:10:21.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                    <SPLIT distance="100" swimtime="00:01:09.94" />
                    <SPLIT distance="150" swimtime="00:01:48.48" />
                    <SPLIT distance="200" swimtime="00:02:27.84" />
                    <SPLIT distance="250" swimtime="00:03:07.32" />
                    <SPLIT distance="300" swimtime="00:03:47.32" />
                    <SPLIT distance="350" swimtime="00:04:27.14" />
                    <SPLIT distance="400" swimtime="00:05:07.45" />
                    <SPLIT distance="450" swimtime="00:05:47.50" />
                    <SPLIT distance="500" swimtime="00:06:28.09" />
                    <SPLIT distance="550" swimtime="00:07:07.99" />
                    <SPLIT distance="600" swimtime="00:07:48.60" />
                    <SPLIT distance="650" swimtime="00:08:28.64" />
                    <SPLIT distance="700" swimtime="00:09:08.77" />
                    <SPLIT distance="750" swimtime="00:09:48.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Kielmas" birthdate="2009-10-16" gender="M" nation="POL" license="102503700187" swrid="5453711" athleteid="18526">
              <RESULTS>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej, a przed sygnałem startu" eventid="1071" reactiontime="+46" status="DSQ" swimtime="00:00:57.53" resultid="18527" heatid="18969" lane="5" entrytime="00:00:54.47" entrycourse="LCM" />
                <RESULT eventid="1095" points="140" reactiontime="+71" swimtime="00:03:35.23" resultid="18528" heatid="18996" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.83" />
                    <SPLIT distance="100" swimtime="00:01:45.65" />
                    <SPLIT distance="150" swimtime="00:02:41.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="138" reactiontime="+55" swimtime="00:07:05.39" resultid="18529" heatid="19009" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.17" />
                    <SPLIT distance="100" swimtime="00:01:39.11" />
                    <SPLIT distance="150" swimtime="00:02:30.77" />
                    <SPLIT distance="200" swimtime="00:03:26.68" />
                    <SPLIT distance="250" swimtime="00:04:21.54" />
                    <SPLIT distance="300" swimtime="00:05:19.24" />
                    <SPLIT distance="350" swimtime="00:06:13.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="115" reactiontime="+98" swimtime="00:00:49.31" resultid="18530" heatid="19034" lane="9" entrytime="00:00:48.56" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Gałązka" birthdate="2009-06-16" gender="M" nation="POL" license="102503700155" swrid="5353675" athleteid="18510">
              <RESULTS>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej, a przed sygnałem startu" eventid="1063" status="DSQ" swimtime="00:00:38.43" resultid="18511" heatid="18956" lane="8" entrytime="00:00:37.08" entrycourse="LCM" />
                <RESULT eventid="1087" points="115" reactiontime="+67" swimtime="00:03:29.59" resultid="18512" heatid="18987" lane="3" entrytime="00:03:30.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.78" />
                    <SPLIT distance="100" swimtime="00:01:41.18" />
                    <SPLIT distance="150" swimtime="00:02:36.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="119" swimtime="00:07:26.28" resultid="18513" heatid="19009" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.06" />
                    <SPLIT distance="100" swimtime="00:01:43.02" />
                    <SPLIT distance="150" swimtime="00:02:40.91" />
                    <SPLIT distance="200" swimtime="00:03:38.15" />
                    <SPLIT distance="250" swimtime="00:04:36.17" />
                    <SPLIT distance="300" swimtime="00:05:35.34" />
                    <SPLIT distance="350" swimtime="00:06:32.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="109" reactiontime="+68" swimtime="00:00:50.15" resultid="18514" heatid="19033" lane="3" entrytime="00:00:50.81" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mieszko" lastname="Nowacki" birthdate="2009-11-06" gender="M" nation="POL" license="102503700136" swrid="5173031" athleteid="18488">
              <RESULTS>
                <RESULT eventid="1063" points="222" reactiontime="+78" swimtime="00:00:34.53" resultid="18489" heatid="18953" lane="1" />
                <RESULT eventid="1095" points="255" reactiontime="+87" swimtime="00:02:56.42" resultid="18490" heatid="18996" lane="6" entrytime="00:03:00.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.99" />
                    <SPLIT distance="100" swimtime="00:01:29.11" />
                    <SPLIT distance="150" swimtime="00:02:15.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="239" reactiontime="+91" swimtime="00:00:38.64" resultid="18491" heatid="19035" lane="6" entrytime="00:00:38.50" entrycourse="LCM" />
                <RESULT eventid="1145" points="245" reactiontime="+81" swimtime="00:03:02.14" resultid="18492" heatid="19053" lane="1" entrytime="00:03:06.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.45" />
                    <SPLIT distance="100" swimtime="00:01:25.56" />
                    <SPLIT distance="150" swimtime="00:02:24.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Adamiec" birthdate="2008-03-01" gender="M" nation="POL" license="102503700205" swrid="5462113" athleteid="18493">
              <RESULTS>
                <RESULT eventid="1063" points="185" reactiontime="+74" swimtime="00:00:36.65" resultid="18494" heatid="18956" lane="1" entrytime="00:00:36.81" entrycourse="LCM" />
                <RESULT eventid="1087" points="163" reactiontime="+77" swimtime="00:03:06.40" resultid="18495" heatid="18988" lane="8" entrytime="00:03:06.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.14" />
                    <SPLIT distance="100" swimtime="00:01:30.97" />
                    <SPLIT distance="150" swimtime="00:02:21.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="78" reactiontime="+81" swimtime="00:00:51.91" resultid="18496" heatid="19020" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dagmara" lastname="Mazurek" birthdate="2009-04-15" gender="F" nation="POL" license="102503600145" swrid="5225190" athleteid="18482">
              <RESULTS>
                <RESULT eventid="1059" points="437" reactiontime="+80" swimtime="00:00:31.19" resultid="18483" heatid="18949" lane="7" entrytime="00:00:31.22" entrycourse="LCM" />
                <RESULT eventid="1083" points="425" reactiontime="+86" swimtime="00:02:30.24" resultid="18484" heatid="18983" lane="3" entrytime="00:02:30.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                    <SPLIT distance="100" swimtime="00:01:13.95" />
                    <SPLIT distance="150" swimtime="00:01:53.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="394" reactiontime="+74" swimtime="00:05:22.35" resultid="18485" heatid="19006" lane="9" entrytime="00:05:18.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                    <SPLIT distance="100" swimtime="00:01:12.73" />
                    <SPLIT distance="150" swimtime="00:01:53.45" />
                    <SPLIT distance="200" swimtime="00:02:34.87" />
                    <SPLIT distance="250" swimtime="00:03:17.66" />
                    <SPLIT distance="300" swimtime="00:04:00.62" />
                    <SPLIT distance="350" swimtime="00:04:42.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="426" reactiontime="+68" swimtime="00:01:08.68" resultid="18486" heatid="19064" lane="9" entrytime="00:01:08.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="400" swimtime="00:10:57.46" resultid="18487" heatid="19096" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                    <SPLIT distance="100" swimtime="00:01:16.84" />
                    <SPLIT distance="150" swimtime="00:01:58.04" />
                    <SPLIT distance="200" swimtime="00:02:39.27" />
                    <SPLIT distance="250" swimtime="00:03:20.66" />
                    <SPLIT distance="300" swimtime="00:04:01.89" />
                    <SPLIT distance="350" swimtime="00:04:43.58" />
                    <SPLIT distance="400" swimtime="00:05:25.68" />
                    <SPLIT distance="450" swimtime="00:06:07.70" />
                    <SPLIT distance="500" swimtime="00:06:49.96" />
                    <SPLIT distance="550" swimtime="00:07:32.35" />
                    <SPLIT distance="600" swimtime="00:08:14.56" />
                    <SPLIT distance="650" swimtime="00:08:57.03" />
                    <SPLIT distance="700" swimtime="00:09:38.30" />
                    <SPLIT distance="750" swimtime="00:10:18.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Liubomyr" lastname="Yaremko" birthdate="2007-03-02" gender="M" nation="POL" license="102503700142" swrid="5339633" athleteid="18503">
              <RESULTS>
                <RESULT eventid="1063" points="265" swimtime="00:00:32.53" resultid="18504" heatid="18953" lane="9" />
                <RESULT eventid="1071" points="348" reactiontime="+73" swimtime="00:00:36.88" resultid="18505" heatid="18973" lane="8" entrytime="00:00:37.81" entrycourse="LCM" />
                <RESULT eventid="1121" points="281" reactiontime="+68" swimtime="00:00:36.62" resultid="18506" heatid="19035" lane="5" entrytime="00:00:36.27" entrycourse="LCM" />
                <RESULT eventid="1137" points="330" reactiontime="+70" swimtime="00:01:22.25" resultid="18507" heatid="19046" lane="2" entrytime="00:01:23.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="275" reactiontime="+75" swimtime="00:01:12.05" resultid="18508" heatid="19067" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="296" reactiontime="+72" swimtime="00:01:17.79" resultid="18509" heatid="19086" lane="2" entrytime="00:01:19.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03603" nation="POL" region="03" clubid="18582" name="Wodniacki UKS SP 30">
          <ATHLETES>
            <ATHLETE firstname="Mateusz" lastname="Hunek" birthdate="2009-11-29" gender="M" nation="POL" license="103603700025" swrid="5353672" athleteid="18613">
              <RESULTS>
                <RESULT eventid="1071" points="232" swimtime="00:00:42.21" resultid="18614" heatid="18972" lane="9" entrytime="00:00:41.80" entrycourse="LCM" />
                <RESULT eventid="1137" points="233" reactiontime="+75" swimtime="00:01:32.33" resultid="18615" heatid="19045" lane="4" entrytime="00:01:33.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="250" reactiontime="+74" swimtime="00:03:20.16" resultid="18616" heatid="19093" lane="6" entrytime="00:03:19.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.17" />
                    <SPLIT distance="100" swimtime="00:01:35.41" />
                    <SPLIT distance="150" swimtime="00:02:28.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Zdanowicz" birthdate="2008-03-15" gender="M" nation="POL" license="103603700046" swrid="5043816" athleteid="18601">
              <RESULTS>
                <RESULT eventid="1063" points="139" reactiontime="+93" swimtime="00:00:40.34" resultid="18602" heatid="18955" lane="6" entrytime="00:00:39.41" entrycourse="LCM" />
                <RESULT eventid="1071" points="106" reactiontime="+92" swimtime="00:00:54.82" resultid="18603" heatid="18970" lane="1" entrytime="00:00:51.05" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daria" lastname="Krysiak" birthdate="2009-07-02" gender="F" nation="POL" license="103603600029" swrid="5288474" athleteid="18583">
              <RESULTS>
                <RESULT eventid="1059" points="149" reactiontime="+84" swimtime="00:00:44.56" resultid="18584" heatid="18946" lane="5" entrytime="00:00:42.02" entrycourse="LCM" />
                <RESULT eventid="1067" points="137" reactiontime="+96" swimtime="00:00:56.90" resultid="18585" heatid="18964" lane="5" entrytime="00:00:54.52" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miłosz" lastname="Parol" birthdate="2009-08-02" gender="M" nation="POL" license="103603700038" swrid="5204669" athleteid="18609">
              <RESULTS>
                <RESULT eventid="1071" points="180" reactiontime="+78" swimtime="00:00:45.90" resultid="18610" heatid="18970" lane="5" entrytime="00:00:46.95" entrycourse="LCM" />
                <RESULT eventid="1137" points="163" reactiontime="+81" swimtime="00:01:43.93" resultid="18611" heatid="19044" lane="7" entrytime="00:01:43.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="165" swimtime="00:03:49.75" resultid="18612" heatid="19092" lane="5" entrytime="00:03:45.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.26" />
                    <SPLIT distance="100" swimtime="00:01:52.31" />
                    <SPLIT distance="150" swimtime="00:02:51.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Remigiusz" lastname="Wójcik" birthdate="2009-02-12" gender="M" nation="POL" license="103603700037" swrid="5204675" athleteid="18604">
              <RESULTS>
                <RESULT eventid="1063" points="294" swimtime="00:00:31.44" resultid="18605" heatid="18959" lane="9" entrytime="00:00:31.18" entrycourse="LCM" />
                <RESULT eventid="1079" points="208" reactiontime="+83" swimtime="00:01:23.52" resultid="18606" heatid="18979" lane="4" entrytime="00:01:21.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="259" swimtime="00:00:34.91" resultid="18607" heatid="19022" lane="0" entrytime="00:00:36.64" entrycourse="LCM" />
                <RESULT eventid="1163" points="282" reactiontime="+77" swimtime="00:01:11.52" resultid="18608" heatid="19072" lane="2" entrytime="00:01:11.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martyna" lastname="Hałas" birthdate="2001-08-03" gender="F" nation="POL" license="103603600073" swrid="5453689" athleteid="18589">
              <RESULTS>
                <RESULT eventid="1059" points="295" reactiontime="+81" swimtime="00:00:35.55" resultid="18590" heatid="18948" lane="1" entrytime="00:00:35.00" entrycourse="LCM" />
                <RESULT eventid="1067" points="221" reactiontime="+83" swimtime="00:00:48.59" resultid="18591" heatid="18965" lane="7" entrytime="00:00:49.06" entrycourse="LCM" />
                <RESULT eventid="1108" points="208" reactiontime="+79" swimtime="00:00:41.22" resultid="18592" heatid="19013" lane="4" />
                <RESULT eventid="1159" points="261" reactiontime="+79" swimtime="00:01:20.86" resultid="18593" heatid="19061" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Błaziak" birthdate="2009-09-26" gender="F" nation="POL" license="103603600039" swrid="5431065" athleteid="18586">
              <RESULTS>
                <RESULT eventid="1059" points="149" reactiontime="+99" swimtime="00:00:44.57" resultid="18587" heatid="18946" lane="6" entrytime="00:00:46.35" entrycourse="LCM" />
                <RESULT eventid="1067" points="175" reactiontime="+99" swimtime="00:00:52.51" resultid="18588" heatid="18964" lane="3" entrytime="00:00:54.95" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Serewa" birthdate="2009-06-01" gender="M" nation="POL" license="103603700033" swrid="5204698" athleteid="18594">
              <RESULTS>
                <RESULT eventid="1063" points="177" swimtime="00:00:37.21" resultid="18595" heatid="18956" lane="9" entrytime="00:00:37.46" entrycourse="LCM" />
                <RESULT eventid="1071" points="124" swimtime="00:00:51.98" resultid="18596" heatid="18970" lane="2" entrytime="00:00:49.33" entrycourse="LCM" />
                <RESULT eventid="1121" points="174" reactiontime="+73" swimtime="00:00:42.96" resultid="18597" heatid="19032" lane="2" />
                <RESULT eventid="1145" points="178" reactiontime="+83" swimtime="00:03:22.57" resultid="18598" heatid="19052" lane="4" entrytime="00:03:19.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.03" />
                    <SPLIT distance="100" swimtime="00:01:39.96" />
                    <SPLIT distance="150" swimtime="00:02:39.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="177" reactiontime="+80" swimtime="00:01:23.43" resultid="18599" heatid="19069" lane="4" entrytime="00:01:22.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="152" reactiontime="+76" swimtime="00:01:37.11" resultid="18600" heatid="19085" lane="2" entrytime="00:01:35.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01709" nation="POL" region="09" clubid="16872" name="iSwim Białystok">
          <ATHLETES>
            <ATHLETE firstname="Dawid" lastname="Świderski" birthdate="1979-02-13" gender="M" nation="POL" license="517/09700108" swrid="5422007" athleteid="16876">
              <RESULTS>
                <RESULT eventid="1063" points="489" reactiontime="+73" status="EXH" swimtime="00:00:26.54" resultid="16877" heatid="18952" lane="2" />
                <RESULT eventid="1079" points="459" reactiontime="+75" status="EXH" swimtime="00:01:04.16" resultid="16878" heatid="18978" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="494" reactiontime="+74" status="EXH" swimtime="00:00:28.16" resultid="16879" heatid="19019" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Iłendo" birthdate="1993-02-09" gender="M" nation="POL" license="117/09700014" swrid="4086405" athleteid="16884">
              <RESULTS>
                <RESULT eventid="1063" points="536" reactiontime="+60" status="EXH" swimtime="00:00:25.74" resultid="16885" heatid="18954" lane="0" />
                <RESULT eventid="1121" points="494" reactiontime="+62" status="EXH" swimtime="00:00:30.35" resultid="16886" heatid="19031" lane="3" />
                <RESULT eventid="1163" status="DNS" swimtime="00:00:00.00" resultid="16887" heatid="19068" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Magdalena" lastname="Iwaniuk-Mróz" birthdate="1979-07-17" gender="F" nation="POL" license="117/09600024" athleteid="16873">
              <RESULTS>
                <RESULT eventid="1059" points="453" reactiontime="+74" status="EXH" swimtime="00:00:30.80" resultid="16874" heatid="18945" lane="1" />
                <RESULT eventid="1108" points="377" reactiontime="+74" status="EXH" swimtime="00:00:33.80" resultid="16875" heatid="19013" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wieńczysław" lastname="Safrończyk" birthdate="1954-08-27" gender="M" nation="POL" license="517/09700079" athleteid="16888">
              <RESULTS>
                <RESULT eventid="1071" points="104" status="EXH" swimtime="00:00:55.17" resultid="16889" heatid="18968" lane="6" />
                <RESULT eventid="1137" points="106" reactiontime="+99" status="EXH" swimtime="00:02:00.14" resultid="18943" heatid="19043" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" status="DNS" swimtime="00:00:00.00" resultid="18944" heatid="19092" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sebastian" lastname="Humbla" birthdate="1979-01-24" gender="M" nation="POL" license="117/09700001" athleteid="16880">
              <RESULTS>
                <RESULT eventid="1063" points="432" reactiontime="+67" status="EXH" swimtime="00:00:27.65" resultid="16881" heatid="18953" lane="2" />
                <RESULT eventid="1071" points="361" reactiontime="+67" status="EXH" swimtime="00:00:36.42" resultid="16882" heatid="18969" lane="0" />
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="16883" heatid="19019" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewa" lastname="Markowska" birthdate="1981-03-20" gender="F" nation="POL" license="117/09600015" athleteid="16891">
              <RESULTS>
                <RESULT eventid="1125" points="191" status="EXH" swimtime="00:06:50.56" resultid="16892" heatid="19005" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.63" />
                    <SPLIT distance="100" swimtime="00:01:32.32" />
                    <SPLIT distance="150" swimtime="00:02:25.32" />
                    <SPLIT distance="200" swimtime="00:03:18.63" />
                    <SPLIT distance="250" swimtime="00:04:13.29" />
                    <SPLIT distance="300" swimtime="00:05:07.23" />
                    <SPLIT distance="350" swimtime="00:06:01.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04403" nation="POL" region="03" clubid="17543" name="MKS AVIA Świdnik">
          <ATHLETES>
            <ATHLETE firstname="Michał" lastname="Piekaruś" birthdate="2007-02-03" gender="M" nation="POL" license="104403700003" swrid="5105303" athleteid="17547">
              <RESULTS>
                <RESULT eventid="1063" points="362" reactiontime="+74" swimtime="00:00:29.32" resultid="17548" heatid="18960" lane="8" entrytime="00:00:28.99" entrycourse="LCM" />
                <RESULT eventid="1087" points="399" reactiontime="+73" swimtime="00:02:18.55" resultid="17549" heatid="18987" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.15" />
                    <SPLIT distance="100" swimtime="00:01:06.63" />
                    <SPLIT distance="150" swimtime="00:01:43.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="391" reactiontime="+74" swimtime="00:00:30.45" resultid="17550" heatid="19020" lane="0" />
                <RESULT comment="K14 - Pływak wykonał kopnięcie nóg w płaszczyźnie pionowej w dół (z wyjątkiem jednego ruchu po starcie lub nawrocie)" eventid="1145" reactiontime="+72" status="DSQ" swimtime="00:02:39.70" resultid="17551" heatid="19052" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.21" />
                    <SPLIT distance="100" swimtime="00:01:14.73" />
                    <SPLIT distance="150" swimtime="00:02:04.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="435" reactiontime="+75" swimtime="00:01:01.87" resultid="17552" heatid="19073" lane="4" entrytime="00:01:03.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Maciocha" birthdate="2006-04-14" gender="M" nation="POL" license="104403700005" swrid="5225177" athleteid="17558">
              <RESULTS>
                <RESULT eventid="1063" points="318" reactiontime="+63" swimtime="00:00:30.61" resultid="17559" heatid="18952" lane="9" />
                <RESULT eventid="1095" points="288" reactiontime="+73" swimtime="00:02:49.37" resultid="17560" heatid="18996" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                    <SPLIT distance="100" swimtime="00:01:20.93" />
                    <SPLIT distance="150" swimtime="00:02:06.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="353" reactiontime="+70" swimtime="00:00:33.95" resultid="17561" heatid="19036" lane="8" entrytime="00:00:34.32" entrycourse="LCM" />
                <RESULT eventid="1171" points="326" reactiontime="+70" swimtime="00:01:15.28" resultid="17562" heatid="19086" lane="5" entrytime="00:01:15.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Czeczko" birthdate="2006-05-11" gender="M" nation="POL" license="104403700002" swrid="4827530" athleteid="17571">
              <RESULTS>
                <RESULT eventid="1079" points="420" reactiontime="+68" swimtime="00:01:06.09" resultid="17572" heatid="18980" lane="1" entrytime="00:01:08.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="407" reactiontime="+66" swimtime="00:05:28.85" resultid="17573" heatid="19001" lane="1" entrytime="00:05:40.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                    <SPLIT distance="100" swimtime="00:01:09.56" />
                    <SPLIT distance="150" swimtime="00:01:53.74" />
                    <SPLIT distance="200" swimtime="00:02:36.41" />
                    <SPLIT distance="250" swimtime="00:03:25.44" />
                    <SPLIT distance="300" swimtime="00:04:14.80" />
                    <SPLIT distance="350" swimtime="00:04:53.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="413" reactiontime="+74" swimtime="00:00:29.90" resultid="17574" heatid="19023" lane="7" entrytime="00:00:30.68" entrycourse="LCM" />
                <RESULT eventid="1145" points="409" reactiontime="+72" swimtime="00:02:33.47" resultid="17575" heatid="19053" lane="4" entrytime="00:02:37.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                    <SPLIT distance="100" swimtime="00:01:11.28" />
                    <SPLIT distance="150" swimtime="00:01:59.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="404" reactiontime="+75" swimtime="00:02:29.76" resultid="17576" heatid="19059" lane="0" entrytime="00:02:43.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.37" />
                    <SPLIT distance="100" swimtime="00:01:09.89" />
                    <SPLIT distance="150" swimtime="00:01:48.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patryk" lastname="Lis" birthdate="1998-03-11" gender="M" nation="POL" license="104403700007" swrid="4435930" athleteid="17563">
              <RESULTS>
                <RESULT eventid="1071" points="602" reactiontime="+75" swimtime="00:00:30.72" resultid="17564" heatid="18974" lane="3" entrytime="00:00:30.73" entrycourse="LCM" />
                <RESULT eventid="1113" points="566" reactiontime="+76" swimtime="00:00:26.92" resultid="17565" heatid="19025" lane="9" entrytime="00:00:27.53" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emil" lastname="Krzykała" birthdate="2001-02-01" gender="M" nation="POL" license="104403700006" swrid="4485610" athleteid="17544">
              <RESULTS>
                <RESULT eventid="1063" points="600" reactiontime="+71" swimtime="00:00:24.79" resultid="17545" heatid="18962" lane="6" entrytime="00:00:24.94" entrycourse="LCM" />
                <RESULT eventid="1113" points="596" reactiontime="+71" swimtime="00:00:26.46" resultid="17546" heatid="19025" lane="3" entrytime="00:00:26.04" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tymoteusz" lastname="Sawka" birthdate="2009-07-09" gender="M" nation="POL" license="104403700001" swrid="5448198" athleteid="17553">
              <RESULTS>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej, a przed sygnałem startu" eventid="1063" status="DSQ" swimtime="00:00:31.63" resultid="17554" heatid="18958" lane="0" entrytime="00:00:32.57" entrycourse="LCM" />
                <RESULT eventid="1087" points="286" reactiontime="+68" swimtime="00:02:34.67" resultid="17555" heatid="18989" lane="1" entrytime="00:02:39.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                    <SPLIT distance="100" swimtime="00:01:14.92" />
                    <SPLIT distance="150" swimtime="00:01:57.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="258" reactiontime="+75" swimtime="00:00:34.94" resultid="17556" heatid="19021" lane="6" entrytime="00:00:39.55" entrycourse="LCM" />
                <RESULT eventid="1163" points="301" reactiontime="+61" swimtime="00:01:09.93" resultid="17557" heatid="19071" lane="3" entrytime="00:01:14.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrian" lastname="Maciąg" birthdate="2007-01-18" gender="M" nation="POL" license="104403700004" swrid="5345132" athleteid="17567">
              <RESULTS>
                <RESULT eventid="1071" points="338" reactiontime="+80" swimtime="00:00:37.25" resultid="17568" heatid="18972" lane="5" entrytime="00:00:38.54" entrycourse="LCM" />
                <RESULT eventid="1137" points="335" reactiontime="+69" swimtime="00:01:21.82" resultid="17569" heatid="19046" lane="7" entrytime="00:01:25.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="351" reactiontime="+67" swimtime="00:02:58.79" resultid="17570" heatid="19094" lane="9" entrytime="00:03:10.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.34" />
                    <SPLIT distance="100" swimtime="00:01:26.41" />
                    <SPLIT distance="150" swimtime="00:02:14.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04103" nation="POL" region="03" clubid="17921" name="Swim Team Lubartów">
          <ATHLETES>
            <ATHLETE firstname="Kaja" lastname="Czakon" birthdate="2009-09-22" gender="F" nation="POL" license="104103600009" swrid="5173255" athleteid="17943">
              <RESULTS>
                <RESULT eventid="1067" points="176" swimtime="00:00:52.43" resultid="17944" heatid="18964" lane="0" />
                <RESULT eventid="1117" points="235" reactiontime="+79" swimtime="00:00:43.68" resultid="17945" heatid="19027" lane="3" entrytime="00:00:43.52" entrycourse="LCM" />
                <RESULT eventid="1133" points="156" reactiontime="+82" swimtime="00:01:59.04" resultid="17946" heatid="19039" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="213" swimtime="00:01:26.57" resultid="17947" heatid="19062" lane="0" entrytime="00:01:25.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="203" reactiontime="+84" swimtime="00:01:37.84" resultid="17948" heatid="19079" lane="4" entrytime="00:01:34.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1091" points="236" reactiontime="+74" status="EXH" swimtime="00:03:19.49" resultid="19108" heatid="18992" lane="6" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.70" />
                    <SPLIT distance="100" swimtime="00:01:40.65" />
                    <SPLIT distance="150" swimtime="00:02:32.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kaja" lastname="Wróblewska" birthdate="2007-11-22" gender="F" nation="POL" license="104103600002" swrid="5082974" athleteid="17956">
              <RESULTS>
                <RESULT eventid="1075" points="399" reactiontime="+76" swimtime="00:01:15.31" resultid="17957" heatid="18976" lane="7" entrytime="00:01:16.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1091" points="425" reactiontime="+81" swimtime="00:02:44.02" resultid="17958" heatid="18993" lane="5" entrytime="00:02:41.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.71" />
                    <SPLIT distance="100" swimtime="00:01:21.54" />
                    <SPLIT distance="150" swimtime="00:02:04.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="454" reactiontime="+74" swimtime="00:00:31.78" resultid="17959" heatid="19016" lane="6" entrytime="00:00:32.59" entrycourse="LCM" />
                <RESULT eventid="1150" points="317" reactiontime="+77" swimtime="00:02:58.48" resultid="17960" heatid="19057" lane="0" entrytime="00:02:59.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.12" />
                    <SPLIT distance="100" swimtime="00:01:25.74" />
                    <SPLIT distance="150" swimtime="00:02:13.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="434" reactiontime="+77" swimtime="00:01:08.28" resultid="17961" heatid="19064" lane="0" entrytime="00:01:08.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="399" reactiontime="+80" status="EXH" swimtime="00:01:18.17" resultid="19113" heatid="19078" lane="7" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karol" lastname="Mika" birthdate="2008-09-15" gender="M" nation="POL" license="104103700003" swrid="5173260" athleteid="17949">
              <RESULTS>
                <RESULT eventid="1071" points="259" reactiontime="+54" swimtime="00:00:40.66" resultid="17950" heatid="18972" lane="0" entrytime="00:00:41.79" entrycourse="LCM" />
                <RESULT eventid="1087" points="195" reactiontime="+77" swimtime="00:02:55.66" resultid="17951" heatid="18987" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.94" />
                    <SPLIT distance="100" swimtime="00:01:23.94" />
                    <SPLIT distance="150" swimtime="00:02:10.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="211" reactiontime="+77" swimtime="00:00:37.40" resultid="17952" heatid="19021" lane="3" entrytime="00:00:38.96" entrycourse="LCM" />
                <RESULT eventid="1137" points="230" reactiontime="+87" swimtime="00:01:32.83" resultid="17953" heatid="19045" lane="3" entrytime="00:01:34.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="205" reactiontime="+79" swimtime="00:01:19.47" resultid="17954" heatid="19070" lane="0" entrytime="00:01:19.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="240" reactiontime="+76" swimtime="00:03:22.86" resultid="17955" heatid="19093" lane="3" entrytime="00:03:19.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.89" />
                    <SPLIT distance="100" swimtime="00:01:36.40" />
                    <SPLIT distance="150" swimtime="00:02:30.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Mierzwińska" birthdate="2009-06-17" gender="F" nation="POL" license="104103600016" swrid="5453738" athleteid="17929">
              <RESULTS>
                <RESULT eventid="1059" points="220" swimtime="00:00:39.18" resultid="17930" heatid="18947" lane="0" entrytime="00:00:40.41" entrycourse="LCM" />
                <RESULT eventid="1067" points="220" swimtime="00:00:48.65" resultid="17931" heatid="18965" lane="0" entrytime="00:00:51.64" entrycourse="LCM" />
                <RESULT eventid="1117" points="237" reactiontime="+67" swimtime="00:00:43.58" resultid="17932" heatid="19027" lane="7" entrytime="00:00:44.89" entrycourse="LCM" />
                <RESULT eventid="1133" points="197" swimtime="00:01:50.06" resultid="17933" heatid="19039" lane="6" entrytime="00:02:01.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="165" swimtime="00:01:34.22" resultid="17934" heatid="19061" lane="6" entrytime="00:01:43.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="185" reactiontime="+80" swimtime="00:01:40.92" resultid="17935" heatid="19079" lane="6" entrytime="00:01:45.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Gajos" birthdate="2007-08-31" gender="F" nation="POL" license="104103600023" swrid="5105253" athleteid="17922">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="17923" heatid="18947" lane="1" entrytime="00:00:37.80" entrycourse="LCM" />
                <RESULT eventid="1067" status="DNS" swimtime="00:00:00.00" resultid="17924" heatid="18965" lane="3" entrytime="00:00:46.21" entrycourse="LCM" />
                <RESULT eventid="1117" points="215" reactiontime="+84" swimtime="00:00:44.97" resultid="17925" heatid="19027" lane="5" entrytime="00:00:41.94" entrycourse="LCM" />
                <RESULT eventid="1133" points="217" reactiontime="+95" swimtime="00:01:46.69" resultid="17926" heatid="19038" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="177" swimtime="00:01:32.03" resultid="17927" heatid="19060" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="157" reactiontime="+95" swimtime="00:01:46.65" resultid="17928" heatid="19079" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="08114" nation="POL" region="14" clubid="16838" name="AZS  KU Uniwersytetu Warszawskiego">
          <ATHLETES>
            <ATHLETE firstname="Krzysztof" lastname="Micorek" birthdate="1993-08-25" gender="M" nation="POL" license="108114700041" swrid="4086676" athleteid="16839">
              <RESULTS>
                <RESULT eventid="1063" points="596" reactiontime="+73" status="EXH" swimtime="00:00:24.84" resultid="16840" heatid="18953" lane="3" />
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="16841" heatid="18979" lane="0" />
                <RESULT eventid="1113" points="555" reactiontime="+76" status="EXH" swimtime="00:00:27.09" resultid="16842" heatid="19025" lane="8" entrytime="00:00:27.00" entrycourse="LCM" />
                <RESULT eventid="1163" points="609" reactiontime="+71" status="EXH" swimtime="00:00:55.33" resultid="16843" heatid="19077" lane="9" entrytime="00:00:56.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Godlewski" birthdate="1996-05-26" gender="M" nation="POL" license="108114700059" swrid="4285522" athleteid="16844">
              <RESULTS>
                <RESULT eventid="1071" points="549" reactiontime="+74" status="EXH" swimtime="00:00:31.69" resultid="16845" heatid="18974" lane="2" entrytime="00:00:31.65" entrycourse="LCM" />
                <RESULT eventid="1137" points="497" reactiontime="+66" status="EXH" swimtime="00:01:11.79" resultid="16846" heatid="19047" lane="2" entrytime="00:01:11.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Rębas" birthdate="1989-12-11" gender="M" nation="POL" license="508114700069" swrid="4251117" athleteid="16847">
              <RESULTS>
                <RESULT eventid="1079" points="590" reactiontime="+75" status="EXH" swimtime="00:00:59.01" resultid="16848" heatid="18981" lane="3" entrytime="00:00:59.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="524" reactiontime="+72" status="EXH" swimtime="00:00:27.61" resultid="16849" heatid="19025" lane="0" entrytime="00:00:27.18" entrycourse="LCM" />
                <RESULT eventid="1163" points="602" reactiontime="+76" status="EXH" swimtime="00:00:55.54" resultid="16850" heatid="19077" lane="7" entrytime="00:00:54.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01503" nation="POL" region="03" clubid="18099" name="Uks &quot;Kraszak&quot;">
          <ATHLETES>
            <ATHLETE firstname="Gabriela" lastname="Sieczko" birthdate="2008-12-06" gender="F" nation="POL" license="101503600019" swrid="5455435" athleteid="18100">
              <RESULTS>
                <RESULT eventid="1059" points="278" reactiontime="+91" swimtime="00:00:36.24" resultid="18101" heatid="18947" lane="3" entrytime="00:00:37.12" entrycourse="LCM" />
                <RESULT eventid="1067" points="224" swimtime="00:00:48.36" resultid="18102" heatid="18965" lane="8" entrytime="00:00:50.12" entrycourse="LCM" />
                <RESULT eventid="1117" points="227" reactiontime="+82" swimtime="00:00:44.18" resultid="18103" heatid="19027" lane="1" entrytime="00:00:45.57" entrycourse="LCM" />
                <RESULT comment="K14 - Pływak wykonał kopnięcie nóg w płaszczyźnie pionowej w dół (z wyjątkiem jednego ruchu po starcie lub nawrocie)" eventid="1133" reactiontime="+93" status="DSQ" swimtime="00:01:43.82" resultid="18104" heatid="19039" lane="3" entrytime="00:01:47.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="230" reactiontime="+86" swimtime="00:01:24.30" resultid="18105" heatid="19062" lane="9" entrytime="00:01:25.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="207" reactiontime="+84" swimtime="00:01:37.22" resultid="18106" heatid="19078" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Toczek" birthdate="2003-10-14" gender="M" nation="POL" license="101503700001" swrid="4980283" athleteid="18132">
              <RESULTS>
                <RESULT eventid="1063" points="479" reactiontime="+75" swimtime="00:00:26.71" resultid="18133" heatid="18961" lane="1" entrytime="00:00:26.78" entrycourse="LCM" />
                <RESULT eventid="1071" points="443" reactiontime="+80" swimtime="00:00:34.04" resultid="18134" heatid="18974" lane="8" entrytime="00:00:33.67" entrycourse="LCM" />
                <RESULT eventid="1113" points="484" reactiontime="+76" swimtime="00:00:28.35" resultid="18135" heatid="19024" lane="0" entrytime="00:00:28.86" entrycourse="LCM" />
                <RESULT eventid="1137" points="440" reactiontime="+77" swimtime="00:01:14.77" resultid="18136" heatid="19047" lane="1" entrytime="00:01:13.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="546" reactiontime="+74" swimtime="00:00:57.37" resultid="18137" heatid="19075" lane="3" entrytime="00:00:58.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="457" reactiontime="+82" swimtime="00:02:43.67" resultid="18138" heatid="19094" lane="2" entrytime="00:02:42.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                    <SPLIT distance="100" swimtime="00:01:18.34" />
                    <SPLIT distance="150" swimtime="00:02:01.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Lustyk" birthdate="2009-07-04" gender="F" nation="POL" license="101503600017" athleteid="18127">
              <RESULTS>
                <RESULT eventid="1059" points="151" reactiontime="+95" swimtime="00:00:44.41" resultid="18128" heatid="18945" lane="5" />
                <RESULT eventid="1067" points="118" reactiontime="+88" swimtime="00:00:59.89" resultid="18129" heatid="18963" lane="3" />
                <RESULT eventid="1117" points="134" reactiontime="+72" swimtime="00:00:52.72" resultid="18130" heatid="19027" lane="9" />
                <RESULT eventid="1159" points="134" reactiontime="+86" swimtime="00:01:40.96" resultid="18131" heatid="19061" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Kołodziejak" birthdate="2007-02-09" gender="F" nation="POL" license="101503600018" swrid="5455432" athleteid="18120">
              <RESULTS>
                <RESULT eventid="1059" points="248" reactiontime="+88" swimtime="00:00:37.63" resultid="18121" heatid="18947" lane="6" entrytime="00:00:37.34" entrycourse="LCM" />
                <RESULT eventid="1067" points="272" reactiontime="+92" swimtime="00:00:45.35" resultid="18122" heatid="18965" lane="5" entrytime="00:00:46.15" entrycourse="LCM" />
                <RESULT eventid="1117" points="237" reactiontime="+76" swimtime="00:00:43.55" resultid="18123" heatid="19027" lane="2" entrytime="00:00:43.86" entrycourse="LCM" />
                <RESULT eventid="1133" points="272" reactiontime="+85" swimtime="00:01:38.95" resultid="18124" heatid="19040" lane="9" entrytime="00:01:39.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="226" reactiontime="+96" swimtime="00:01:24.79" resultid="18125" heatid="19061" lane="5" entrytime="00:01:28.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="273" swimtime="00:03:34.30" resultid="18126" heatid="19090" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.03" />
                    <SPLIT distance="100" swimtime="00:01:42.21" />
                    <SPLIT distance="150" swimtime="00:02:38.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patrycja" lastname="Chwedoruk" birthdate="2008-09-17" gender="F" nation="POL" license="101503600014" swrid="5085424" athleteid="18107">
              <RESULTS>
                <RESULT eventid="1059" points="224" swimtime="00:00:38.97" resultid="18108" heatid="18947" lane="9" entrytime="00:00:40.71" entrycourse="LCM" />
                <RESULT eventid="1075" points="150" reactiontime="+99" swimtime="00:01:44.20" resultid="18109" heatid="18975" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="189" reactiontime="+83" swimtime="00:00:42.51" resultid="18110" heatid="19014" lane="5" entrytime="00:00:47.21" entrycourse="LCM" />
                <RESULT eventid="1141" points="221" reactiontime="+84" swimtime="00:03:28.41" resultid="18111" heatid="19048" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.26" />
                    <SPLIT distance="100" swimtime="00:01:38.80" />
                    <SPLIT distance="150" swimtime="00:02:39.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="200" reactiontime="+80" swimtime="00:01:28.36" resultid="18112" heatid="19061" lane="3" entrytime="00:01:34.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="207" reactiontime="+94" swimtime="00:01:37.25" resultid="18113" heatid="19078" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Chwedoruk" birthdate="2003-10-23" gender="F" nation="POL" license="101503600023" swrid="5455429" athleteid="18114">
              <RESULTS>
                <RESULT eventid="1059" points="283" reactiontime="+71" swimtime="00:00:36.04" resultid="18115" heatid="18947" lane="5" entrytime="00:00:36.82" entrycourse="LCM" />
                <RESULT eventid="1067" points="209" reactiontime="+87" swimtime="00:00:49.50" resultid="18116" heatid="18965" lane="1" entrytime="00:00:49.88" entrycourse="LCM" />
                <RESULT eventid="1108" points="254" reactiontime="+87" swimtime="00:00:38.53" resultid="18117" heatid="19015" lane="8" entrytime="00:00:40.94" entrycourse="LCM" />
                <RESULT eventid="1117" points="233" reactiontime="+89" swimtime="00:00:43.79" resultid="18118" heatid="19026" lane="4" />
                <RESULT eventid="1159" points="269" reactiontime="+76" swimtime="00:01:20.07" resultid="18119" heatid="19062" lane="1" entrytime="00:01:23.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04303" nation="POL" region="03" clubid="17525" name="Masters Avia Świdnik">
          <ATHLETES>
            <ATHLETE firstname="Cezary" lastname="Lipiński" birthdate="1972-04-11" gender="M" nation="POL" license="104303700002" swrid="5449345" athleteid="17526">
              <RESULTS>
                <RESULT eventid="1063" points="317" reactiontime="+73" swimtime="00:00:30.64" resultid="17527" heatid="18953" lane="7" />
                <RESULT eventid="1087" points="298" reactiontime="+73" swimtime="00:02:32.59" resultid="17528" heatid="18986" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="100" swimtime="00:01:12.14" />
                    <SPLIT distance="150" swimtime="00:01:51.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="316" reactiontime="+76" swimtime="00:05:22.84" resultid="17529" heatid="19008" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.97" />
                    <SPLIT distance="100" swimtime="00:01:16.73" />
                    <SPLIT distance="150" swimtime="00:01:57.13" />
                    <SPLIT distance="200" swimtime="00:02:36.98" />
                    <SPLIT distance="250" swimtime="00:03:17.86" />
                    <SPLIT distance="300" swimtime="00:03:59.25" />
                    <SPLIT distance="350" swimtime="00:04:41.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="282" reactiontime="+62" swimtime="00:00:33.96" resultid="17530" heatid="19019" lane="9" />
                <RESULT eventid="1163" points="323" reactiontime="+73" swimtime="00:01:08.30" resultid="17531" heatid="19067" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Sitkowski" birthdate="1974-10-05" gender="M" nation="POL" license="504303700001" swrid="5439542" athleteid="17532">
              <RESULTS>
                <RESULT eventid="1063" points="414" reactiontime="+81" swimtime="00:00:28.04" resultid="17533" heatid="18952" lane="1" />
                <RESULT eventid="1095" points="291" reactiontime="+80" swimtime="00:02:48.84" resultid="17534" heatid="18995" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.13" />
                    <SPLIT distance="100" swimtime="00:01:20.28" />
                    <SPLIT distance="150" swimtime="00:02:05.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="352" reactiontime="+69" swimtime="00:00:33.99" resultid="17535" heatid="19033" lane="7" />
                <RESULT eventid="1145" points="267" reactiontime="+85" swimtime="00:02:56.86" resultid="17536" heatid="19051" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.17" />
                    <SPLIT distance="100" swimtime="00:01:21.12" />
                    <SPLIT distance="150" swimtime="00:02:14.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="331" reactiontime="+75" swimtime="00:01:14.95" resultid="17537" heatid="19083" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Zielonka" birthdate="1986-05-26" gender="M" nation="POL" license="104303700006" swrid="4061691" athleteid="17538">
              <RESULTS>
                <RESULT eventid="1063" points="501" reactiontime="+77" swimtime="00:00:26.31" resultid="17539" heatid="18954" lane="1" />
                <RESULT eventid="1079" points="365" reactiontime="+76" swimtime="00:01:09.21" resultid="17540" heatid="18979" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="463" reactiontime="+79" swimtime="00:00:28.77" resultid="17541" heatid="19020" lane="1" />
                <RESULT eventid="1163" points="517" reactiontime="+76" swimtime="00:00:58.43" resultid="17542" heatid="19067" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02103" nation="POL" region="03" clubid="17503" name="LUKS Orlik">
          <ATHLETES>
            <ATHLETE firstname="Bartosz" lastname="Pawluk" birthdate="2009-10-09" gender="M" nation="POL" license="102103700055" swrid="5204699" athleteid="17511">
              <RESULTS>
                <RESULT eventid="1063" points="151" swimtime="00:00:39.21" resultid="17512" heatid="18953" lane="0" />
                <RESULT eventid="1071" points="116" swimtime="00:00:53.06" resultid="17513" heatid="18970" lane="0" entrytime="00:00:52.19" entrycourse="LCM" />
                <RESULT eventid="1121" points="170" swimtime="00:00:43.30" resultid="17514" heatid="19035" lane="0" entrytime="00:00:43.20" entrycourse="LCM" />
                <RESULT eventid="1137" points="115" reactiontime="+92" swimtime="00:01:56.89" resultid="17515" heatid="19042" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="128" swimtime="00:01:32.92" resultid="17516" heatid="19069" lane="8" entrytime="00:01:31.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="121" swimtime="00:01:44.55" resultid="17517" heatid="19085" lane="9" entrytime="00:01:42.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davyd" lastname="Bubnov" birthdate="2009-01-03" gender="M" nation="POL" license="102103700056" swrid="5172976" athleteid="17518">
              <RESULTS>
                <RESULT eventid="1071" points="224" reactiontime="+92" swimtime="00:00:42.67" resultid="17519" heatid="18971" lane="6" entrytime="00:00:43.17" entrycourse="LCM" />
                <RESULT eventid="1087" points="206" reactiontime="+93" swimtime="00:02:52.45" resultid="17520" heatid="18988" lane="6" entrytime="00:02:53.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                    <SPLIT distance="100" swimtime="00:01:24.67" />
                    <SPLIT distance="150" swimtime="00:02:10.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="187" reactiontime="+91" swimtime="00:00:38.90" resultid="17521" heatid="19018" lane="4" />
                <RESULT eventid="1137" points="212" reactiontime="+87" swimtime="00:01:35.39" resultid="17522" heatid="19046" lane="9" entrytime="00:01:32.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="214" reactiontime="+81" swimtime="00:01:18.42" resultid="17523" heatid="19070" lane="2" entrytime="00:01:17.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="211" reactiontime="+79" swimtime="00:03:31.62" resultid="17524" heatid="19093" lane="1" entrytime="00:03:25.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.92" />
                    <SPLIT distance="100" swimtime="00:01:41.85" />
                    <SPLIT distance="150" swimtime="00:02:37.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ernest" lastname="Czechowski" birthdate="2009-03-25" gender="M" nation="POL" license="102103700057" swrid="5204717" athleteid="17504">
              <RESULTS>
                <RESULT eventid="1063" status="DNS" swimtime="00:00:00.00" resultid="17505" heatid="18956" lane="3" entrytime="00:00:35.21" entrycourse="LCM" />
                <RESULT eventid="1087" points="246" reactiontime="+80" swimtime="00:02:42.58" resultid="17506" heatid="18988" lane="7" entrytime="00:02:59.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                    <SPLIT distance="100" swimtime="00:01:17.08" />
                    <SPLIT distance="150" swimtime="00:02:00.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="17507" heatid="19021" lane="0" entrytime="00:00:43.72" entrycourse="LCM" />
                <RESULT eventid="1121" status="DNS" swimtime="00:00:00.00" resultid="17508" heatid="19034" lane="7" entrytime="00:00:46.60" entrycourse="LCM" />
                <RESULT eventid="1163" points="238" reactiontime="+77" swimtime="00:01:15.63" resultid="17509" heatid="19071" lane="7" entrytime="00:01:14.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" status="DNS" swimtime="00:00:00.00" resultid="17510" heatid="19085" lane="5" entrytime="00:01:30.43" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01703" nation="POL" region="03" clubid="17764" name="RWKS Sparta Biłgoraj">
          <ATHLETES>
            <ATHLETE firstname="Kornel" lastname="Kulanin" birthdate="2009-04-29" gender="M" nation="POL" license="101703700133" swrid="5199320" athleteid="17800">
              <RESULTS>
                <RESULT eventid="1063" points="287" reactiontime="+70" swimtime="00:00:31.69" resultid="17801" heatid="18959" lane="7" entrytime="00:00:30.82" entrycourse="LCM" />
                <RESULT eventid="1079" points="294" reactiontime="+62" swimtime="00:01:14.42" resultid="17802" heatid="18980" lane="9" entrytime="00:01:14.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="277" reactiontime="+71" swimtime="00:05:37.31" resultid="17803" heatid="19009" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                    <SPLIT distance="100" swimtime="00:01:16.51" />
                    <SPLIT distance="150" swimtime="00:01:59.58" />
                    <SPLIT distance="200" swimtime="00:02:42.57" />
                    <SPLIT distance="250" swimtime="00:03:26.10" />
                    <SPLIT distance="300" swimtime="00:04:10.51" />
                    <SPLIT distance="350" swimtime="00:04:54.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="340" swimtime="00:00:31.89" resultid="17804" heatid="19023" lane="9" entrytime="00:00:31.88" entrycourse="LCM" />
                <RESULT eventid="1155" points="264" reactiontime="+61" swimtime="00:02:52.53" resultid="17805" heatid="19059" lane="9" entrytime="00:03:00.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                    <SPLIT distance="100" swimtime="00:01:19.59" />
                    <SPLIT distance="150" swimtime="00:02:05.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="291" reactiontime="+42" swimtime="00:01:10.72" resultid="17806" heatid="19073" lane="8" entrytime="00:01:07.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Mazur" birthdate="2009-03-17" gender="M" nation="POL" license="101703700129" swrid="5199327" athleteid="17807">
              <RESULTS>
                <RESULT eventid="1063" points="197" swimtime="00:00:35.92" resultid="17808" heatid="18956" lane="2" entrytime="00:00:35.68" entrycourse="LCM" />
                <RESULT eventid="1087" points="123" reactiontime="+90" swimtime="00:03:24.92" resultid="17809" heatid="18987" lane="4" entrytime="00:03:19.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.11" />
                    <SPLIT distance="100" swimtime="00:01:38.24" />
                    <SPLIT distance="150" swimtime="00:02:33.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="141" reactiontime="+79" swimtime="00:00:42.75" resultid="17810" heatid="19021" lane="7" entrytime="00:00:42.06" entrycourse="LCM" />
                <RESULT eventid="1137" points="109" reactiontime="+81" swimtime="00:01:59.06" resultid="17811" heatid="19043" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="152" reactiontime="+83" swimtime="00:01:27.88" resultid="17812" heatid="19069" lane="7" entrytime="00:01:27.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="108" reactiontime="+72" swimtime="00:01:48.80" resultid="17813" heatid="19085" lane="8" entrytime="00:01:42.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nataniel" lastname="Kobak" birthdate="2008-01-04" gender="M" nation="POL" license="101703700121" swrid="5173002" athleteid="17864">
              <RESULTS>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej, a przed sygnałem startu" eventid="1087" reactiontime="+46" status="DSQ" swimtime="00:02:16.20" resultid="17865" heatid="18990" lane="6" entrytime="00:02:15.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                    <SPLIT distance="100" swimtime="00:01:05.49" />
                    <SPLIT distance="150" swimtime="00:01:41.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6365" points="448" reactiontime="+71" swimtime="00:09:50.80" resultid="17866" heatid="19002" lane="6" entrytime="00:10:20.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                    <SPLIT distance="100" swimtime="00:01:09.59" />
                    <SPLIT distance="150" swimtime="00:01:47.28" />
                    <SPLIT distance="200" swimtime="00:02:24.42" />
                    <SPLIT distance="250" swimtime="00:03:02.27" />
                    <SPLIT distance="300" swimtime="00:03:39.64" />
                    <SPLIT distance="350" swimtime="00:04:17.53" />
                    <SPLIT distance="400" swimtime="00:04:55.13" />
                    <SPLIT distance="450" swimtime="00:05:32.86" />
                    <SPLIT distance="500" swimtime="00:06:10.60" />
                    <SPLIT distance="550" swimtime="00:06:48.36" />
                    <SPLIT distance="600" swimtime="00:07:26.06" />
                    <SPLIT distance="650" swimtime="00:08:03.89" />
                    <SPLIT distance="700" swimtime="00:08:40.72" />
                    <SPLIT distance="750" swimtime="00:09:16.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="441" reactiontime="+63" swimtime="00:04:48.95" resultid="17867" heatid="19010" lane="3" entrytime="00:04:50.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.53" />
                    <SPLIT distance="100" swimtime="00:01:07.79" />
                    <SPLIT distance="150" swimtime="00:01:44.49" />
                    <SPLIT distance="200" swimtime="00:02:22.02" />
                    <SPLIT distance="250" swimtime="00:02:59.34" />
                    <SPLIT distance="300" swimtime="00:03:37.21" />
                    <SPLIT distance="350" swimtime="00:04:13.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="404" reactiontime="+68" swimtime="00:00:32.46" resultid="17868" heatid="19037" lane="9" entrytime="00:00:33.01" entrycourse="LCM" />
                <RESULT eventid="1163" points="432" reactiontime="+57" swimtime="00:01:02.01" resultid="17869" heatid="19073" lane="5" entrytime="00:01:03.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="387" reactiontime="+67" swimtime="00:01:11.11" resultid="17870" heatid="19087" lane="4" entrytime="00:01:09.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Giruć" birthdate="2009-01-28" gender="M" nation="POL" license="101703700125" swrid="5158182" athleteid="17842">
              <RESULTS>
                <RESULT eventid="1071" points="303" reactiontime="+76" swimtime="00:00:38.62" resultid="17843" heatid="18973" lane="1" entrytime="00:00:37.71" entrycourse="LCM" />
                <RESULT eventid="6365" points="261" reactiontime="+89" swimtime="00:11:47.03" resultid="17844" heatid="19002" lane="1" entrytime="00:11:28.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.01" />
                    <SPLIT distance="100" swimtime="00:01:20.76" />
                    <SPLIT distance="150" swimtime="00:02:04.63" />
                    <SPLIT distance="200" swimtime="00:02:49.36" />
                    <SPLIT distance="250" swimtime="00:03:34.53" />
                    <SPLIT distance="300" swimtime="00:04:18.81" />
                    <SPLIT distance="350" swimtime="00:05:03.58" />
                    <SPLIT distance="400" swimtime="00:05:48.07" />
                    <SPLIT distance="450" swimtime="00:06:33.77" />
                    <SPLIT distance="500" swimtime="00:07:19.01" />
                    <SPLIT distance="550" swimtime="00:08:05.37" />
                    <SPLIT distance="600" swimtime="00:08:51.12" />
                    <SPLIT distance="650" swimtime="00:09:37.05" />
                    <SPLIT distance="700" swimtime="00:10:20.53" />
                    <SPLIT distance="750" swimtime="00:11:04.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1137" points="332" reactiontime="+82" swimtime="00:01:22.08" resultid="17845" heatid="19046" lane="3" entrytime="00:01:20.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="297" reactiontime="+97" swimtime="00:02:50.80" resultid="17846" heatid="19053" lane="6" entrytime="00:02:48.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                    <SPLIT distance="100" swimtime="00:01:21.45" />
                    <SPLIT distance="150" swimtime="00:02:08.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="248" reactiontime="+70" swimtime="00:01:14.58" resultid="17847" heatid="19072" lane="6" entrytime="00:01:10.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" status="DNS" swimtime="00:00:00.00" resultid="17848" heatid="19086" lane="7" entrytime="00:01:20.62" entrycourse="LCM" />
                <RESULT eventid="1179" points="349" reactiontime="+81" swimtime="00:02:59.11" resultid="17849" heatid="19094" lane="0" entrytime="00:02:54.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.12" />
                    <SPLIT distance="100" swimtime="00:01:25.56" />
                    <SPLIT distance="150" swimtime="00:02:12.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcel" lastname="Jonczak" birthdate="2009-03-12" gender="M" nation="POL" license="101703700130" swrid="5204273" athleteid="17878">
              <RESULTS>
                <RESULT eventid="1087" points="308" reactiontime="+66" swimtime="00:02:30.95" resultid="17879" heatid="18987" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                    <SPLIT distance="100" swimtime="00:01:11.00" />
                    <SPLIT distance="150" swimtime="00:01:51.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="293" reactiontime="+67" swimtime="00:06:07.05" resultid="17880" heatid="19001" lane="0" entrytime="00:05:59.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                    <SPLIT distance="100" swimtime="00:01:19.12" />
                    <SPLIT distance="150" swimtime="00:02:07.28" />
                    <SPLIT distance="200" swimtime="00:02:52.70" />
                    <SPLIT distance="250" swimtime="00:03:49.91" />
                    <SPLIT distance="300" swimtime="00:04:45.10" />
                    <SPLIT distance="350" swimtime="00:05:27.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="349" reactiontime="+48" swimtime="00:00:31.63" resultid="17881" heatid="19023" lane="0" entrytime="00:00:31.23" entrycourse="LCM" />
                <RESULT eventid="1121" points="363" reactiontime="+69" swimtime="00:00:33.63" resultid="17882" heatid="19036" lane="6" entrytime="00:00:33.28" entrycourse="LCM" />
                <RESULT eventid="1163" points="345" reactiontime="+67" swimtime="00:01:06.85" resultid="17883" heatid="19073" lane="6" entrytime="00:01:04.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="298" reactiontime="+66" swimtime="00:01:17.57" resultid="17884" heatid="19087" lane="8" entrytime="00:01:13.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Bury" birthdate="2007-07-02" gender="M" nation="POL" license="101703700095" swrid="5098668" athleteid="17828">
              <RESULTS>
                <RESULT eventid="1071" points="400" reactiontime="+47" swimtime="00:00:35.21" resultid="17829" heatid="18974" lane="0" entrytime="00:00:34.92" entrycourse="LCM" />
                <RESULT eventid="1103" points="460" reactiontime="+76" swimtime="00:05:15.76" resultid="17830" heatid="19001" lane="6" entrytime="00:05:16.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                    <SPLIT distance="100" swimtime="00:01:12.13" />
                    <SPLIT distance="150" swimtime="00:01:54.80" />
                    <SPLIT distance="200" swimtime="00:02:38.71" />
                    <SPLIT distance="250" swimtime="00:03:21.94" />
                    <SPLIT distance="300" swimtime="00:04:07.18" />
                    <SPLIT distance="350" swimtime="00:04:43.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1137" points="418" reactiontime="+65" swimtime="00:01:16.03" resultid="17831" heatid="19047" lane="0" entrytime="00:01:15.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="455" reactiontime="+56" swimtime="00:02:28.16" resultid="17832" heatid="19054" lane="8" entrytime="00:02:23.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.45" />
                    <SPLIT distance="100" swimtime="00:01:11.43" />
                    <SPLIT distance="150" swimtime="00:01:55.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="415" reactiontime="+69" swimtime="00:01:09.49" resultid="17833" heatid="19088" lane="9" entrytime="00:01:08.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="463" reactiontime="+69" swimtime="00:02:42.99" resultid="17834" heatid="19094" lane="7" entrytime="00:02:45.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.08" />
                    <SPLIT distance="100" swimtime="00:01:19.21" />
                    <SPLIT distance="150" swimtime="00:02:02.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="449" reactiontime="+59" status="EXH" swimtime="00:00:27.30" resultid="19107" heatid="18958" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartłomiej" lastname="Obszyński" birthdate="2007-04-28" gender="M" nation="POL" license="101703700108" swrid="5098679" athleteid="17850">
              <RESULTS>
                <RESULT eventid="1079" points="389" reactiontime="+69" swimtime="00:01:07.79" resultid="17851" heatid="18980" lane="8" entrytime="00:01:09.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6365" points="471" reactiontime="+77" swimtime="00:09:40.83" resultid="17852" heatid="19002" lane="3" entrytime="00:10:15.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.20" />
                    <SPLIT distance="100" swimtime="00:01:06.85" />
                    <SPLIT distance="150" swimtime="00:01:43.06" />
                    <SPLIT distance="200" swimtime="00:02:19.46" />
                    <SPLIT distance="250" swimtime="00:02:55.78" />
                    <SPLIT distance="300" swimtime="00:03:33.08" />
                    <SPLIT distance="350" swimtime="00:04:10.02" />
                    <SPLIT distance="400" swimtime="00:04:47.62" />
                    <SPLIT distance="450" swimtime="00:05:24.64" />
                    <SPLIT distance="500" swimtime="00:06:01.34" />
                    <SPLIT distance="550" swimtime="00:06:38.03" />
                    <SPLIT distance="600" swimtime="00:07:16.08" />
                    <SPLIT distance="650" swimtime="00:07:52.66" />
                    <SPLIT distance="700" swimtime="00:08:29.32" />
                    <SPLIT distance="750" swimtime="00:09:04.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="449" reactiontime="+71" swimtime="00:04:47.29" resultid="17853" heatid="19010" lane="5" entrytime="00:04:47.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                    <SPLIT distance="100" swimtime="00:01:07.35" />
                    <SPLIT distance="150" swimtime="00:01:44.81" />
                    <SPLIT distance="200" swimtime="00:02:21.74" />
                    <SPLIT distance="250" swimtime="00:02:58.71" />
                    <SPLIT distance="300" swimtime="00:03:35.99" />
                    <SPLIT distance="350" swimtime="00:04:12.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="395" reactiontime="+77" swimtime="00:00:30.34" resultid="17854" heatid="19023" lane="1" entrytime="00:00:30.90" entrycourse="LCM" />
                <RESULT eventid="1163" points="423" reactiontime="+71" swimtime="00:01:02.46" resultid="17855" heatid="19074" lane="0" entrytime="00:01:03.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="494" reactiontime="+73" swimtime="00:18:21.48" resultid="17856" heatid="19099" lane="5" entrytime="00:19:24.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                    <SPLIT distance="100" swimtime="00:01:07.68" />
                    <SPLIT distance="150" swimtime="00:01:44.39" />
                    <SPLIT distance="200" swimtime="00:02:21.03" />
                    <SPLIT distance="250" swimtime="00:02:58.52" />
                    <SPLIT distance="300" swimtime="00:03:35.70" />
                    <SPLIT distance="350" swimtime="00:04:13.18" />
                    <SPLIT distance="400" swimtime="00:04:50.94" />
                    <SPLIT distance="450" swimtime="00:05:28.44" />
                    <SPLIT distance="500" swimtime="00:06:05.53" />
                    <SPLIT distance="550" swimtime="00:06:42.57" />
                    <SPLIT distance="600" swimtime="00:07:19.69" />
                    <SPLIT distance="650" swimtime="00:07:57.91" />
                    <SPLIT distance="700" swimtime="00:08:35.34" />
                    <SPLIT distance="750" swimtime="00:09:11.67" />
                    <SPLIT distance="800" swimtime="00:09:48.42" />
                    <SPLIT distance="850" swimtime="00:10:25.64" />
                    <SPLIT distance="900" swimtime="00:11:02.35" />
                    <SPLIT distance="950" swimtime="00:11:39.51" />
                    <SPLIT distance="1000" swimtime="00:12:16.69" />
                    <SPLIT distance="1050" swimtime="00:12:53.69" />
                    <SPLIT distance="1100" swimtime="00:13:30.47" />
                    <SPLIT distance="1150" swimtime="00:14:07.37" />
                    <SPLIT distance="1200" swimtime="00:14:44.55" />
                    <SPLIT distance="1250" swimtime="00:15:21.58" />
                    <SPLIT distance="1300" swimtime="00:15:58.45" />
                    <SPLIT distance="1350" swimtime="00:16:36.20" />
                    <SPLIT distance="1400" swimtime="00:17:12.90" />
                    <SPLIT distance="1450" swimtime="00:17:47.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miłosz" lastname="Jagosiak" birthdate="2008-08-04" gender="M" nation="POL" license="101703700115" swrid="5148626" athleteid="17885">
              <RESULTS>
                <RESULT eventid="1095" points="348" reactiontime="+58" swimtime="00:02:39.06" resultid="17886" heatid="18997" lane="9" entrytime="00:02:40.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                    <SPLIT distance="100" swimtime="00:01:17.05" />
                    <SPLIT distance="150" swimtime="00:01:59.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6365" points="350" reactiontime="+82" swimtime="00:10:41.34" resultid="17887" heatid="19002" lane="2" entrytime="00:10:48.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                    <SPLIT distance="100" swimtime="00:01:11.81" />
                    <SPLIT distance="150" swimtime="00:01:51.56" />
                    <SPLIT distance="200" swimtime="00:02:32.05" />
                    <SPLIT distance="250" swimtime="00:03:13.14" />
                    <SPLIT distance="300" swimtime="00:03:54.29" />
                    <SPLIT distance="350" swimtime="00:04:35.40" />
                    <SPLIT distance="400" swimtime="00:05:17.06" />
                    <SPLIT distance="450" swimtime="00:05:58.42" />
                    <SPLIT distance="500" swimtime="00:06:39.49" />
                    <SPLIT distance="550" swimtime="00:07:20.84" />
                    <SPLIT distance="600" swimtime="00:08:01.03" />
                    <SPLIT distance="650" swimtime="00:08:41.96" />
                    <SPLIT distance="700" swimtime="00:09:22.10" />
                    <SPLIT distance="750" swimtime="00:10:01.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="392" reactiontime="+82" swimtime="00:05:00.56" resultid="17888" heatid="19010" lane="6" entrytime="00:04:59.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                    <SPLIT distance="100" swimtime="00:01:09.97" />
                    <SPLIT distance="150" swimtime="00:01:48.90" />
                    <SPLIT distance="200" swimtime="00:02:27.88" />
                    <SPLIT distance="250" swimtime="00:03:07.21" />
                    <SPLIT distance="300" swimtime="00:03:46.23" />
                    <SPLIT distance="350" swimtime="00:04:25.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="379" reactiontime="+67" swimtime="00:00:33.16" resultid="17889" heatid="19036" lane="3" entrytime="00:00:33.24" entrycourse="LCM" />
                <RESULT eventid="1163" points="379" reactiontime="+85" swimtime="00:01:04.81" resultid="17890" heatid="19073" lane="3" entrytime="00:01:04.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="331" reactiontime="+74" swimtime="00:01:14.93" resultid="17891" heatid="19087" lane="1" entrytime="00:01:13.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Duńko" birthdate="2007-12-11" gender="F" nation="POL" license="101703600097" swrid="5112635" athleteid="17821">
              <RESULTS>
                <RESULT eventid="1067" points="507" reactiontime="+79" swimtime="00:00:36.86" resultid="17822" heatid="18967" lane="8" entrytime="00:00:36.25" entrycourse="LCM" />
                <RESULT eventid="1075" points="487" reactiontime="+94" swimtime="00:01:10.49" resultid="17823" heatid="18977" lane="0" entrytime="00:01:10.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="435" reactiontime="+80" swimtime="00:00:32.24" resultid="17824" heatid="19016" lane="4" entrytime="00:00:31.65" entrycourse="LCM" />
                <RESULT eventid="1133" points="497" reactiontime="+66" swimtime="00:01:20.92" resultid="17825" heatid="19041" lane="8" entrytime="00:01:19.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="517" reactiontime="+85" swimtime="00:01:04.41" resultid="17826" heatid="19065" lane="5" entrytime="00:01:03.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="529" reactiontime="+79" swimtime="00:02:51.99" resultid="17827" heatid="19091" lane="7" entrytime="00:02:54.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.69" />
                    <SPLIT distance="100" swimtime="00:01:22.63" />
                    <SPLIT distance="150" swimtime="00:02:07.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Radosław" lastname="Oszajca" birthdate="2007-04-18" gender="M" nation="POL" license="101703700109" swrid="5098680" athleteid="17786">
              <RESULTS>
                <RESULT eventid="1063" points="323" reactiontime="+78" swimtime="00:00:30.45" resultid="17787" heatid="18958" lane="3" entrytime="00:00:31.35" entrycourse="LCM" />
                <RESULT eventid="1071" points="352" reactiontime="+82" swimtime="00:00:36.74" resultid="17788" heatid="18973" lane="3" entrytime="00:00:36.13" entrycourse="LCM" />
                <RESULT eventid="1113" points="325" reactiontime="+81" swimtime="00:00:32.37" resultid="17789" heatid="19022" lane="5" entrytime="00:00:32.33" entrycourse="LCM" />
                <RESULT eventid="1137" points="321" reactiontime="+85" swimtime="00:01:23.04" resultid="17790" heatid="19046" lane="5" entrytime="00:01:20.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="334" reactiontime="+81" swimtime="00:01:07.56" resultid="17791" heatid="19072" lane="4" entrytime="00:01:08.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="346" reactiontime="+66" swimtime="00:02:59.48" resultid="17792" heatid="19094" lane="8" entrytime="00:02:52.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.31" />
                    <SPLIT distance="100" swimtime="00:01:26.53" />
                    <SPLIT distance="150" swimtime="00:02:14.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kinga" lastname="Cich" birthdate="2007-10-21" gender="F" nation="POL" license="101703600100" swrid="5148624" athleteid="17765">
              <RESULTS>
                <RESULT eventid="1059" points="478" swimtime="00:00:30.27" resultid="17766" heatid="18950" lane="9" entrytime="00:00:30.25" entrycourse="LCM" />
                <RESULT eventid="1091" points="519" reactiontime="+71" swimtime="00:02:33.44" resultid="17767" heatid="18994" lane="1" entrytime="00:02:32.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.69" />
                    <SPLIT distance="100" swimtime="00:01:13.75" />
                    <SPLIT distance="150" swimtime="00:01:52.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="510" reactiontime="+82" swimtime="00:04:55.90" resultid="17768" heatid="19006" lane="6" entrytime="00:04:56.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                    <SPLIT distance="100" swimtime="00:01:07.39" />
                    <SPLIT distance="150" swimtime="00:01:44.04" />
                    <SPLIT distance="200" swimtime="00:02:21.66" />
                    <SPLIT distance="250" swimtime="00:02:59.86" />
                    <SPLIT distance="300" swimtime="00:03:38.49" />
                    <SPLIT distance="350" swimtime="00:04:18.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6361" points="479" reactiontime="+90" swimtime="00:19:36.28" resultid="17769" heatid="19055" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.00" />
                    <SPLIT distance="100" swimtime="00:01:10.87" />
                    <SPLIT distance="150" swimtime="00:01:48.52" />
                    <SPLIT distance="200" swimtime="00:02:27.26" />
                    <SPLIT distance="250" swimtime="00:03:06.25" />
                    <SPLIT distance="300" swimtime="00:03:45.16" />
                    <SPLIT distance="350" swimtime="00:04:24.16" />
                    <SPLIT distance="400" swimtime="00:05:03.34" />
                    <SPLIT distance="450" swimtime="00:05:42.78" />
                    <SPLIT distance="500" swimtime="00:06:22.61" />
                    <SPLIT distance="550" swimtime="00:07:01.83" />
                    <SPLIT distance="600" swimtime="00:07:41.61" />
                    <SPLIT distance="650" swimtime="00:08:21.52" />
                    <SPLIT distance="700" swimtime="00:09:01.19" />
                    <SPLIT distance="750" swimtime="00:09:40.78" />
                    <SPLIT distance="800" swimtime="00:10:20.71" />
                    <SPLIT distance="850" swimtime="00:11:01.04" />
                    <SPLIT distance="900" swimtime="00:11:40.90" />
                    <SPLIT distance="950" swimtime="00:12:20.50" />
                    <SPLIT distance="1000" swimtime="00:13:01.27" />
                    <SPLIT distance="1050" swimtime="00:13:41.06" />
                    <SPLIT distance="1100" swimtime="00:14:20.89" />
                    <SPLIT distance="1150" swimtime="00:15:00.59" />
                    <SPLIT distance="1200" swimtime="00:15:40.62" />
                    <SPLIT distance="1250" swimtime="00:16:20.05" />
                    <SPLIT distance="1300" swimtime="00:16:59.74" />
                    <SPLIT distance="1350" swimtime="00:17:39.19" />
                    <SPLIT distance="1400" swimtime="00:18:18.95" />
                    <SPLIT distance="1450" swimtime="00:18:58.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="501" reactiontime="+77" swimtime="00:01:12.44" resultid="17770" heatid="19081" lane="6" entrytime="00:01:12.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="500" reactiontime="+84" swimtime="00:10:10.43" resultid="17771" heatid="19096" lane="2" entrytime="00:11:17.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                    <SPLIT distance="100" swimtime="00:01:09.97" />
                    <SPLIT distance="150" swimtime="00:01:47.68" />
                    <SPLIT distance="200" swimtime="00:02:25.66" />
                    <SPLIT distance="250" swimtime="00:03:03.75" />
                    <SPLIT distance="300" swimtime="00:03:42.37" />
                    <SPLIT distance="350" swimtime="00:04:21.36" />
                    <SPLIT distance="400" swimtime="00:05:00.70" />
                    <SPLIT distance="450" swimtime="00:05:39.58" />
                    <SPLIT distance="500" swimtime="00:06:18.58" />
                    <SPLIT distance="550" swimtime="00:06:57.64" />
                    <SPLIT distance="600" swimtime="00:07:36.68" />
                    <SPLIT distance="650" swimtime="00:08:15.30" />
                    <SPLIT distance="700" swimtime="00:08:54.81" />
                    <SPLIT distance="750" swimtime="00:09:33.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" status="DNS" swimtime="00:00:00.00" resultid="19101" heatid="19026" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Damian" lastname="Błaszczyk" birthdate="2006-04-25" gender="M" nation="POL" license="101703700084" swrid="5014987" athleteid="17835">
              <RESULTS>
                <RESULT eventid="1071" points="524" reactiontime="+67" swimtime="00:00:32.18" resultid="17836" heatid="18969" lane="9" />
                <RESULT eventid="1079" points="474" reactiontime="+74" swimtime="00:01:03.47" resultid="17837" heatid="18981" lane="0" entrytime="00:01:03.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="493" reactiontime="+65" swimtime="00:00:28.18" resultid="17838" heatid="19024" lane="7" entrytime="00:00:28.19" entrycourse="LCM" />
                <RESULT eventid="1137" points="475" reactiontime="+68" swimtime="00:01:12.87" resultid="17839" heatid="19047" lane="8" entrytime="00:01:14.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="503" reactiontime="+73" swimtime="00:00:58.95" resultid="17840" heatid="19075" lane="7" entrytime="00:00:59.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.27" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K11 - Pływak wykonał nierównoczesne lub naprzemienne ruchy nóg" eventid="1179" reactiontime="+74" status="DSQ" swimtime="00:02:45.76" resultid="17841" heatid="19092" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                    <SPLIT distance="100" swimtime="00:01:17.18" />
                    <SPLIT distance="150" swimtime="00:02:01.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maksymilian" lastname="Pawlos" birthdate="2007-10-20" gender="M" nation="POL" license="101703700096" swrid="5193083" athleteid="17857">
              <RESULTS>
                <RESULT eventid="1079" points="340" reactiontime="+75" swimtime="00:01:10.87" resultid="17858" heatid="18980" lane="0" entrytime="00:01:11.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="339" reactiontime="+92" swimtime="00:02:40.43" resultid="17859" heatid="18996" lane="3" entrytime="00:02:51.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                    <SPLIT distance="100" swimtime="00:01:18.95" />
                    <SPLIT distance="150" swimtime="00:02:00.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="367" reactiontime="+72" swimtime="00:00:31.10" resultid="17860" heatid="19022" lane="4" entrytime="00:00:31.89" entrycourse="LCM" />
                <RESULT eventid="1121" points="336" reactiontime="+87" swimtime="00:00:34.50" resultid="17861" heatid="19035" lane="4" entrytime="00:00:36.17" entrycourse="LCM" />
                <RESULT eventid="1155" points="256" reactiontime="+75" swimtime="00:02:54.37" resultid="17862" heatid="19058" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.13" />
                    <SPLIT distance="100" swimtime="00:01:23.97" />
                    <SPLIT distance="150" swimtime="00:02:10.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="339" reactiontime="+83" swimtime="00:01:14.30" resultid="17863" heatid="19087" lane="0" entrytime="00:01:13.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Konrad" lastname="Szendała" birthdate="2009-08-09" gender="M" nation="POL" license="101703700128" swrid="5158167" athleteid="17814">
              <RESULTS>
                <RESULT eventid="1063" points="145" reactiontime="+64" swimtime="00:00:39.79" resultid="17815" heatid="18955" lane="3" entrytime="00:00:38.57" entrycourse="LCM" />
                <RESULT eventid="1071" points="128" swimtime="00:00:51.36" resultid="17816" heatid="18970" lane="9" entrytime="00:00:52.21" entrycourse="LCM" />
                <RESULT eventid="1121" points="127" reactiontime="+69" swimtime="00:00:47.65" resultid="17817" heatid="19034" lane="1" entrytime="00:00:47.55" entrycourse="LCM" />
                <RESULT eventid="1137" points="116" swimtime="00:01:56.44" resultid="17818" heatid="19044" lane="8" entrytime="00:01:53.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="116" swimtime="00:01:36.07" resultid="17819" heatid="19069" lane="9" entrytime="00:01:32.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="108" reactiontime="+79" swimtime="00:01:48.61" resultid="17820" heatid="19085" lane="0" entrytime="00:01:42.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Grasza" birthdate="2009-05-29" gender="M" nation="POL" license="101703700132" swrid="5225171" athleteid="17793">
              <RESULTS>
                <RESULT eventid="1063" points="262" reactiontime="+81" swimtime="00:00:32.64" resultid="17794" heatid="18957" lane="1" entrytime="00:00:33.85" entrycourse="LCM" />
                <RESULT eventid="1071" points="244" reactiontime="+81" swimtime="00:00:41.52" resultid="17795" heatid="18971" lane="4" entrytime="00:00:41.82" entrycourse="LCM" />
                <RESULT eventid="1137" points="231" reactiontime="+72" swimtime="00:01:32.65" resultid="17796" heatid="19045" lane="1" entrytime="00:01:36.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="193" reactiontime="+79" swimtime="00:03:16.96" resultid="17797" heatid="19053" lane="0" entrytime="00:03:08.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.65" />
                    <SPLIT distance="100" swimtime="00:01:39.68" />
                    <SPLIT distance="150" swimtime="00:02:34.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" status="DNS" swimtime="00:00:00.00" resultid="17798" heatid="19071" lane="6" entrytime="00:01:14.55" entrycourse="LCM" />
                <RESULT eventid="1179" points="227" reactiontime="+82" swimtime="00:03:26.48" resultid="17799" heatid="19093" lane="7" entrytime="00:03:24.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.39" />
                    <SPLIT distance="100" swimtime="00:01:40.11" />
                    <SPLIT distance="150" swimtime="00:02:35.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Kowalik" birthdate="2009-08-29" gender="M" nation="POL" license="101703700131" swrid="5199338" athleteid="17871">
              <RESULTS>
                <RESULT eventid="1087" points="135" reactiontime="+67" swimtime="00:03:18.81" resultid="17872" heatid="18986" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.49" />
                    <SPLIT distance="100" swimtime="00:01:31.66" />
                    <SPLIT distance="150" swimtime="00:02:26.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="154" reactiontime="+65" swimtime="00:03:28.66" resultid="17873" heatid="18996" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.37" />
                    <SPLIT distance="100" swimtime="00:01:42.36" />
                    <SPLIT distance="150" swimtime="00:02:37.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="137" reactiontime="+70" swimtime="00:00:46.52" resultid="17874" heatid="19034" lane="6" entrytime="00:00:44.99" entrycourse="LCM" />
                <RESULT eventid="1137" points="133" reactiontime="+67" swimtime="00:01:51.39" resultid="17875" heatid="19043" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="136" reactiontime="+76" swimtime="00:01:31.05" resultid="17876" heatid="19069" lane="2" entrytime="00:01:25.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="129" reactiontime="+68" swimtime="00:01:42.37" resultid="17877" heatid="19085" lane="7" entrytime="00:01:38.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03903" nation="POL" region="03" clubid="17213" name="KS Narwal Międzyrzec Podl.">
          <ATHLETES>
            <ATHLETE firstname="Filip" lastname="Pocztarski" birthdate="2008-01-20" gender="M" nation="POL" license="103903700004" swrid="5255452" athleteid="17234">
              <RESULTS>
                <RESULT eventid="1063" points="441" reactiontime="+62" swimtime="00:00:27.46" resultid="17235" heatid="18961" lane="0" entrytime="00:00:27.06" entrycourse="LCM" />
                <RESULT eventid="1087" points="349" reactiontime="+67" swimtime="00:02:24.79" resultid="17236" heatid="18990" lane="8" entrytime="00:02:20.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                    <SPLIT distance="100" swimtime="00:01:10.30" />
                    <SPLIT distance="150" swimtime="00:01:49.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="270" reactiontime="+54" swimtime="00:00:34.44" resultid="17237" heatid="19022" lane="9" entrytime="00:00:36.95" entrycourse="LCM" />
                <RESULT eventid="1121" points="314" reactiontime="+72" swimtime="00:00:35.28" resultid="17238" heatid="19036" lane="9" entrytime="00:00:34.49" entrycourse="LCM" />
                <RESULT eventid="1163" points="427" reactiontime="+69" swimtime="00:01:02.27" resultid="17239" heatid="19074" lane="6" entrytime="00:01:01.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="272" reactiontime="+70" swimtime="00:01:19.93" resultid="17240" heatid="19086" lane="6" entrytime="00:01:18.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Jakimiak" birthdate="2003-04-15" gender="M" nation="POL" license="103903700010" swrid="4931187" athleteid="17221">
              <RESULTS>
                <RESULT eventid="1063" points="669" reactiontime="+63" swimtime="00:00:23.90" resultid="17222" heatid="18962" lane="4" entrytime="00:00:23.38" entrycourse="LCM" />
                <RESULT eventid="1087" points="722" reactiontime="+64" swimtime="00:01:53.66" resultid="17223" heatid="18991" lane="4" entrytime="00:01:53.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.51" />
                    <SPLIT distance="100" swimtime="00:00:56.67" />
                    <SPLIT distance="150" swimtime="00:01:25.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="736" reactiontime="+69" swimtime="00:04:03.67" resultid="17224" heatid="19012" lane="3" entrytime="00:04:08.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.78" />
                    <SPLIT distance="100" swimtime="00:00:59.62" />
                    <SPLIT distance="150" swimtime="00:01:30.95" />
                    <SPLIT distance="200" swimtime="00:02:02.13" />
                    <SPLIT distance="250" swimtime="00:02:33.24" />
                    <SPLIT distance="300" swimtime="00:03:04.48" />
                    <SPLIT distance="350" swimtime="00:03:35.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="620" reactiontime="+67" swimtime="00:00:26.11" resultid="17225" heatid="19025" lane="5" entrytime="00:00:25.80" entrycourse="LCM" />
                <RESULT eventid="1163" points="741" reactiontime="+63" swimtime="00:00:51.82" resultid="17226" heatid="19077" lane="4" entrytime="00:00:52.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cezary" lastname="Cap" birthdate="2007-03-14" gender="M" nation="POL" license="103903700003" swrid="5200026" athleteid="17214">
              <RESULTS>
                <RESULT eventid="1063" points="469" reactiontime="+60" swimtime="00:00:26.91" resultid="17215" heatid="18961" lane="9" entrytime="00:00:27.56" entrycourse="LCM" />
                <RESULT eventid="1087" points="348" reactiontime="+76" swimtime="00:02:24.89" resultid="17216" heatid="18989" lane="3" entrytime="00:02:28.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                    <SPLIT distance="100" swimtime="00:01:08.49" />
                    <SPLIT distance="150" swimtime="00:01:48.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="331" reactiontime="+78" swimtime="00:05:17.86" resultid="17217" heatid="19009" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.15" />
                    <SPLIT distance="100" swimtime="00:01:13.70" />
                    <SPLIT distance="150" swimtime="00:01:53.91" />
                    <SPLIT distance="200" swimtime="00:02:36.01" />
                    <SPLIT distance="250" swimtime="00:03:17.01" />
                    <SPLIT distance="300" swimtime="00:03:59.13" />
                    <SPLIT distance="350" swimtime="00:04:40.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="410" reactiontime="+74" swimtime="00:00:32.28" resultid="17218" heatid="19036" lane="2" entrytime="00:00:33.58" entrycourse="LCM" />
                <RESULT eventid="1163" points="460" reactiontime="+71" swimtime="00:01:00.74" resultid="17219" heatid="19074" lane="1" entrytime="00:01:02.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="296" reactiontime="+74" swimtime="00:01:17.74" resultid="17220" heatid="19086" lane="3" entrytime="00:01:15.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Mironiuk" birthdate="2007-07-06" gender="M" nation="POL" license="103903700002" swrid="5255413" athleteid="17248">
              <RESULTS>
                <RESULT eventid="1063" points="446" reactiontime="+61" swimtime="00:00:27.36" resultid="17249" heatid="18960" lane="5" entrytime="00:00:28.20" entrycourse="LCM" />
                <RESULT eventid="1095" points="391" reactiontime="+61" swimtime="00:02:32.96" resultid="17250" heatid="18997" lane="0" entrytime="00:02:35.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.91" />
                    <SPLIT distance="150" swimtime="00:01:55.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="386" reactiontime="+53" swimtime="00:00:30.57" resultid="17251" heatid="19019" lane="2" />
                <RESULT eventid="1121" points="481" reactiontime="+65" swimtime="00:00:30.63" resultid="17252" heatid="19037" lane="7" entrytime="00:00:30.35" entrycourse="LCM" />
                <RESULT eventid="1163" status="DNS" swimtime="00:00:00.00" resultid="17253" heatid="19073" lane="0" entrytime="00:01:07.56" entrycourse="LCM" />
                <RESULT eventid="1171" points="437" reactiontime="+62" swimtime="00:01:08.30" resultid="17254" heatid="19088" lane="0" entrytime="00:01:08.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Franciszek" lastname="Korulczyk" birthdate="2006-12-11" gender="M" nation="POL" license="103903700025" swrid="5165778" athleteid="17227">
              <RESULTS>
                <RESULT eventid="1063" points="495" reactiontime="+58" swimtime="00:00:26.43" resultid="17228" heatid="18962" lane="0" entrytime="00:00:25.93" entrycourse="LCM" />
                <RESULT eventid="1079" points="436" reactiontime="+62" swimtime="00:01:05.24" resultid="17229" heatid="18980" lane="6" entrytime="00:01:06.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="442" reactiontime="+62" swimtime="00:00:29.22" resultid="17230" heatid="19020" lane="6" />
                <RESULT eventid="1121" points="458" reactiontime="+62" swimtime="00:00:31.12" resultid="17231" heatid="19037" lane="6" entrytime="00:00:30.10" entrycourse="LCM" />
                <RESULT eventid="1163" points="522" reactiontime="+59" swimtime="00:00:58.23" resultid="17232" heatid="19075" lane="4" entrytime="00:00:58.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="400" reactiontime="+64" swimtime="00:01:10.35" resultid="17233" heatid="19087" lane="6" entrytime="00:01:12.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Morgunowicz" birthdate="2008-09-05" gender="M" nation="POL" license="103903700030" swrid="5429176" athleteid="17241">
              <RESULTS>
                <RESULT eventid="1063" points="270" reactiontime="+59" swimtime="00:00:32.32" resultid="17242" heatid="18958" lane="2" entrytime="00:00:32.03" entrycourse="LCM" />
                <RESULT eventid="1071" points="198" reactiontime="+63" swimtime="00:00:44.45" resultid="17243" heatid="18970" lane="4" entrytime="00:00:46.16" entrycourse="LCM" />
                <RESULT eventid="1121" points="181" reactiontime="+84" swimtime="00:00:42.36" resultid="17244" heatid="19035" lane="1" entrytime="00:00:40.29" entrycourse="LCM" />
                <RESULT eventid="1137" points="168" reactiontime="+73" swimtime="00:01:42.90" resultid="17245" heatid="19043" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="260" reactiontime="+66" swimtime="00:01:13.41" resultid="17246" heatid="19072" lane="8" entrytime="00:01:12.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="156" reactiontime="+79" swimtime="00:01:36.25" resultid="17247" heatid="19085" lane="6" entrytime="00:01:35.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="07614" nation="POL" region="14" clubid="18457" name="UKS GOS Raszyn">
          <ATHLETES>
            <ATHLETE firstname="Julia" lastname="Kulik" birthdate="2005-02-11" gender="F" nation="POL" license="107614600014" swrid="5083156" athleteid="18464">
              <RESULTS>
                <RESULT eventid="1059" points="653" reactiontime="+70" status="EXH" swimtime="00:00:27.28" resultid="18465" heatid="18951" lane="6" entrytime="00:00:27.10" entrycourse="LCM" />
                <RESULT eventid="1083" points="674" reactiontime="+71" status="EXH" swimtime="00:02:08.85" resultid="18466" heatid="18985" lane="5" entrytime="00:02:03.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.63" />
                    <SPLIT distance="100" swimtime="00:01:02.98" />
                    <SPLIT distance="150" swimtime="00:01:35.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="643" reactiontime="+75" status="EXH" swimtime="00:04:33.90" resultid="18467" heatid="19007" lane="5" entrytime="00:04:21.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.37" />
                    <SPLIT distance="100" swimtime="00:01:04.10" />
                    <SPLIT distance="150" swimtime="00:01:38.92" />
                    <SPLIT distance="200" swimtime="00:02:14.06" />
                    <SPLIT distance="250" swimtime="00:02:48.91" />
                    <SPLIT distance="300" swimtime="00:03:24.58" />
                    <SPLIT distance="350" swimtime="00:03:59.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="682" reactiontime="+70" status="EXH" swimtime="00:00:58.73" resultid="18468" heatid="19066" lane="5" entrytime="00:00:56.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="663" reactiontime="+75" status="EXH" swimtime="00:09:15.82" resultid="18469" heatid="19097" lane="5" entrytime="00:09:22.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                    <SPLIT distance="100" swimtime="00:01:06.02" />
                    <SPLIT distance="150" swimtime="00:01:40.34" />
                    <SPLIT distance="200" swimtime="00:02:15.18" />
                    <SPLIT distance="250" swimtime="00:02:50.27" />
                    <SPLIT distance="300" swimtime="00:03:25.19" />
                    <SPLIT distance="350" swimtime="00:04:00.03" />
                    <SPLIT distance="400" swimtime="00:04:35.40" />
                    <SPLIT distance="450" swimtime="00:05:10.32" />
                    <SPLIT distance="500" swimtime="00:05:45.68" />
                    <SPLIT distance="550" swimtime="00:06:21.20" />
                    <SPLIT distance="600" swimtime="00:06:56.97" />
                    <SPLIT distance="650" swimtime="00:07:31.31" />
                    <SPLIT distance="700" swimtime="00:08:06.57" />
                    <SPLIT distance="750" swimtime="00:08:41.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Owerko" birthdate="2002-09-02" gender="F" nation="POL" license="107614600016" swrid="5106999" athleteid="18470">
              <RESULTS>
                <RESULT eventid="1067" points="601" reactiontime="+67" status="EXH" swimtime="00:00:34.83" resultid="18471" heatid="18967" lane="7" entrytime="00:00:35.45" entrycourse="LCM" />
                <RESULT eventid="1133" points="497" reactiontime="+64" status="EXH" swimtime="00:01:20.95" resultid="18472" heatid="19041" lane="2" entrytime="00:01:18.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="442" reactiontime="+71" status="EXH" swimtime="00:03:02.60" resultid="18473" heatid="19091" lane="8" entrytime="00:02:57.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.96" />
                    <SPLIT distance="100" swimtime="00:01:28.95" />
                    <SPLIT distance="150" swimtime="00:02:16.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Polańska" birthdate="2000-09-24" gender="F" nation="POL" license="107614600027" swrid="4585041" athleteid="18458">
              <RESULTS>
                <RESULT eventid="1059" points="711" reactiontime="+72" status="EXH" swimtime="00:00:26.52" resultid="18459" heatid="18951" lane="4" entrytime="00:00:26.22" entrycourse="LCM" />
                <RESULT eventid="1083" points="793" reactiontime="+76" status="EXH" swimtime="00:02:02.02" resultid="18460" heatid="18985" lane="4" entrytime="00:01:59.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.28" />
                    <SPLIT distance="100" swimtime="00:00:59.21" />
                    <SPLIT distance="150" swimtime="00:01:30.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="730" reactiontime="+74" status="EXH" swimtime="00:04:22.61" resultid="18461" heatid="19007" lane="4" entrytime="00:04:15.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.35" />
                    <SPLIT distance="100" swimtime="00:01:01.85" />
                    <SPLIT distance="150" swimtime="00:01:35.03" />
                    <SPLIT distance="200" swimtime="00:02:08.16" />
                    <SPLIT distance="250" swimtime="00:02:41.48" />
                    <SPLIT distance="300" swimtime="00:03:15.24" />
                    <SPLIT distance="350" swimtime="00:03:49.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="773" reactiontime="+71" status="EXH" swimtime="00:00:56.32" resultid="18462" heatid="19066" lane="4" entrytime="00:00:55.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="750" reactiontime="+77" status="EXH" swimtime="00:08:53.54" resultid="18463" heatid="19097" lane="4" entrytime="00:08:53.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.53" />
                    <SPLIT distance="100" swimtime="00:01:04.26" />
                    <SPLIT distance="150" swimtime="00:01:38.34" />
                    <SPLIT distance="200" swimtime="00:02:12.56" />
                    <SPLIT distance="250" swimtime="00:02:46.41" />
                    <SPLIT distance="300" swimtime="00:03:20.06" />
                    <SPLIT distance="350" swimtime="00:03:53.74" />
                    <SPLIT distance="400" swimtime="00:04:27.22" />
                    <SPLIT distance="450" swimtime="00:05:00.88" />
                    <SPLIT distance="500" swimtime="00:05:34.51" />
                    <SPLIT distance="550" swimtime="00:06:08.28" />
                    <SPLIT distance="600" swimtime="00:06:42.01" />
                    <SPLIT distance="650" swimtime="00:07:15.16" />
                    <SPLIT distance="700" swimtime="00:07:48.23" />
                    <SPLIT distance="750" swimtime="00:08:21.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00605" nation="POL" region="05" clubid="18572" name="UKS SP-149 Łódź">
          <ATHLETES>
            <ATHLETE firstname="Nina" lastname="Ostrowska" birthdate="2006-02-25" gender="F" nation="POL" license="100605600295" swrid="5025337" athleteid="18573">
              <RESULTS>
                <RESULT eventid="6361" status="DNS" swimtime="00:00:00.00" resultid="18574" heatid="19055" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03103" nation="POL" region="03" clubid="17255" name="KU AZS UMCS Lublin">
          <ATHLETES>
            <ATHLETE firstname="Kamil" lastname="Chycki" birthdate="2005-03-17" gender="M" nation="POL" license="103103700179" swrid="5228586" athleteid="17398">
              <RESULTS>
                <RESULT eventid="1063" points="473" reactiontime="+73" swimtime="00:00:26.83" resultid="17399" heatid="18961" lane="6" entrytime="00:00:26.64" entrycourse="LCM" />
                <RESULT eventid="1087" points="534" reactiontime="+75" swimtime="00:02:05.67" resultid="17400" heatid="18991" lane="0" entrytime="00:02:04.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.78" />
                    <SPLIT distance="100" swimtime="00:01:01.41" />
                    <SPLIT distance="150" swimtime="00:01:34.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="508" reactiontime="+71" swimtime="00:04:35.74" resultid="17401" heatid="19011" lane="1" entrytime="00:04:33.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.32" />
                    <SPLIT distance="100" swimtime="00:01:04.57" />
                    <SPLIT distance="150" swimtime="00:01:39.48" />
                    <SPLIT distance="200" swimtime="00:02:14.54" />
                    <SPLIT distance="250" swimtime="00:02:50.66" />
                    <SPLIT distance="300" swimtime="00:03:26.30" />
                    <SPLIT distance="350" swimtime="00:04:02.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="554" reactiontime="+73" swimtime="00:00:57.09" resultid="17402" heatid="19076" lane="5" entrytime="00:00:56.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Burdyn" birthdate="2005-03-06" gender="F" nation="POL" license="103103600116" swrid="5066543" athleteid="17443">
              <RESULTS>
                <RESULT eventid="1075" points="607" reactiontime="+70" swimtime="00:01:05.52" resultid="17444" heatid="18977" lane="3" entrytime="00:01:05.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="564" reactiontime="+66" swimtime="00:02:16.67" resultid="17445" heatid="18984" lane="3" entrytime="00:02:15.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.90" />
                    <SPLIT distance="100" swimtime="00:01:06.84" />
                    <SPLIT distance="150" swimtime="00:01:42.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="562" reactiontime="+69" swimtime="00:04:46.39" resultid="17446" heatid="19007" lane="0" entrytime="00:04:43.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.92" />
                    <SPLIT distance="100" swimtime="00:01:07.40" />
                    <SPLIT distance="150" swimtime="00:01:43.57" />
                    <SPLIT distance="200" swimtime="00:02:20.47" />
                    <SPLIT distance="250" swimtime="00:02:57.80" />
                    <SPLIT distance="300" swimtime="00:03:34.51" />
                    <SPLIT distance="350" swimtime="00:04:11.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="565" reactiontime="+66" swimtime="00:02:32.52" resultid="17447" heatid="19050" lane="7" entrytime="00:02:31.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.96" />
                    <SPLIT distance="100" swimtime="00:01:10.66" />
                    <SPLIT distance="150" swimtime="00:01:57.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1150" points="490" reactiontime="+67" swimtime="00:02:34.48" resultid="17448" heatid="19057" lane="5" entrytime="00:02:30.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.88" />
                    <SPLIT distance="100" swimtime="00:01:12.40" />
                    <SPLIT distance="150" swimtime="00:01:53.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="536" reactiontime="+71" swimtime="00:09:56.69" resultid="17449" heatid="19095" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.88" />
                    <SPLIT distance="100" swimtime="00:01:10.48" />
                    <SPLIT distance="150" swimtime="00:01:47.81" />
                    <SPLIT distance="200" swimtime="00:02:24.89" />
                    <SPLIT distance="250" swimtime="00:03:02.00" />
                    <SPLIT distance="300" swimtime="00:03:39.13" />
                    <SPLIT distance="350" swimtime="00:04:16.92" />
                    <SPLIT distance="400" swimtime="00:04:54.76" />
                    <SPLIT distance="450" swimtime="00:05:32.84" />
                    <SPLIT distance="500" swimtime="00:06:11.03" />
                    <SPLIT distance="550" swimtime="00:06:49.10" />
                    <SPLIT distance="600" swimtime="00:07:27.11" />
                    <SPLIT distance="650" swimtime="00:08:05.35" />
                    <SPLIT distance="700" swimtime="00:08:43.30" />
                    <SPLIT distance="750" swimtime="00:09:20.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Mróz" birthdate="2003-05-27" gender="M" nation="POL" license="103103700118" swrid="4744845" athleteid="17477">
              <RESULTS>
                <RESULT eventid="1079" points="578" reactiontime="+73" swimtime="00:00:59.41" resultid="17478" heatid="18981" lane="6" entrytime="00:00:59.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6365" points="662" reactiontime="+74" swimtime="00:08:38.53" resultid="17479" heatid="19003" lane="3" entrytime="00:08:36.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                    <SPLIT distance="100" swimtime="00:01:01.39" />
                    <SPLIT distance="150" swimtime="00:01:33.81" />
                    <SPLIT distance="200" swimtime="00:02:06.44" />
                    <SPLIT distance="250" swimtime="00:02:39.07" />
                    <SPLIT distance="300" swimtime="00:03:11.81" />
                    <SPLIT distance="350" swimtime="00:03:44.31" />
                    <SPLIT distance="400" swimtime="00:04:17.16" />
                    <SPLIT distance="450" swimtime="00:04:49.36" />
                    <SPLIT distance="500" swimtime="00:05:22.22" />
                    <SPLIT distance="550" swimtime="00:05:54.86" />
                    <SPLIT distance="600" swimtime="00:06:27.74" />
                    <SPLIT distance="650" swimtime="00:07:00.39" />
                    <SPLIT distance="700" swimtime="00:07:33.38" />
                    <SPLIT distance="750" swimtime="00:08:06.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="601" reactiontime="+70" swimtime="00:04:20.74" resultid="17480" heatid="19012" lane="7" entrytime="00:04:14.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.21" />
                    <SPLIT distance="100" swimtime="00:01:01.77" />
                    <SPLIT distance="150" swimtime="00:01:35.41" />
                    <SPLIT distance="200" swimtime="00:02:08.93" />
                    <SPLIT distance="250" swimtime="00:02:42.17" />
                    <SPLIT distance="300" swimtime="00:03:15.44" />
                    <SPLIT distance="350" swimtime="00:03:48.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="554" reactiontime="+75" swimtime="00:02:18.79" resultid="17481" heatid="19054" lane="2" entrytime="00:02:19.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.30" />
                    <SPLIT distance="100" swimtime="00:01:06.18" />
                    <SPLIT distance="150" swimtime="00:01:46.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="626" reactiontime="+79" swimtime="00:02:09.44" resultid="17482" heatid="19059" lane="4" entrytime="00:02:04.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.56" />
                    <SPLIT distance="100" swimtime="00:01:01.93" />
                    <SPLIT distance="150" swimtime="00:01:36.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Błażej" lastname="Fronczek" birthdate="2009-07-31" gender="M" nation="POL" license="103103700087" swrid="5225188" athleteid="17367">
              <RESULTS>
                <RESULT eventid="1063" points="220" reactiontime="+68" swimtime="00:00:34.60" resultid="17368" heatid="18954" lane="4" entrytime="00:00:41.44" entrycourse="LCM" />
                <RESULT eventid="1095" points="244" reactiontime="+68" swimtime="00:02:58.91" resultid="17369" heatid="18996" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.07" />
                    <SPLIT distance="100" swimtime="00:01:26.78" />
                    <SPLIT distance="150" swimtime="00:02:14.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="244" reactiontime="+68" swimtime="00:05:52.06" resultid="17370" heatid="19008" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.33" />
                    <SPLIT distance="100" swimtime="00:01:21.96" />
                    <SPLIT distance="150" swimtime="00:02:08.48" />
                    <SPLIT distance="200" swimtime="00:02:55.17" />
                    <SPLIT distance="250" swimtime="00:03:40.66" />
                    <SPLIT distance="300" swimtime="00:04:26.43" />
                    <SPLIT distance="350" swimtime="00:05:10.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="236" reactiontime="+67" swimtime="00:00:38.82" resultid="17371" heatid="19035" lane="9" entrytime="00:00:43.25" entrycourse="LCM" />
                <RESULT eventid="1163" points="207" reactiontime="+60" swimtime="00:01:19.21" resultid="17372" heatid="19070" lane="5" entrytime="00:01:16.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Norbert" lastname="Zacharzyński" birthdate="2003-06-06" gender="M" nation="POL" license="103103700158" swrid="4837459" athleteid="17430">
              <RESULTS>
                <RESULT eventid="1071" points="676" reactiontime="+65" swimtime="00:00:29.56" resultid="17431" heatid="18974" lane="5" entrytime="00:00:29.85" entrycourse="LCM" />
                <RESULT eventid="1113" points="581" reactiontime="+64" swimtime="00:00:26.68" resultid="17432" heatid="19025" lane="6" entrytime="00:00:26.42" entrycourse="LCM" />
                <RESULT eventid="1137" points="664" reactiontime="+65" swimtime="00:01:05.19" resultid="17433" heatid="19047" lane="4" entrytime="00:01:05.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="671" reactiontime="+67" swimtime="00:02:10.21" resultid="17434" heatid="19054" lane="4" entrytime="00:02:08.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.99" />
                    <SPLIT distance="100" swimtime="00:01:03.39" />
                    <SPLIT distance="150" swimtime="00:01:40.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="679" reactiontime="+68" swimtime="00:02:23.47" resultid="17435" heatid="19094" lane="4" entrytime="00:02:21.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.73" />
                    <SPLIT distance="100" swimtime="00:01:10.01" />
                    <SPLIT distance="150" swimtime="00:01:47.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alicja" lastname="Pyszniak" birthdate="2005-02-05" gender="F" nation="POL" license="103103600154" swrid="4973772" athleteid="17276">
              <RESULTS>
                <RESULT eventid="1059" points="473" reactiontime="+71" swimtime="00:00:30.36" resultid="17277" heatid="18949" lane="4" entrytime="00:00:30.50" entrycourse="LCM" />
                <RESULT eventid="1083" points="511" reactiontime="+74" swimtime="00:02:21.26" resultid="17278" heatid="18984" lane="2" entrytime="00:02:19.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                    <SPLIT distance="100" swimtime="00:01:08.16" />
                    <SPLIT distance="150" swimtime="00:01:45.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="498" reactiontime="+76" swimtime="00:04:58.23" resultid="17279" heatid="19006" lane="3" entrytime="00:04:55.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                    <SPLIT distance="100" swimtime="00:01:10.22" />
                    <SPLIT distance="150" swimtime="00:01:47.68" />
                    <SPLIT distance="200" swimtime="00:02:25.55" />
                    <SPLIT distance="250" swimtime="00:03:03.53" />
                    <SPLIT distance="300" swimtime="00:03:41.68" />
                    <SPLIT distance="350" swimtime="00:04:20.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="504" reactiontime="+71" swimtime="00:01:04.94" resultid="17280" heatid="19065" lane="8" entrytime="00:01:05.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="495" reactiontime="+75" swimtime="00:10:12.70" resultid="17281" heatid="19095" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                    <SPLIT distance="100" swimtime="00:01:12.53" />
                    <SPLIT distance="150" swimtime="00:01:50.83" />
                    <SPLIT distance="200" swimtime="00:02:29.09" />
                    <SPLIT distance="250" swimtime="00:03:07.54" />
                    <SPLIT distance="300" swimtime="00:03:45.86" />
                    <SPLIT distance="350" swimtime="00:04:24.19" />
                    <SPLIT distance="400" swimtime="00:05:02.67" />
                    <SPLIT distance="450" swimtime="00:05:41.42" />
                    <SPLIT distance="500" swimtime="00:06:20.28" />
                    <SPLIT distance="550" swimtime="00:06:59.60" />
                    <SPLIT distance="600" swimtime="00:07:38.89" />
                    <SPLIT distance="650" swimtime="00:08:17.55" />
                    <SPLIT distance="700" swimtime="00:08:56.88" />
                    <SPLIT distance="750" swimtime="00:09:35.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Łoboda" birthdate="2002-11-04" gender="M" nation="POL" license="103103700098" swrid="5083376" athleteid="17335">
              <RESULTS>
                <RESULT eventid="1063" points="640" reactiontime="+70" swimtime="00:00:24.26" resultid="17336" heatid="18962" lane="5" entrytime="00:00:24.17" entrycourse="LCM" />
                <RESULT eventid="1079" points="660" reactiontime="+68" swimtime="00:00:56.83" resultid="17337" heatid="18981" lane="4" entrytime="00:00:56.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="666" reactiontime="+65" swimtime="00:00:25.49" resultid="17338" heatid="19025" lane="4" entrytime="00:00:25.10" entrycourse="LCM" />
                <RESULT eventid="1121" points="551" reactiontime="+80" swimtime="00:00:29.26" resultid="17339" heatid="19037" lane="4" entrytime="00:00:29.09" entrycourse="LCM" />
                <RESULT eventid="1163" points="585" reactiontime="+64" swimtime="00:00:56.08" resultid="17340" heatid="19077" lane="8" entrytime="00:00:55.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Cioch-Gradzik" birthdate="2003-07-12" gender="F" nation="POL" license="103103600114" swrid="4809210" athleteid="17456">
              <RESULTS>
                <RESULT eventid="1075" points="576" reactiontime="+75" swimtime="00:01:06.65" resultid="17457" heatid="18977" lane="2" entrytime="00:01:06.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="545" reactiontime="+81" swimtime="00:02:18.25" resultid="17458" heatid="18985" lane="1" entrytime="00:02:12.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                    <SPLIT distance="100" swimtime="00:01:07.58" />
                    <SPLIT distance="150" swimtime="00:01:43.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="498" reactiontime="+86" swimtime="00:04:58.12" resultid="17459" heatid="19007" lane="6" entrytime="00:04:36.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.00" />
                    <SPLIT distance="100" swimtime="00:01:11.29" />
                    <SPLIT distance="150" swimtime="00:01:49.53" />
                    <SPLIT distance="200" swimtime="00:02:27.54" />
                    <SPLIT distance="250" swimtime="00:03:04.47" />
                    <SPLIT distance="300" swimtime="00:03:42.30" />
                    <SPLIT distance="350" swimtime="00:04:20.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Śledź" birthdate="2005-10-27" gender="M" nation="POL" license="103103700193" swrid="4931032" athleteid="17392">
              <RESULTS>
                <RESULT eventid="1087" points="518" reactiontime="+61" swimtime="00:02:06.96" resultid="17394" heatid="18990" lane="4" entrytime="00:02:07.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.87" />
                    <SPLIT distance="100" swimtime="00:01:01.43" />
                    <SPLIT distance="150" swimtime="00:01:34.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6365" points="511" reactiontime="+61" swimtime="00:09:25.35" resultid="17395" heatid="19002" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                    <SPLIT distance="100" swimtime="00:01:08.00" />
                    <SPLIT distance="150" swimtime="00:01:44.52" />
                    <SPLIT distance="200" swimtime="00:02:20.83" />
                    <SPLIT distance="250" swimtime="00:02:57.46" />
                    <SPLIT distance="300" swimtime="00:03:33.50" />
                    <SPLIT distance="350" swimtime="00:04:09.48" />
                    <SPLIT distance="400" swimtime="00:04:45.15" />
                    <SPLIT distance="450" swimtime="00:05:21.20" />
                    <SPLIT distance="500" swimtime="00:05:56.95" />
                    <SPLIT distance="550" swimtime="00:06:32.89" />
                    <SPLIT distance="600" swimtime="00:07:08.22" />
                    <SPLIT distance="650" swimtime="00:07:43.73" />
                    <SPLIT distance="700" swimtime="00:08:19.04" />
                    <SPLIT distance="750" swimtime="00:08:52.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="573" reactiontime="+65" swimtime="00:04:24.94" resultid="17396" heatid="19011" lane="5" entrytime="00:04:27.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.77" />
                    <SPLIT distance="100" swimtime="00:01:02.77" />
                    <SPLIT distance="150" swimtime="00:01:37.00" />
                    <SPLIT distance="200" swimtime="00:02:11.05" />
                    <SPLIT distance="250" swimtime="00:02:45.42" />
                    <SPLIT distance="300" swimtime="00:03:19.77" />
                    <SPLIT distance="350" swimtime="00:03:54.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="502" reactiontime="+48" swimtime="00:00:58.99" resultid="17397" heatid="19067" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martyna" lastname="Piesko" birthdate="2003-05-13" gender="F" nation="POL" license="103103600119" swrid="4621520" athleteid="17301">
              <RESULTS>
                <RESULT eventid="1059" points="635" reactiontime="+62" swimtime="00:00:27.53" resultid="17302" heatid="18951" lane="2" entrytime="00:00:27.44" entrycourse="LCM" />
                <RESULT eventid="1091" points="652" reactiontime="+63" swimtime="00:02:22.19" resultid="17303" heatid="18994" lane="5" entrytime="00:02:24.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                    <SPLIT distance="100" swimtime="00:01:09.39" />
                    <SPLIT distance="150" swimtime="00:01:46.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kinga" lastname="Żydek" birthdate="2005-12-06" gender="F" nation="POL" license="103103600180" swrid="5109094" athleteid="17407">
              <RESULTS>
                <RESULT eventid="1067" points="569" reactiontime="+69" swimtime="00:00:35.46" resultid="17408" heatid="18967" lane="1" entrytime="00:00:35.84" entrycourse="LCM" />
                <RESULT eventid="1133" points="593" reactiontime="+62" swimtime="00:01:16.32" resultid="17409" heatid="19041" lane="5" entrytime="00:01:17.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="509" reactiontime="+66" swimtime="00:02:37.87" resultid="17410" heatid="19049" lane="5" entrytime="00:02:42.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.75" />
                    <SPLIT distance="100" swimtime="00:01:19.22" />
                    <SPLIT distance="150" swimtime="00:02:01.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="633" reactiontime="+66" swimtime="00:02:42.01" resultid="17411" heatid="19091" lane="5" entrytime="00:02:45.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                    <SPLIT distance="100" swimtime="00:01:20.35" />
                    <SPLIT distance="150" swimtime="00:02:01.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="420" reactiontime="+76" swimtime="00:10:47.22" resultid="17412" heatid="19096" lane="4" entrytime="00:10:38.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                    <SPLIT distance="100" swimtime="00:01:15.39" />
                    <SPLIT distance="150" swimtime="00:01:57.08" />
                    <SPLIT distance="200" swimtime="00:02:37.51" />
                    <SPLIT distance="250" swimtime="00:03:17.30" />
                    <SPLIT distance="300" swimtime="00:03:57.94" />
                    <SPLIT distance="350" swimtime="00:04:39.07" />
                    <SPLIT distance="400" swimtime="00:05:18.91" />
                    <SPLIT distance="450" swimtime="00:06:00.21" />
                    <SPLIT distance="500" swimtime="00:06:41.34" />
                    <SPLIT distance="550" swimtime="00:07:23.79" />
                    <SPLIT distance="600" swimtime="00:08:04.17" />
                    <SPLIT distance="650" swimtime="00:08:46.07" />
                    <SPLIT distance="700" swimtime="00:09:26.75" />
                    <SPLIT distance="750" swimtime="00:10:07.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Chodulski" birthdate="2000-03-06" gender="M" nation="POL" license="103103700073" swrid="4395632" athleteid="17491">
              <RESULTS>
                <RESULT eventid="1087" points="676" reactiontime="+65" swimtime="00:01:56.19" resultid="17492" heatid="18991" lane="5" entrytime="00:01:55.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.56" />
                    <SPLIT distance="100" swimtime="00:00:56.92" />
                    <SPLIT distance="150" swimtime="00:01:26.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6365" points="689" reactiontime="+66" swimtime="00:08:31.86" resultid="17493" heatid="19003" lane="4" entrytime="00:08:21.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.19" />
                    <SPLIT distance="100" swimtime="00:01:01.07" />
                    <SPLIT distance="150" swimtime="00:01:33.52" />
                    <SPLIT distance="200" swimtime="00:02:05.65" />
                    <SPLIT distance="250" swimtime="00:02:38.35" />
                    <SPLIT distance="300" swimtime="00:03:10.87" />
                    <SPLIT distance="350" swimtime="00:03:43.48" />
                    <SPLIT distance="400" swimtime="00:04:15.98" />
                    <SPLIT distance="450" swimtime="00:04:48.33" />
                    <SPLIT distance="500" swimtime="00:05:20.53" />
                    <SPLIT distance="550" swimtime="00:05:53.09" />
                    <SPLIT distance="600" swimtime="00:06:25.28" />
                    <SPLIT distance="650" swimtime="00:06:57.20" />
                    <SPLIT distance="700" swimtime="00:07:28.90" />
                    <SPLIT distance="750" swimtime="00:08:00.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="730" reactiontime="+65" swimtime="00:04:04.37" resultid="17494" heatid="19012" lane="4" entrytime="00:04:00.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.24" />
                    <SPLIT distance="100" swimtime="00:00:58.75" />
                    <SPLIT distance="150" swimtime="00:01:29.67" />
                    <SPLIT distance="200" swimtime="00:02:00.89" />
                    <SPLIT distance="250" swimtime="00:02:31.90" />
                    <SPLIT distance="300" swimtime="00:03:03.03" />
                    <SPLIT distance="350" swimtime="00:03:34.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="597" reactiontime="+68" swimtime="00:00:55.71" resultid="17495" heatid="19077" lane="6" entrytime="00:00:53.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="734" reactiontime="+68" swimtime="00:16:05.37" resultid="17496" heatid="19100" lane="4" entrytime="00:16:03.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.82" />
                    <SPLIT distance="100" swimtime="00:01:00.13" />
                    <SPLIT distance="150" swimtime="00:01:32.02" />
                    <SPLIT distance="200" swimtime="00:02:04.05" />
                    <SPLIT distance="250" swimtime="00:02:36.57" />
                    <SPLIT distance="300" swimtime="00:03:08.71" />
                    <SPLIT distance="350" swimtime="00:03:40.73" />
                    <SPLIT distance="400" swimtime="00:04:13.05" />
                    <SPLIT distance="450" swimtime="00:04:45.47" />
                    <SPLIT distance="500" swimtime="00:05:18.25" />
                    <SPLIT distance="550" swimtime="00:05:50.52" />
                    <SPLIT distance="600" swimtime="00:06:23.13" />
                    <SPLIT distance="650" swimtime="00:06:55.69" />
                    <SPLIT distance="700" swimtime="00:07:28.26" />
                    <SPLIT distance="750" swimtime="00:08:00.61" />
                    <SPLIT distance="800" swimtime="00:08:33.10" />
                    <SPLIT distance="850" swimtime="00:09:05.35" />
                    <SPLIT distance="900" swimtime="00:09:37.78" />
                    <SPLIT distance="950" swimtime="00:10:10.20" />
                    <SPLIT distance="1000" swimtime="00:10:42.69" />
                    <SPLIT distance="1050" swimtime="00:11:15.24" />
                    <SPLIT distance="1100" swimtime="00:11:47.92" />
                    <SPLIT distance="1150" swimtime="00:12:20.33" />
                    <SPLIT distance="1200" swimtime="00:12:52.96" />
                    <SPLIT distance="1250" swimtime="00:13:25.64" />
                    <SPLIT distance="1300" swimtime="00:13:58.18" />
                    <SPLIT distance="1350" swimtime="00:14:30.60" />
                    <SPLIT distance="1400" swimtime="00:15:02.78" />
                    <SPLIT distance="1450" swimtime="00:15:34.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henry" lastname="Radzikowski" birthdate="2002-01-16" gender="M" nation="POL" license="103103700176" swrid="5378200" athleteid="17341">
              <RESULTS>
                <RESULT eventid="1063" points="633" reactiontime="+68" swimtime="00:00:24.35" resultid="17342" heatid="18953" lane="5" />
                <RESULT eventid="1087" points="679" reactiontime="+68" swimtime="00:01:56.03" resultid="17343" heatid="18991" lane="3" entrytime="00:01:55.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.59" />
                    <SPLIT distance="100" swimtime="00:00:55.19" />
                    <SPLIT distance="150" swimtime="00:01:25.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6365" points="632" reactiontime="+72" swimtime="00:08:46.71" resultid="17344" heatid="19003" lane="5" entrytime="00:08:30.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                    <SPLIT distance="100" swimtime="00:01:01.28" />
                    <SPLIT distance="150" swimtime="00:01:33.74" />
                    <SPLIT distance="200" swimtime="00:02:06.29" />
                    <SPLIT distance="250" swimtime="00:02:38.94" />
                    <SPLIT distance="300" swimtime="00:03:12.05" />
                    <SPLIT distance="350" swimtime="00:03:45.14" />
                    <SPLIT distance="400" swimtime="00:04:18.31" />
                    <SPLIT distance="450" swimtime="00:04:51.45" />
                    <SPLIT distance="500" swimtime="00:05:25.13" />
                    <SPLIT distance="550" swimtime="00:05:58.74" />
                    <SPLIT distance="600" swimtime="00:06:33.10" />
                    <SPLIT distance="650" swimtime="00:07:06.86" />
                    <SPLIT distance="700" swimtime="00:07:41.16" />
                    <SPLIT distance="750" swimtime="00:08:14.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="720" reactiontime="+70" swimtime="00:04:05.52" resultid="17345" heatid="19012" lane="5" entrytime="00:04:06.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.09" />
                    <SPLIT distance="100" swimtime="00:00:58.92" />
                    <SPLIT distance="150" swimtime="00:01:29.93" />
                    <SPLIT distance="200" swimtime="00:02:01.08" />
                    <SPLIT distance="250" swimtime="00:02:32.04" />
                    <SPLIT distance="300" swimtime="00:03:03.18" />
                    <SPLIT distance="350" swimtime="00:03:34.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="683" reactiontime="+66" swimtime="00:00:53.26" resultid="17346" heatid="19077" lane="3" entrytime="00:00:53.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Wiśniewska" birthdate="2004-10-23" gender="F" nation="POL" license="103103600133" swrid="5172971" athleteid="17282">
              <RESULTS>
                <RESULT eventid="1059" points="571" reactiontime="+64" swimtime="00:00:28.52" resultid="17283" heatid="18951" lane="0" entrytime="00:00:28.12" entrycourse="LCM" />
                <RESULT eventid="1083" points="606" reactiontime="+80" swimtime="00:02:13.45" resultid="17284" heatid="18984" lane="5" entrytime="00:02:14.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.06" />
                    <SPLIT distance="100" swimtime="00:01:04.67" />
                    <SPLIT distance="150" swimtime="00:01:39.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="631" reactiontime="+64" swimtime="00:00:31.45" resultid="17285" heatid="19030" lane="3" entrytime="00:00:31.25" entrycourse="LCM" />
                <RESULT eventid="1141" points="555" reactiontime="+88" swimtime="00:02:33.39" resultid="17286" heatid="19048" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.06" />
                    <SPLIT distance="100" swimtime="00:01:10.22" />
                    <SPLIT distance="150" swimtime="00:01:57.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="629" reactiontime="+65" swimtime="00:01:07.16" resultid="17287" heatid="19082" lane="3" entrytime="00:01:07.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="495" reactiontime="+84" swimtime="00:10:12.48" resultid="17288" heatid="19095" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                    <SPLIT distance="100" swimtime="00:01:10.76" />
                    <SPLIT distance="150" swimtime="00:01:48.54" />
                    <SPLIT distance="200" swimtime="00:02:26.14" />
                    <SPLIT distance="250" swimtime="00:03:04.28" />
                    <SPLIT distance="300" swimtime="00:03:42.42" />
                    <SPLIT distance="350" swimtime="00:04:21.32" />
                    <SPLIT distance="400" swimtime="00:05:00.20" />
                    <SPLIT distance="450" swimtime="00:05:39.41" />
                    <SPLIT distance="500" swimtime="00:06:18.65" />
                    <SPLIT distance="550" swimtime="00:06:58.05" />
                    <SPLIT distance="600" swimtime="00:07:36.93" />
                    <SPLIT distance="650" swimtime="00:08:16.38" />
                    <SPLIT distance="700" swimtime="00:08:55.18" />
                    <SPLIT distance="750" swimtime="00:09:34.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Kafarska" birthdate="2009-06-28" gender="F" nation="POL" license="103103600105" swrid="5243531" athleteid="18619">
              <RESULTS>
                <RESULT eventid="1059" points="325" reactiontime="+72" swimtime="00:00:34.41" resultid="18620" heatid="18946" lane="1" />
                <RESULT eventid="1091" points="245" reactiontime="+69" status="EXH" swimtime="00:03:17.09" resultid="19109" heatid="18992" lane="7" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.02" />
                    <SPLIT distance="100" swimtime="00:01:39.86" />
                    <SPLIT distance="150" swimtime="00:02:31.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Sławacki" birthdate="2005-01-04" gender="M" nation="POL" license="103103700159" swrid="4780103" athleteid="17379">
              <RESULTS>
                <RESULT eventid="1063" points="627" reactiontime="+70" swimtime="00:00:24.42" resultid="17380" heatid="18962" lane="3" entrytime="00:00:24.22" entrycourse="LCM" />
                <RESULT eventid="1087" points="674" reactiontime="+71" swimtime="00:01:56.28" resultid="17381" heatid="18991" lane="6" entrytime="00:01:55.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.68" />
                    <SPLIT distance="100" swimtime="00:00:57.46" />
                    <SPLIT distance="150" swimtime="00:01:27.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="685" reactiontime="+71" swimtime="00:04:09.62" resultid="17382" heatid="19012" lane="6" entrytime="00:04:11.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.96" />
                    <SPLIT distance="100" swimtime="00:00:58.97" />
                    <SPLIT distance="150" swimtime="00:01:30.44" />
                    <SPLIT distance="200" swimtime="00:02:02.11" />
                    <SPLIT distance="250" swimtime="00:02:34.41" />
                    <SPLIT distance="300" swimtime="00:03:06.40" />
                    <SPLIT distance="350" swimtime="00:03:38.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="639" reactiontime="+71" swimtime="00:02:12.35" resultid="17383" heatid="19054" lane="5" entrytime="00:02:11.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.23" />
                    <SPLIT distance="100" swimtime="00:01:03.15" />
                    <SPLIT distance="150" swimtime="00:01:41.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="685" reactiontime="+70" swimtime="00:00:53.21" resultid="17384" heatid="19077" lane="5" entrytime="00:00:53.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Karwowska" birthdate="2004-09-08" gender="F" nation="POL" license="103103600223" swrid="5019889" athleteid="17269">
              <RESULTS>
                <RESULT eventid="1059" points="572" reactiontime="+67" swimtime="00:00:28.50" resultid="17270" heatid="18951" lane="9" entrytime="00:00:28.47" entrycourse="LCM" />
                <RESULT eventid="1083" points="589" reactiontime="+83" swimtime="00:02:14.76" resultid="17271" heatid="18985" lane="7" entrytime="00:02:12.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                    <SPLIT distance="100" swimtime="00:01:05.39" />
                    <SPLIT distance="150" swimtime="00:01:40.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="572" reactiontime="+85" swimtime="00:04:44.71" resultid="17272" heatid="19007" lane="7" entrytime="00:04:39.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                    <SPLIT distance="100" swimtime="00:01:06.73" />
                    <SPLIT distance="150" swimtime="00:01:43.10" />
                    <SPLIT distance="200" swimtime="00:02:18.72" />
                    <SPLIT distance="250" swimtime="00:02:55.27" />
                    <SPLIT distance="300" swimtime="00:03:32.22" />
                    <SPLIT distance="350" swimtime="00:04:08.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="598" reactiontime="+73" swimtime="00:00:32.01" resultid="17273" heatid="19030" lane="7" entrytime="00:00:32.25" entrycourse="LCM" />
                <RESULT eventid="1159" points="568" reactiontime="+80" swimtime="00:01:02.43" resultid="17274" heatid="19066" lane="8" entrytime="00:01:01.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="542" reactiontime="+82" swimtime="00:09:54.32" resultid="17275" heatid="19095" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.00" />
                    <SPLIT distance="100" swimtime="00:01:10.42" />
                    <SPLIT distance="150" swimtime="00:01:48.13" />
                    <SPLIT distance="200" swimtime="00:02:25.60" />
                    <SPLIT distance="250" swimtime="00:03:03.51" />
                    <SPLIT distance="300" swimtime="00:03:41.43" />
                    <SPLIT distance="350" swimtime="00:04:19.52" />
                    <SPLIT distance="400" swimtime="00:04:57.52" />
                    <SPLIT distance="450" swimtime="00:05:35.46" />
                    <SPLIT distance="500" swimtime="00:06:13.20" />
                    <SPLIT distance="550" swimtime="00:06:50.73" />
                    <SPLIT distance="600" swimtime="00:07:28.16" />
                    <SPLIT distance="650" swimtime="00:08:05.31" />
                    <SPLIT distance="700" swimtime="00:08:42.27" />
                    <SPLIT distance="750" swimtime="00:09:18.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="571" reactiontime="+75" status="EXH" swimtime="00:01:09.39" resultid="19114" heatid="19082" lane="4" entrytime="00:01:13.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Weronika" lastname="Żmuda" birthdate="2000-03-26" gender="F" nation="POL" license="103103600005" swrid="4353669" athleteid="17403">
              <RESULTS>
                <RESULT eventid="1067" points="699" reactiontime="+65" swimtime="00:00:33.12" resultid="17404" heatid="18967" lane="4" entrytime="00:00:33.14" entrycourse="LCM" />
                <RESULT eventid="1075" points="610" reactiontime="+69" swimtime="00:01:05.41" resultid="17405" heatid="18977" lane="4" entrytime="00:01:04.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="651" reactiontime="+66" swimtime="00:01:13.98" resultid="17406" heatid="19041" lane="4" entrytime="00:01:13.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Lewtak" birthdate="2004-05-20" gender="M" nation="POL" license="103103700131" swrid="5056726" athleteid="17467">
              <RESULTS>
                <RESULT eventid="1079" points="479" reactiontime="+65" swimtime="00:01:03.23" resultid="17468" heatid="18981" lane="9" entrytime="00:01:03.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="430" reactiontime="+73" swimtime="00:00:29.49" resultid="17469" heatid="19023" lane="3" entrytime="00:00:29.91" entrycourse="LCM" />
                <RESULT eventid="1155" points="497" reactiontime="+70" swimtime="00:02:19.70" resultid="17470" heatid="19059" lane="2" entrytime="00:02:19.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.27" />
                    <SPLIT distance="100" swimtime="00:01:06.97" />
                    <SPLIT distance="150" swimtime="00:01:43.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Kowalska" birthdate="2005-11-14" gender="F" nation="POL" license="103103600177" swrid="4931027" athleteid="17484">
              <RESULTS>
                <RESULT eventid="1083" points="586" reactiontime="+72" swimtime="00:02:14.99" resultid="17485" heatid="18985" lane="9" entrytime="00:02:14.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                    <SPLIT distance="100" swimtime="00:01:05.19" />
                    <SPLIT distance="150" swimtime="00:01:40.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="526" reactiontime="+73" swimtime="00:05:29.77" resultid="17486" heatid="18999" lane="6" entrytime="00:05:14.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                    <SPLIT distance="100" swimtime="00:01:15.31" />
                    <SPLIT distance="150" swimtime="00:01:58.14" />
                    <SPLIT distance="200" swimtime="00:02:39.26" />
                    <SPLIT distance="250" swimtime="00:03:28.29" />
                    <SPLIT distance="300" swimtime="00:04:16.83" />
                    <SPLIT distance="350" swimtime="00:04:53.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="574" reactiontime="+73" swimtime="00:04:44.48" resultid="17487" heatid="19006" lane="5" entrytime="00:04:48.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                    <SPLIT distance="100" swimtime="00:01:08.38" />
                    <SPLIT distance="150" swimtime="00:01:44.83" />
                    <SPLIT distance="200" swimtime="00:02:21.31" />
                    <SPLIT distance="250" swimtime="00:02:57.70" />
                    <SPLIT distance="300" swimtime="00:03:33.78" />
                    <SPLIT distance="350" swimtime="00:04:09.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="542" reactiontime="+71" swimtime="00:02:34.68" resultid="17488" heatid="19050" lane="9" entrytime="00:02:34.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                    <SPLIT distance="100" swimtime="00:01:14.83" />
                    <SPLIT distance="150" swimtime="00:01:58.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="551" reactiontime="+71" swimtime="00:01:03.07" resultid="17489" heatid="19066" lane="9" entrytime="00:01:02.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="582" reactiontime="+61" swimtime="00:09:40.36" resultid="17490" heatid="19095" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.78" />
                    <SPLIT distance="100" swimtime="00:01:10.70" />
                    <SPLIT distance="150" swimtime="00:01:47.55" />
                    <SPLIT distance="200" swimtime="00:02:24.47" />
                    <SPLIT distance="250" swimtime="00:03:01.39" />
                    <SPLIT distance="300" swimtime="00:03:38.30" />
                    <SPLIT distance="350" swimtime="00:04:15.07" />
                    <SPLIT distance="400" swimtime="00:04:51.78" />
                    <SPLIT distance="450" swimtime="00:05:28.34" />
                    <SPLIT distance="500" swimtime="00:06:04.88" />
                    <SPLIT distance="550" swimtime="00:06:41.41" />
                    <SPLIT distance="600" swimtime="00:07:17.88" />
                    <SPLIT distance="650" swimtime="00:07:54.31" />
                    <SPLIT distance="700" swimtime="00:08:30.19" />
                    <SPLIT distance="750" swimtime="00:09:05.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Dragan" birthdate="2008-12-26" gender="M" nation="POL" license="103103700078" swrid="5009209" athleteid="17360">
              <RESULTS>
                <RESULT eventid="1063" points="253" swimtime="00:00:33.05" resultid="17361" heatid="18957" lane="2" entrytime="00:00:33.64" entrycourse="LCM" />
                <RESULT eventid="1071" points="175" swimtime="00:00:46.36" resultid="17362" heatid="18971" lane="0" entrytime="00:00:44.92" entrycourse="LCM" />
                <RESULT eventid="1137" points="167" swimtime="00:01:43.09" resultid="17363" heatid="19045" lane="9" entrytime="00:01:38.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="185" swimtime="00:03:19.92" resultid="17364" heatid="19051" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.09" />
                    <SPLIT distance="100" swimtime="00:01:38.19" />
                    <SPLIT distance="150" swimtime="00:02:36.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="259" reactiontime="+73" swimtime="00:01:13.53" resultid="17365" heatid="19070" lane="4" entrytime="00:01:16.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="221" swimtime="00:03:28.50" resultid="17366" heatid="19093" lane="8" entrytime="00:03:26.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.83" />
                    <SPLIT distance="100" swimtime="00:01:42.01" />
                    <SPLIT distance="150" swimtime="00:02:35.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nikodem" lastname="Chołżyński" birthdate="2003-03-30" gender="M" nation="POL" license="103103700124" swrid="4744862" athleteid="17463">
              <RESULTS>
                <RESULT eventid="1079" points="555" reactiontime="+63" swimtime="00:01:00.20" resultid="17464" heatid="18981" lane="8" entrytime="00:01:01.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="517" reactiontime="+66" swimtime="00:00:27.73" resultid="17465" heatid="19024" lane="3" entrytime="00:00:27.72" entrycourse="LCM" />
                <RESULT eventid="1163" points="515" reactiontime="+69" swimtime="00:00:58.52" resultid="17466" heatid="19075" lane="1" entrytime="00:00:59.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Iga" lastname="Banach" birthdate="2008-06-04" gender="F" nation="POL" license="103103600081" swrid="5286984" athleteid="17317">
              <RESULTS>
                <RESULT eventid="1059" points="318" swimtime="00:00:34.65" resultid="17318" heatid="18948" lane="2" entrytime="00:00:33.75" entrycourse="LCM" />
                <RESULT eventid="1067" points="310" reactiontime="+61" swimtime="00:00:43.41" resultid="17319" heatid="18966" lane="0" entrytime="00:00:42.69" entrycourse="LCM" />
                <RESULT eventid="1108" points="260" reactiontime="+72" swimtime="00:00:38.23" resultid="17320" heatid="19015" lane="1" entrytime="00:00:39.08" entrycourse="LCM" />
                <RESULT comment="K4 - Pływak wykonał cykl ruchowy inny niż jeden ruch ramion i jedno kopnięcie nogami (z wyjątkiem ostatniego cyklu przed nawrotem lub zakończeniem wyścigu)" eventid="1133" reactiontime="+77" status="DSQ" swimtime="00:01:36.26" resultid="17321" heatid="19040" lane="0" entrytime="00:01:37.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="333" reactiontime="+77" swimtime="00:01:14.58" resultid="17322" heatid="19062" lane="5" entrytime="00:01:18.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="298" reactiontime="+86" swimtime="00:03:28.25" resultid="19110" heatid="19090" lane="0" entrytime="00:03:55.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.76" />
                    <SPLIT distance="100" swimtime="00:01:39.90" />
                    <SPLIT distance="150" swimtime="00:02:35.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Sagan" birthdate="2002-10-14" gender="M" nation="POL" license="103103700110" swrid="4440789" athleteid="17426">
              <RESULTS>
                <RESULT eventid="1071" points="677" reactiontime="+63" swimtime="00:00:29.55" resultid="17427" heatid="18974" lane="4" entrytime="00:00:29.65" entrycourse="LCM" />
                <RESULT eventid="1137" points="640" reactiontime="+65" swimtime="00:01:05.99" resultid="17428" heatid="19047" lane="5" entrytime="00:01:05.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="629" reactiontime="+56" swimtime="00:01:00.51" resultid="17429" heatid="19088" lane="6" entrytime="00:01:02.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emilia" lastname="Łuszczewska" birthdate="2005-05-07" gender="F" nation="POL" license="103103600184" swrid="5164146" athleteid="17497">
              <RESULTS>
                <RESULT eventid="1091" points="512" reactiontime="+62" swimtime="00:02:34.11" resultid="17498" heatid="18994" lane="7" entrytime="00:02:31.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.60" />
                    <SPLIT distance="100" swimtime="00:01:16.10" />
                    <SPLIT distance="150" swimtime="00:01:55.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="521" reactiontime="+61" swimtime="00:00:33.51" resultid="17499" heatid="19030" lane="8" entrytime="00:00:32.72" entrycourse="LCM" />
                <RESULT eventid="1141" points="510" reactiontime="+69" swimtime="00:02:37.81" resultid="17500" heatid="19050" lane="1" entrytime="00:02:32.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                    <SPLIT distance="100" swimtime="00:01:15.24" />
                    <SPLIT distance="150" swimtime="00:02:03.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="486" reactiontime="+62" swimtime="00:01:13.18" resultid="17501" heatid="19082" lane="0" entrytime="00:01:09.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Dwojak" birthdate="2004-05-28" gender="F" nation="POL" license="103103600132" swrid="4910045" athleteid="17256">
              <RESULTS>
                <RESULT eventid="1059" points="682" reactiontime="+71" swimtime="00:00:26.89" resultid="17257" heatid="18951" lane="3" entrytime="00:00:26.93" entrycourse="LCM" />
                <RESULT eventid="1067" points="652" reactiontime="+71" swimtime="00:00:33.89" resultid="17258" heatid="18967" lane="5" entrytime="00:00:33.64" entrycourse="LCM" />
                <RESULT eventid="1108" points="545" reactiontime="+69" swimtime="00:00:29.90" resultid="17259" heatid="19014" lane="1" />
                <RESULT eventid="1141" points="655" reactiontime="+70" swimtime="00:02:25.16" resultid="17260" heatid="19050" lane="5" entrytime="00:02:23.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.21" />
                    <SPLIT distance="100" swimtime="00:01:10.47" />
                    <SPLIT distance="150" swimtime="00:01:51.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="656" reactiontime="+75" swimtime="00:00:59.50" resultid="17261" heatid="19066" lane="2" entrytime="00:00:59.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="591" reactiontime="+71" swimtime="00:09:37.55" resultid="17262" heatid="19095" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                    <SPLIT distance="100" swimtime="00:01:09.52" />
                    <SPLIT distance="150" swimtime="00:01:46.65" />
                    <SPLIT distance="200" swimtime="00:02:23.87" />
                    <SPLIT distance="250" swimtime="00:03:00.83" />
                    <SPLIT distance="300" swimtime="00:03:37.60" />
                    <SPLIT distance="350" swimtime="00:04:14.67" />
                    <SPLIT distance="400" swimtime="00:04:51.19" />
                    <SPLIT distance="450" swimtime="00:05:27.53" />
                    <SPLIT distance="500" swimtime="00:06:04.05" />
                    <SPLIT distance="550" swimtime="00:06:40.97" />
                    <SPLIT distance="600" swimtime="00:07:17.28" />
                    <SPLIT distance="650" swimtime="00:07:53.89" />
                    <SPLIT distance="700" swimtime="00:08:28.93" />
                    <SPLIT distance="750" swimtime="00:09:03.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kornelia" lastname="Samuła" birthdate="2003-10-25" gender="F" nation="POL" license="103103600121" swrid="4744827" athleteid="17295">
              <RESULTS>
                <RESULT eventid="1059" points="482" reactiontime="+74" swimtime="00:00:30.18" resultid="17296" heatid="18950" lane="6" entrytime="00:00:29.54" entrycourse="LCM" />
                <RESULT eventid="1091" points="546" reactiontime="+67" swimtime="00:02:30.88" resultid="17297" heatid="18994" lane="6" entrytime="00:02:28.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                    <SPLIT distance="100" swimtime="00:01:12.89" />
                    <SPLIT distance="150" swimtime="00:01:52.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="571" reactiontime="+73" swimtime="00:00:32.52" resultid="17298" heatid="19030" lane="1" entrytime="00:00:32.66" entrycourse="LCM" />
                <RESULT eventid="1141" points="467" reactiontime="+75" swimtime="00:02:42.49" resultid="17299" heatid="19048" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                    <SPLIT distance="100" swimtime="00:01:13.77" />
                    <SPLIT distance="150" swimtime="00:02:03.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="518" reactiontime="+66" swimtime="00:01:11.66" resultid="17300" heatid="19082" lane="1" entrytime="00:01:09.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mikołaj" lastname="Kubiniec" birthdate="2004-08-29" gender="M" nation="POL" license="103103700128" swrid="5109071" athleteid="17385">
              <RESULTS>
                <RESULT eventid="1063" points="544" reactiontime="+65" swimtime="00:00:25.61" resultid="17386" heatid="18962" lane="7" entrytime="00:00:25.58" entrycourse="LCM" />
                <RESULT eventid="1079" points="410" reactiontime="+65" swimtime="00:01:06.60" resultid="17387" heatid="18979" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1087" points="545" reactiontime="+66" swimtime="00:02:04.82" resultid="17388" heatid="18991" lane="7" entrytime="00:02:01.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.75" />
                    <SPLIT distance="100" swimtime="00:00:59.81" />
                    <SPLIT distance="150" swimtime="00:01:32.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6365" points="572" reactiontime="+64" swimtime="00:09:04.45" resultid="17389" heatid="19003" lane="6" entrytime="00:08:58.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.45" />
                    <SPLIT distance="100" swimtime="00:01:02.97" />
                    <SPLIT distance="150" swimtime="00:01:38.09" />
                    <SPLIT distance="200" swimtime="00:02:13.36" />
                    <SPLIT distance="250" swimtime="00:02:48.19" />
                    <SPLIT distance="300" swimtime="00:03:22.79" />
                    <SPLIT distance="350" swimtime="00:03:57.59" />
                    <SPLIT distance="400" swimtime="00:04:32.77" />
                    <SPLIT distance="450" swimtime="00:05:06.58" />
                    <SPLIT distance="500" swimtime="00:05:41.08" />
                    <SPLIT distance="550" swimtime="00:06:15.15" />
                    <SPLIT distance="600" swimtime="00:06:48.68" />
                    <SPLIT distance="650" swimtime="00:07:22.23" />
                    <SPLIT distance="700" swimtime="00:07:56.43" />
                    <SPLIT distance="750" swimtime="00:08:30.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="574" reactiontime="+64" swimtime="00:04:24.69" resultid="17390" heatid="19012" lane="1" entrytime="00:04:18.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.85" />
                    <SPLIT distance="100" swimtime="00:00:59.50" />
                    <SPLIT distance="150" swimtime="00:01:32.87" />
                    <SPLIT distance="200" swimtime="00:02:07.70" />
                    <SPLIT distance="250" swimtime="00:02:42.20" />
                    <SPLIT distance="300" swimtime="00:03:16.75" />
                    <SPLIT distance="350" swimtime="00:03:51.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="570" reactiontime="+64" swimtime="00:00:56.57" resultid="17391" heatid="19077" lane="0" entrytime="00:00:55.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Dwojak" birthdate="2004-05-28" gender="F" nation="POL" license="103103600137" swrid="4910044" athleteid="17263">
              <RESULTS>
                <RESULT eventid="1059" points="602" reactiontime="+78" swimtime="00:00:28.03" resultid="17264" heatid="18951" lane="8" entrytime="00:00:28.10" entrycourse="LCM" />
                <RESULT eventid="1091" points="622" reactiontime="+93" swimtime="00:02:24.46" resultid="17265" heatid="18994" lane="4" entrytime="00:02:23.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.00" />
                    <SPLIT distance="100" swimtime="00:01:10.81" />
                    <SPLIT distance="150" swimtime="00:01:48.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="594" reactiontime="+83" swimtime="00:04:41.16" resultid="17266" heatid="19007" lane="9" entrytime="00:04:43.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.75" />
                    <SPLIT distance="100" swimtime="00:01:06.91" />
                    <SPLIT distance="150" swimtime="00:01:42.91" />
                    <SPLIT distance="200" swimtime="00:02:18.76" />
                    <SPLIT distance="250" swimtime="00:02:54.92" />
                    <SPLIT distance="300" swimtime="00:03:30.99" />
                    <SPLIT distance="350" swimtime="00:04:06.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="605" reactiontime="+64" swimtime="00:01:08.05" resultid="17267" heatid="19082" lane="6" entrytime="00:01:08.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="575" reactiontime="+81" swimtime="00:09:42.89" resultid="17268" heatid="19095" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.63" />
                    <SPLIT distance="100" swimtime="00:01:09.69" />
                    <SPLIT distance="150" swimtime="00:01:46.93" />
                    <SPLIT distance="200" swimtime="00:02:23.85" />
                    <SPLIT distance="250" swimtime="00:03:00.86" />
                    <SPLIT distance="300" swimtime="00:03:37.66" />
                    <SPLIT distance="350" swimtime="00:04:14.37" />
                    <SPLIT distance="400" swimtime="00:04:51.41" />
                    <SPLIT distance="450" swimtime="00:05:28.02" />
                    <SPLIT distance="500" swimtime="00:06:04.59" />
                    <SPLIT distance="550" swimtime="00:06:41.57" />
                    <SPLIT distance="600" swimtime="00:07:18.27" />
                    <SPLIT distance="650" swimtime="00:07:55.04" />
                    <SPLIT distance="700" swimtime="00:08:31.69" />
                    <SPLIT distance="750" swimtime="00:09:08.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Kozak" birthdate="2004-08-19" gender="F" nation="POL" license="103103600122" swrid="4892188" athleteid="17450">
              <RESULTS>
                <RESULT eventid="1075" points="510" reactiontime="+67" swimtime="00:01:09.44" resultid="17451" heatid="18977" lane="8" entrytime="00:01:09.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="501" reactiontime="+73" swimtime="00:02:22.25" resultid="17452" heatid="18984" lane="6" entrytime="00:02:15.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                    <SPLIT distance="100" swimtime="00:01:07.84" />
                    <SPLIT distance="150" swimtime="00:01:45.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="485" reactiontime="+74" swimtime="00:00:31.09" resultid="17453" heatid="19017" lane="8" entrytime="00:00:30.69" entrycourse="LCM" />
                <RESULT comment="G1 - Pływak nie złamał powierzchni wody głową przed lub na linii 15 m po starcie lub nawrocie" eventid="1117" reactiontime="+58" status="DSQ" swimtime="00:00:33.77" resultid="17454" heatid="19029" lane="3" entrytime="00:00:33.13" entrycourse="LCM" />
                <RESULT eventid="1150" points="517" reactiontime="+73" swimtime="00:02:31.75" resultid="17455" heatid="19057" lane="3" entrytime="00:02:33.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                    <SPLIT distance="100" swimtime="00:01:12.09" />
                    <SPLIT distance="150" swimtime="00:01:52.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Adamczyk" birthdate="2003-02-16" gender="M" nation="POL" license="103103700117" swrid="4621512" athleteid="17419">
              <RESULTS>
                <RESULT eventid="1071" points="527" reactiontime="+62" swimtime="00:00:32.11" resultid="17420" heatid="18969" lane="2" />
                <RESULT eventid="1087" points="545" reactiontime="+66" swimtime="00:02:04.84" resultid="17421" heatid="18991" lane="2" entrytime="00:01:58.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.03" />
                    <SPLIT distance="100" swimtime="00:01:01.11" />
                    <SPLIT distance="150" swimtime="00:01:33.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="645" reactiontime="+62" swimtime="00:04:14.68" resultid="17422" heatid="19012" lane="8" entrytime="00:04:20.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.72" />
                    <SPLIT distance="100" swimtime="00:00:58.25" />
                    <SPLIT distance="150" swimtime="00:01:30.80" />
                    <SPLIT distance="200" swimtime="00:02:03.50" />
                    <SPLIT distance="250" swimtime="00:02:36.75" />
                    <SPLIT distance="300" swimtime="00:03:09.59" />
                    <SPLIT distance="350" swimtime="00:03:42.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1137" points="513" reactiontime="+66" swimtime="00:01:11.05" resultid="17423" heatid="19047" lane="7" entrytime="00:01:12.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="562" reactiontime="+65" swimtime="00:00:56.83" resultid="17424" heatid="19077" lane="2" entrytime="00:00:54.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="553" reactiontime="+72" swimtime="00:02:33.62" resultid="17425" heatid="19094" lane="3" entrytime="00:02:37.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                    <SPLIT distance="100" swimtime="00:01:14.87" />
                    <SPLIT distance="150" swimtime="00:01:54.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Tomaszewski" birthdate="2005-09-16" gender="M" nation="POL" license="103103700178" swrid="4973779" athleteid="17471">
              <RESULTS>
                <RESULT eventid="1079" points="633" reactiontime="+75" swimtime="00:00:57.65" resultid="17472" heatid="18981" lane="5" entrytime="00:00:58.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="602" reactiontime="+75" swimtime="00:04:48.72" resultid="17473" heatid="19001" lane="4" entrytime="00:04:47.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.98" />
                    <SPLIT distance="100" swimtime="00:01:03.69" />
                    <SPLIT distance="150" swimtime="00:01:41.49" />
                    <SPLIT distance="200" swimtime="00:02:18.73" />
                    <SPLIT distance="250" swimtime="00:03:00.39" />
                    <SPLIT distance="300" swimtime="00:03:42.40" />
                    <SPLIT distance="350" swimtime="00:04:16.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="606" reactiontime="+73" swimtime="00:00:26.31" resultid="17474" heatid="19025" lane="2" entrytime="00:00:26.45" entrycourse="LCM" />
                <RESULT eventid="1145" points="602" reactiontime="+76" swimtime="00:02:14.97" resultid="17475" heatid="19054" lane="3" entrytime="00:02:15.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.65" />
                    <SPLIT distance="100" swimtime="00:01:02.72" />
                    <SPLIT distance="150" swimtime="00:01:43.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="670" reactiontime="+70" swimtime="00:00:59.24" resultid="17476" heatid="19088" lane="4" entrytime="00:00:59.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Starkiewicz" birthdate="2009-12-02" gender="F" nation="POL" license="103103600076" swrid="5286992" athleteid="17323">
              <RESULTS>
                <RESULT eventid="1059" points="336" swimtime="00:00:34.04" resultid="17324" heatid="18946" lane="9" />
                <RESULT eventid="1083" points="293" reactiontime="+86" swimtime="00:02:50.04" resultid="17325" heatid="18982" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.88" />
                    <SPLIT distance="100" swimtime="00:01:21.98" />
                    <SPLIT distance="150" swimtime="00:02:08.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="242" reactiontime="+93" swimtime="00:06:19.43" resultid="17326" heatid="19004" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.79" />
                    <SPLIT distance="100" swimtime="00:01:24.71" />
                    <SPLIT distance="150" swimtime="00:02:15.46" />
                    <SPLIT distance="200" swimtime="00:03:06.23" />
                    <SPLIT distance="250" swimtime="00:03:57.56" />
                    <SPLIT distance="300" swimtime="00:04:48.13" />
                    <SPLIT distance="350" swimtime="00:05:37.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="239" reactiontime="+84" swimtime="00:03:23.21" resultid="17327" heatid="19048" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.78" />
                    <SPLIT distance="100" swimtime="00:01:37.71" />
                    <SPLIT distance="150" swimtime="00:02:41.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="280" reactiontime="+83" swimtime="00:01:18.99" resultid="17328" heatid="19062" lane="4" entrytime="00:01:15.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jeremi" lastname="Siuda" birthdate="2008-08-01" gender="M" nation="POL" license="103103700091" swrid="5353688" athleteid="17373">
              <RESULTS>
                <RESULT eventid="1063" points="245" swimtime="00:00:33.38" resultid="17374" heatid="18957" lane="0" entrytime="00:00:34.25" entrycourse="LCM" />
                <RESULT eventid="1071" points="246" reactiontime="+71" swimtime="00:00:41.37" resultid="17375" heatid="18970" lane="3" entrytime="00:00:48.01" entrycourse="LCM" />
                <RESULT eventid="1121" points="179" reactiontime="+76" swimtime="00:00:42.54" resultid="17376" heatid="19033" lane="6" entrytime="00:00:52.24" entrycourse="LCM" />
                <RESULT eventid="1137" points="228" swimtime="00:01:33.07" resultid="17377" heatid="19045" lane="5" entrytime="00:01:34.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="226" reactiontime="+70" swimtime="00:01:16.98" resultid="17378" heatid="19070" lane="3" entrytime="00:01:17.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marika" lastname="Wieczorek" birthdate="2003-05-07" gender="F" nation="POL" license="103103600138" swrid="4947511" athleteid="17314">
              <RESULTS>
                <RESULT eventid="1059" points="504" swimtime="00:00:29.73" resultid="17315" heatid="18945" lane="2" />
                <RESULT eventid="1159" points="510" swimtime="00:01:04.72" resultid="17316" heatid="19061" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Domoradzka" birthdate="2003-07-07" gender="F" nation="POL" license="103103600136" swrid="4907098" athleteid="17308">
              <RESULTS>
                <RESULT eventid="1059" points="520" reactiontime="+69" swimtime="00:00:29.42" resultid="17309" heatid="18950" lane="3" entrytime="00:00:28.91" entrycourse="LCM" />
                <RESULT eventid="1083" points="600" reactiontime="+70" swimtime="00:02:13.93" resultid="17310" heatid="18985" lane="6" entrytime="00:02:11.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.16" />
                    <SPLIT distance="100" swimtime="00:01:05.52" />
                    <SPLIT distance="150" swimtime="00:01:40.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="580" reactiontime="+74" swimtime="00:04:43.47" resultid="17311" heatid="19007" lane="2" entrytime="00:04:37.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                    <SPLIT distance="100" swimtime="00:01:09.03" />
                    <SPLIT distance="150" swimtime="00:01:45.70" />
                    <SPLIT distance="200" swimtime="00:02:22.27" />
                    <SPLIT distance="250" swimtime="00:02:58.24" />
                    <SPLIT distance="300" swimtime="00:03:34.40" />
                    <SPLIT distance="350" swimtime="00:04:09.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="520" reactiontime="+71" swimtime="00:01:04.27" resultid="17312" heatid="19066" lane="0" entrytime="00:01:02.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="578" reactiontime="+73" swimtime="00:09:41.74" resultid="17313" heatid="19095" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                    <SPLIT distance="100" swimtime="00:01:10.70" />
                    <SPLIT distance="150" swimtime="00:01:48.11" />
                    <SPLIT distance="200" swimtime="00:02:25.12" />
                    <SPLIT distance="250" swimtime="00:03:02.05" />
                    <SPLIT distance="300" swimtime="00:03:38.34" />
                    <SPLIT distance="350" swimtime="00:04:15.32" />
                    <SPLIT distance="400" swimtime="00:04:52.09" />
                    <SPLIT distance="450" swimtime="00:05:28.70" />
                    <SPLIT distance="500" swimtime="00:06:05.32" />
                    <SPLIT distance="550" swimtime="00:06:42.24" />
                    <SPLIT distance="600" swimtime="00:07:19.38" />
                    <SPLIT distance="650" swimtime="00:07:56.21" />
                    <SPLIT distance="700" swimtime="00:08:32.20" />
                    <SPLIT distance="750" swimtime="00:09:07.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Skoczylas" birthdate="2009-04-27" gender="M" nation="POL" license="103103700074" swrid="5225165" athleteid="17354">
              <RESULTS>
                <RESULT eventid="1063" points="290" reactiontime="+64" swimtime="00:00:31.59" resultid="17355" heatid="18958" lane="7" entrytime="00:00:32.36" entrycourse="LCM" />
                <RESULT eventid="6365" points="325" reactiontime="+58" swimtime="00:10:57.59" resultid="17356" heatid="19002" lane="7" entrytime="00:11:00.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                    <SPLIT distance="100" swimtime="00:01:17.05" />
                    <SPLIT distance="150" swimtime="00:01:58.79" />
                    <SPLIT distance="200" swimtime="00:02:40.42" />
                    <SPLIT distance="250" swimtime="00:03:22.46" />
                    <SPLIT distance="300" swimtime="00:04:04.94" />
                    <SPLIT distance="350" swimtime="00:04:46.95" />
                    <SPLIT distance="400" swimtime="00:05:29.12" />
                    <SPLIT distance="450" swimtime="00:06:11.46" />
                    <SPLIT distance="500" swimtime="00:06:53.61" />
                    <SPLIT distance="550" swimtime="00:07:35.18" />
                    <SPLIT distance="600" swimtime="00:08:17.15" />
                    <SPLIT distance="650" swimtime="00:08:58.30" />
                    <SPLIT distance="700" swimtime="00:09:38.90" />
                    <SPLIT distance="750" swimtime="00:10:19.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="243" swimtime="00:00:35.66" resultid="17357" heatid="19021" lane="2" entrytime="00:00:39.60" entrycourse="LCM" />
                <RESULT eventid="1145" points="269" reactiontime="+64" swimtime="00:02:56.57" resultid="17358" heatid="19052" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.58" />
                    <SPLIT distance="100" swimtime="00:01:24.86" />
                    <SPLIT distance="150" swimtime="00:02:18.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="168" reactiontime="+64" swimtime="00:03:20.50" resultid="17359" heatid="19058" lane="4" entrytime="00:03:18.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.44" />
                    <SPLIT distance="100" swimtime="00:01:32.66" />
                    <SPLIT distance="150" swimtime="00:02:28.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miłosz" lastname="Fronczek" birthdate="2008-01-31" gender="M" nation="POL" license="103103700086" swrid="5225191" athleteid="17413">
              <RESULTS>
                <RESULT eventid="1071" points="252" reactiontime="+76" swimtime="00:00:41.04" resultid="17414" heatid="18971" lane="3" entrytime="00:00:43.00" entrycourse="LCM" />
                <RESULT eventid="1087" points="344" reactiontime="+63" swimtime="00:02:25.57" resultid="17415" heatid="18990" lane="9" entrytime="00:02:26.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                    <SPLIT distance="100" swimtime="00:01:10.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="355" reactiontime="+76" swimtime="00:05:10.67" resultid="17416" heatid="19009" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                    <SPLIT distance="100" swimtime="00:01:14.93" />
                    <SPLIT distance="150" swimtime="00:01:54.75" />
                    <SPLIT distance="200" swimtime="00:02:34.68" />
                    <SPLIT distance="250" swimtime="00:03:14.88" />
                    <SPLIT distance="300" swimtime="00:03:54.97" />
                    <SPLIT distance="350" swimtime="00:04:33.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="290" reactiontime="+69" swimtime="00:00:36.25" resultid="17417" heatid="19032" lane="5" />
                <RESULT eventid="1163" points="331" swimtime="00:01:07.78" resultid="17418" heatid="19072" lane="5" entrytime="00:01:09.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Sobolewski" birthdate="2008-07-13" gender="M" nation="POL" license="103103700084" swrid="5340910" athleteid="17347">
              <RESULTS>
                <RESULT eventid="1063" points="145" swimtime="00:00:39.78" resultid="17348" heatid="18955" lane="0" entrytime="00:00:40.46" entrycourse="LCM" />
                <RESULT eventid="1071" points="126" reactiontime="+92" swimtime="00:00:51.73" resultid="17349" heatid="18969" lane="4" entrytime="00:00:53.11" entrycourse="LCM" />
                <RESULT eventid="1121" points="117" reactiontime="+75" swimtime="00:00:49.04" resultid="17350" heatid="19033" lane="5" entrytime="00:00:50.75" entrycourse="LCM" />
                <RESULT eventid="1137" points="121" reactiontime="+82" swimtime="00:01:54.72" resultid="17351" heatid="19043" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="133" reactiontime="+65" swimtime="00:01:31.74" resultid="17352" heatid="19069" lane="0" entrytime="00:01:32.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="140" reactiontime="+84" swimtime="00:04:02.70" resultid="17353" heatid="19092" lane="3" entrytime="00:04:00.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.95" />
                    <SPLIT distance="100" swimtime="00:01:57.61" />
                    <SPLIT distance="150" swimtime="00:03:01.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulina" lastname="Warchałowska" birthdate="2005-01-30" gender="F" nation="POL" license="103103600157" swrid="4930974" athleteid="17436">
              <RESULTS>
                <RESULT eventid="1075" points="586" reactiontime="+72" swimtime="00:01:06.28" resultid="17437" heatid="18977" lane="5" entrytime="00:01:05.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="544" reactiontime="+74" swimtime="00:02:18.39" resultid="17438" heatid="18985" lane="0" entrytime="00:02:14.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.95" />
                    <SPLIT distance="100" swimtime="00:01:06.63" />
                    <SPLIT distance="150" swimtime="00:01:42.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="493" reactiontime="+76" swimtime="00:04:59.32" resultid="17439" heatid="19007" lane="1" entrytime="00:04:40.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                    <SPLIT distance="100" swimtime="00:01:11.48" />
                    <SPLIT distance="150" swimtime="00:01:49.27" />
                    <SPLIT distance="200" swimtime="00:02:27.29" />
                    <SPLIT distance="250" swimtime="00:03:05.14" />
                    <SPLIT distance="300" swimtime="00:03:43.50" />
                    <SPLIT distance="350" swimtime="00:04:21.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="445" swimtime="00:00:31.98" resultid="17440" heatid="19017" lane="0" entrytime="00:00:31.32" entrycourse="LCM" />
                <RESULT eventid="1150" points="549" reactiontime="+75" swimtime="00:02:28.74" resultid="17441" heatid="19057" lane="4" entrytime="00:02:25.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                    <SPLIT distance="100" swimtime="00:01:10.10" />
                    <SPLIT distance="150" swimtime="00:01:49.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="508" reactiontime="+75" swimtime="00:01:04.79" resultid="17442" heatid="19065" lane="6" entrytime="00:01:03.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Szubzda" birthdate="2004-02-25" gender="F" nation="POL" license="103103600130" swrid="4792826" athleteid="17289">
              <RESULTS>
                <RESULT eventid="1059" points="540" reactiontime="+71" swimtime="00:00:29.06" resultid="17290" heatid="18950" lane="5" entrytime="00:00:28.91" entrycourse="LCM" />
                <RESULT eventid="1075" points="557" reactiontime="+73" swimtime="00:01:07.39" resultid="17291" heatid="18977" lane="6" entrytime="00:01:06.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="570" reactiontime="+73" swimtime="00:00:29.45" resultid="17292" heatid="19017" lane="3" entrytime="00:00:29.27" entrycourse="LCM" />
                <RESULT eventid="1117" points="633" reactiontime="+62" swimtime="00:00:31.41" resultid="17293" heatid="19030" lane="6" entrytime="00:00:31.53" entrycourse="LCM" />
                <RESULT eventid="1167" points="592" reactiontime="+59" swimtime="00:01:08.55" resultid="17294" heatid="19082" lane="2" entrytime="00:01:08.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00603" nation="POL" region="03" clubid="17076" name="KS ,,Wisła&apos;&apos; Puławy">
          <ATHLETES>
            <ATHLETE firstname="Klaudia" lastname="Deputat" birthdate="2008-12-31" gender="F" nation="POL" license="100603600170" swrid="5314167" athleteid="17095">
              <RESULTS>
                <RESULT eventid="1059" points="350" swimtime="00:00:33.56" resultid="17096" heatid="18946" lane="0" />
                <RESULT eventid="1091" points="339" reactiontime="+72" swimtime="00:02:56.77" resultid="17097" heatid="18993" lane="0" entrytime="00:03:10.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.33" />
                    <SPLIT distance="100" swimtime="00:01:25.10" />
                    <SPLIT distance="150" swimtime="00:02:12.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="322" reactiontime="+81" swimtime="00:05:44.81" resultid="17098" heatid="19004" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="100" swimtime="00:01:17.48" />
                    <SPLIT distance="150" swimtime="00:02:02.41" />
                    <SPLIT distance="200" swimtime="00:02:46.96" />
                    <SPLIT distance="250" swimtime="00:03:33.39" />
                    <SPLIT distance="300" swimtime="00:04:17.82" />
                    <SPLIT distance="350" swimtime="00:05:03.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="384" reactiontime="+75" swimtime="00:00:37.11" resultid="17099" heatid="19028" lane="9" entrytime="00:00:40.28" entrycourse="LCM" />
                <RESULT eventid="1167" points="366" reactiontime="+72" swimtime="00:01:20.41" resultid="17100" heatid="19078" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartłomiej" lastname="Rymkiewicz" birthdate="2009-09-11" gender="M" nation="POL" license="100603700181" swrid="5405574" athleteid="17135">
              <RESULTS>
                <RESULT eventid="1071" points="173" reactiontime="+63" swimtime="00:00:46.52" resultid="17136" heatid="18968" lane="4" />
                <RESULT eventid="1095" points="269" reactiontime="+62" swimtime="00:02:53.34" resultid="17137" heatid="18996" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.38" />
                    <SPLIT distance="100" swimtime="00:01:26.54" />
                    <SPLIT distance="150" swimtime="00:02:10.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="242" reactiontime="+63" swimtime="00:00:38.46" resultid="17138" heatid="19035" lane="2" entrytime="00:00:38.53" entrycourse="LCM" />
                <RESULT comment="K11 - Pływak wykonał nierównoczesne lub naprzemienne ruchy nóg" eventid="1145" status="DSQ" swimtime="00:03:02.36" resultid="17139" heatid="19053" lane="8" entrytime="00:03:06.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.91" />
                    <SPLIT distance="100" swimtime="00:01:26.73" />
                    <SPLIT distance="150" swimtime="00:02:22.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="244" reactiontime="+58" swimtime="00:01:22.93" resultid="17140" heatid="19086" lane="9" entrytime="00:01:25.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Pecio" birthdate="2005-01-26" gender="F" nation="POL" license="100603600089" swrid="4999904" athleteid="17115">
              <RESULTS>
                <RESULT eventid="1067" points="555" reactiontime="+67" swimtime="00:00:35.76" resultid="17116" heatid="18967" lane="3" entrytime="00:00:34.59" entrycourse="LCM" />
                <RESULT eventid="1083" points="426" reactiontime="+68" swimtime="00:02:30.15" resultid="17117" heatid="18982" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                    <SPLIT distance="100" swimtime="00:01:11.42" />
                    <SPLIT distance="150" swimtime="00:01:51.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="402" reactiontime="+53" swimtime="00:00:33.10" resultid="17118" heatid="19014" lane="2" />
                <RESULT eventid="1133" points="383" reactiontime="+69" swimtime="00:01:28.27" resultid="17119" heatid="19041" lane="9" entrytime="00:01:21.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="414" reactiontime="+68" swimtime="00:01:09.35" resultid="17120" heatid="19065" lane="2" entrytime="00:01:04.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="356" reactiontime="+68" swimtime="00:03:16.13" resultid="17121" heatid="19090" lane="4" entrytime="00:03:06.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.01" />
                    <SPLIT distance="100" swimtime="00:01:36.91" />
                    <SPLIT distance="150" swimtime="00:02:29.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Gawełko" birthdate="2006-05-27" gender="F" nation="POL" license="100603600183" swrid="5112642" athleteid="17122">
              <RESULTS>
                <RESULT eventid="1067" points="495" reactiontime="+67" swimtime="00:00:37.16" resultid="17123" heatid="18966" lane="5" entrytime="00:00:36.88" entrycourse="LCM" />
                <RESULT eventid="1083" points="514" reactiontime="+71" swimtime="00:02:21.01" resultid="17124" heatid="18984" lane="7" entrytime="00:02:20.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                    <SPLIT distance="100" swimtime="00:01:08.84" />
                    <SPLIT distance="150" swimtime="00:01:45.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="510" reactiontime="+69" swimtime="00:04:55.94" resultid="17125" heatid="19006" lane="2" entrytime="00:04:58.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                    <SPLIT distance="100" swimtime="00:01:09.08" />
                    <SPLIT distance="150" swimtime="00:01:46.74" />
                    <SPLIT distance="200" swimtime="00:02:24.61" />
                    <SPLIT distance="250" swimtime="00:03:02.99" />
                    <SPLIT distance="300" swimtime="00:03:41.23" />
                    <SPLIT distance="350" swimtime="00:04:19.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="494" reactiontime="+69" swimtime="00:01:21.12" resultid="17126" heatid="19041" lane="1" entrytime="00:01:19.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="498" reactiontime="+72" swimtime="00:01:05.21" resultid="17127" heatid="19065" lane="1" entrytime="00:01:05.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="485" reactiontime="+71" swimtime="00:02:56.95" resultid="17128" heatid="19091" lane="2" entrytime="00:02:53.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.74" />
                    <SPLIT distance="100" swimtime="00:01:25.10" />
                    <SPLIT distance="150" swimtime="00:02:11.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hubert" lastname="Żaczek" birthdate="2008-01-02" gender="M" nation="POL" license="100603700158" swrid="5243444" athleteid="17148">
              <RESULTS>
                <RESULT eventid="1079" points="333" reactiontime="+71" swimtime="00:01:11.35" resultid="17149" heatid="18978" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="M10 - Pływak nie dotknął ściany dwiema dłońmi przy nawrocie lub na zakończenie wyścigu" eventid="1103" reactiontime="+70" status="DSQ" swimtime="00:05:27.94" resultid="17150" heatid="19001" lane="2" entrytime="00:05:34.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                    <SPLIT distance="100" swimtime="00:01:14.70" />
                    <SPLIT distance="150" swimtime="00:01:56.94" />
                    <SPLIT distance="200" swimtime="00:02:37.83" />
                    <SPLIT distance="250" swimtime="00:03:25.64" />
                    <SPLIT distance="300" swimtime="00:04:13.34" />
                    <SPLIT distance="350" swimtime="00:04:51.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="391" reactiontime="+63" swimtime="00:00:32.80" resultid="17151" heatid="19036" lane="1" entrytime="00:00:33.75" entrycourse="LCM" />
                <RESULT eventid="1145" points="415" reactiontime="+55" swimtime="00:02:32.72" resultid="17152" heatid="19053" lane="5" entrytime="00:02:38.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                    <SPLIT distance="100" swimtime="00:01:12.45" />
                    <SPLIT distance="150" swimtime="00:01:58.68" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej, a przed sygnałem startu" eventid="1171" reactiontime="+42" status="DSQ" swimtime="00:01:12.06" resultid="17153" heatid="19087" lane="7" entrytime="00:01:12.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nikola" lastname="Jasik" birthdate="2006-07-17" gender="F" nation="POL" license="100603600131" swrid="4416128" athleteid="17082">
              <RESULTS>
                <RESULT eventid="1059" points="534" reactiontime="+70" swimtime="00:00:29.16" resultid="17083" heatid="18950" lane="4" entrytime="00:00:28.50" entrycourse="LCM" />
                <RESULT eventid="1075" points="487" reactiontime="+73" swimtime="00:01:10.47" resultid="17084" heatid="18977" lane="7" entrytime="00:01:07.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="525" reactiontime="+72" swimtime="00:00:30.27" resultid="17085" heatid="19017" lane="7" entrytime="00:00:29.83" entrycourse="LCM" />
                <RESULT eventid="1133" points="460" reactiontime="+73" swimtime="00:01:23.03" resultid="17086" heatid="19040" lane="4" entrytime="00:01:22.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="511" reactiontime="+72" swimtime="00:01:04.64" resultid="17087" heatid="19065" lane="3" entrytime="00:01:03.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" status="DNS" swimtime="00:00:00.00" resultid="17088" heatid="19089" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Król" birthdate="2006-02-27" gender="F" nation="POL" license="100603600123" swrid="4909923" athleteid="17108">
              <RESULTS>
                <RESULT eventid="1067" points="600" reactiontime="+64" swimtime="00:00:34.84" resultid="17109" heatid="18967" lane="6" entrytime="00:00:35.33" entrycourse="LCM" />
                <RESULT eventid="1099" points="684" reactiontime="+67" swimtime="00:05:02.20" resultid="17110" heatid="18999" lane="5" entrytime="00:05:08.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.85" />
                    <SPLIT distance="100" swimtime="00:01:08.90" />
                    <SPLIT distance="150" swimtime="00:01:49.16" />
                    <SPLIT distance="200" swimtime="00:02:27.40" />
                    <SPLIT distance="250" swimtime="00:03:10.63" />
                    <SPLIT distance="300" swimtime="00:03:53.82" />
                    <SPLIT distance="350" swimtime="00:04:28.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="702" reactiontime="+59" swimtime="00:00:30.35" resultid="17111" heatid="19030" lane="4" entrytime="00:00:29.97" entrycourse="LCM" />
                <RESULT eventid="1141" points="666" reactiontime="+72" swimtime="00:02:24.41" resultid="17112" heatid="19050" lane="4" entrytime="00:02:23.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                    <SPLIT distance="100" swimtime="00:01:08.80" />
                    <SPLIT distance="150" swimtime="00:01:52.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="657" reactiontime="+71" swimtime="00:00:59.47" resultid="17113" heatid="19066" lane="3" entrytime="00:00:58.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="564" reactiontime="+72" swimtime="00:02:48.31" resultid="17114" heatid="19091" lane="3" entrytime="00:02:48.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                    <SPLIT distance="100" swimtime="00:01:21.68" />
                    <SPLIT distance="150" swimtime="00:02:05.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Damian" lastname="Baraban" birthdate="2008-05-07" gender="M" nation="POL" license="100603700171" swrid="5314175" athleteid="17101">
              <RESULTS>
                <RESULT eventid="1063" points="231" reactiontime="+78" swimtime="00:00:34.07" resultid="17102" heatid="18957" lane="7" entrytime="00:00:33.68" entrycourse="LCM" />
                <RESULT eventid="1079" points="149" swimtime="00:01:33.32" resultid="17103" heatid="18979" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="250" reactiontime="+53" swimtime="00:05:49.16" resultid="17104" heatid="19010" lane="8" entrytime="00:05:45.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.10" />
                    <SPLIT distance="100" swimtime="00:01:21.78" />
                    <SPLIT distance="150" swimtime="00:02:06.53" />
                    <SPLIT distance="200" swimtime="00:02:50.79" />
                    <SPLIT distance="250" swimtime="00:03:36.29" />
                    <SPLIT distance="300" swimtime="00:04:20.97" />
                    <SPLIT distance="350" swimtime="00:05:06.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1137" points="162" reactiontime="+82" swimtime="00:01:44.22" resultid="17105" heatid="19044" lane="3" entrytime="00:01:41.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="184" reactiontime="+68" swimtime="00:03:14.62" resultid="17106" heatid="19058" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.61" />
                    <SPLIT distance="100" swimtime="00:01:32.89" />
                    <SPLIT distance="150" swimtime="00:02:26.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="232" reactiontime="+60" swimtime="00:01:16.32" resultid="17107" heatid="19070" lane="8" entrytime="00:01:18.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwia" lastname="Wit" birthdate="2008-03-08" gender="F" nation="POL" license="100603600194" swrid="5322634" athleteid="17089">
              <RESULTS>
                <RESULT eventid="1059" points="439" reactiontime="+52" swimtime="00:00:31.13" resultid="17090" heatid="18949" lane="9" entrytime="00:00:31.72" entrycourse="LCM" />
                <RESULT eventid="1083" points="386" reactiontime="+68" swimtime="00:02:35.06" resultid="17091" heatid="18983" lane="8" entrytime="00:02:34.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                    <SPLIT distance="100" swimtime="00:01:14.53" />
                    <SPLIT distance="150" swimtime="00:01:55.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="357" reactiontime="+73" swimtime="00:05:33.32" resultid="17092" heatid="19005" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.91" />
                    <SPLIT distance="100" swimtime="00:01:17.02" />
                    <SPLIT distance="150" swimtime="00:01:59.73" />
                    <SPLIT distance="200" swimtime="00:02:42.73" />
                    <SPLIT distance="250" swimtime="00:03:25.06" />
                    <SPLIT distance="300" swimtime="00:04:09.29" />
                    <SPLIT distance="350" swimtime="00:04:50.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="248" reactiontime="+70" swimtime="00:00:38.84" resultid="17093" heatid="19015" lane="7" entrytime="00:00:37.96" entrycourse="LCM" />
                <RESULT eventid="1159" points="381" reactiontime="+71" swimtime="00:01:11.30" resultid="17094" heatid="19063" lane="7" entrytime="00:01:10.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Bocianowska" birthdate="2008-09-01" gender="F" nation="POL" license="100603600151" swrid="5233350" athleteid="17141">
              <RESULTS>
                <RESULT eventid="1075" points="346" reactiontime="+94" swimtime="00:01:18.98" resultid="17142" heatid="18975" lane="4" entrytime="00:01:21.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="359" reactiontime="+87" swimtime="00:06:14.73" resultid="17143" heatid="18998" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                    <SPLIT distance="100" swimtime="00:01:20.82" />
                    <SPLIT distance="150" swimtime="00:02:12.71" />
                    <SPLIT distance="200" swimtime="00:03:00.36" />
                    <SPLIT distance="250" swimtime="00:03:55.04" />
                    <SPLIT distance="300" swimtime="00:04:49.62" />
                    <SPLIT distance="350" swimtime="00:05:32.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="382" reactiontime="+92" swimtime="00:00:33.66" resultid="17144" heatid="19015" lane="6" entrytime="00:00:36.26" entrycourse="LCM" />
                <RESULT eventid="1141" points="352" reactiontime="+93" swimtime="00:02:58.53" resultid="17145" heatid="19048" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.25" />
                    <SPLIT distance="100" swimtime="00:01:23.40" />
                    <SPLIT distance="150" swimtime="00:02:16.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="323" reactiontime="+91" swimtime="00:01:15.29" resultid="17146" heatid="19063" lane="9" entrytime="00:01:14.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="270" reactiontime="+80" swimtime="00:01:29.04" resultid="17147" heatid="19080" lane="0" entrytime="00:01:28.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Sala" birthdate="2008-01-06" gender="M" nation="POL" license="100603700156" swrid="5243443" athleteid="17129">
              <RESULTS>
                <RESULT eventid="1071" points="369" reactiontime="+70" swimtime="00:00:36.16" resultid="17130" heatid="18973" lane="7" entrytime="00:00:37.48" entrycourse="LCM" />
                <RESULT eventid="1103" points="296" reactiontime="+73" swimtime="00:06:05.82" resultid="17131" heatid="19000" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.74" />
                    <SPLIT distance="100" swimtime="00:01:25.82" />
                    <SPLIT distance="150" swimtime="00:02:16.43" />
                    <SPLIT distance="200" swimtime="00:03:02.41" />
                    <SPLIT distance="250" swimtime="00:03:50.74" />
                    <SPLIT distance="300" swimtime="00:04:39.66" />
                    <SPLIT distance="350" swimtime="00:05:22.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="330" reactiontime="+68" swimtime="00:00:32.21" resultid="17132" heatid="19022" lane="3" entrytime="00:00:32.45" entrycourse="LCM" />
                <RESULT eventid="1137" points="343" reactiontime="+70" swimtime="00:01:21.23" resultid="17133" heatid="19046" lane="1" entrytime="00:01:25.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="341" reactiontime="+68" swimtime="00:03:00.49" resultid="17134" heatid="19093" lane="4" entrytime="00:03:10.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.37" />
                    <SPLIT distance="100" swimtime="00:01:27.60" />
                    <SPLIT distance="150" swimtime="00:02:16.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Słotwińska" birthdate="2005-11-29" gender="F" nation="POL" license="100603600094" swrid="4909922" athleteid="17077">
              <RESULTS>
                <RESULT eventid="1059" points="421" reactiontime="+90" swimtime="00:00:31.56" resultid="17078" heatid="18949" lane="3" entrytime="00:00:30.68" entrycourse="LCM" />
                <RESULT eventid="1083" points="437" reactiontime="+93" swimtime="00:02:28.88" resultid="17079" heatid="18983" lane="4" entrytime="00:02:27.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.54" />
                    <SPLIT distance="100" swimtime="00:01:14.14" />
                    <SPLIT distance="150" swimtime="00:01:53.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="323" reactiontime="+85" swimtime="00:00:35.59" resultid="17080" heatid="19014" lane="3" />
                <RESULT eventid="1159" points="374" reactiontime="+92" swimtime="00:01:11.71" resultid="17081" heatid="19063" lane="4" entrytime="00:01:08.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01203" nation="POL" region="03" clubid="18339" name="UKS ,,Trójka&apos;&apos; Puławy">
          <ATHLETES>
            <ATHLETE firstname="Sebastian" lastname="Gogacz" birthdate="1976-10-28" gender="M" nation="POL" license="501203700057" swrid="4754646" athleteid="18359">
              <RESULTS>
                <RESULT eventid="1079" points="381" reactiontime="+80" swimtime="00:01:08.24" resultid="18360" heatid="18979" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="354" reactiontime="+84" swimtime="00:05:11.03" resultid="18361" heatid="19008" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                    <SPLIT distance="100" swimtime="00:01:15.36" />
                    <SPLIT distance="150" swimtime="00:01:55.10" />
                    <SPLIT distance="200" swimtime="00:02:34.30" />
                    <SPLIT distance="250" swimtime="00:03:13.15" />
                    <SPLIT distance="300" swimtime="00:03:52.76" />
                    <SPLIT distance="350" swimtime="00:04:32.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="323" reactiontime="+84" swimtime="00:02:46.14" resultid="18362" heatid="19052" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                    <SPLIT distance="100" swimtime="00:01:20.77" />
                    <SPLIT distance="150" swimtime="00:02:07.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Przybylska" birthdate="2009-09-03" gender="F" nation="POL" license="101203600063" swrid="5322645" athleteid="18340">
              <RESULTS>
                <RESULT eventid="1059" points="237" swimtime="00:00:38.24" resultid="18341" heatid="18948" lane="9" entrytime="00:00:36.19" entrycourse="LCM" />
                <RESULT eventid="1091" points="205" reactiontime="+70" swimtime="00:03:28.91" resultid="18342" heatid="18992" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.08" />
                    <SPLIT distance="100" swimtime="00:01:44.23" />
                    <SPLIT distance="150" swimtime="00:02:38.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="178" swimtime="00:00:43.39" resultid="18343" heatid="19015" lane="0" entrytime="00:00:42.19" entrycourse="LCM" />
                <RESULT eventid="1117" points="215" reactiontime="+71" swimtime="00:00:44.97" resultid="18344" heatid="19027" lane="6" entrytime="00:00:43.72" entrycourse="LCM" />
                <RESULT eventid="1159" points="251" swimtime="00:01:21.94" resultid="18345" heatid="19062" lane="2" entrytime="00:01:20.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="203" reactiontime="+72" swimtime="00:01:37.81" resultid="18346" heatid="19079" lane="3" entrytime="00:01:37.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tymoteusz" lastname="Bielawski" birthdate="2006-10-16" gender="M" nation="POL" license="101203700049" swrid="5009216" athleteid="18352">
              <RESULTS>
                <RESULT eventid="1063" points="389" reactiontime="+75" swimtime="00:00:28.62" resultid="18353" heatid="18960" lane="1" entrytime="00:00:28.75" entrycourse="LCM" />
                <RESULT eventid="1071" points="302" reactiontime="+77" swimtime="00:00:38.67" resultid="18354" heatid="18972" lane="4" entrytime="00:00:38.27" entrycourse="LCM" />
                <RESULT eventid="1113" points="355" reactiontime="+74" swimtime="00:00:31.44" resultid="18355" heatid="19023" lane="8" entrytime="00:00:31.13" entrycourse="LCM" />
                <RESULT eventid="1121" points="311" reactiontime="+73" swimtime="00:00:35.40" resultid="18356" heatid="19033" lane="8" />
                <RESULT eventid="1163" status="DNS" swimtime="00:00:00.00" resultid="18357" heatid="19074" lane="9" entrytime="00:01:03.64" entrycourse="LCM" />
                <RESULT eventid="1171" status="DNS" swimtime="00:00:00.00" resultid="18358" heatid="19084" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karina" lastname="Surowiecka" birthdate="2008-08-02" gender="F" nation="POL" license="101203600098" swrid="5461064" athleteid="18347">
              <RESULTS>
                <RESULT eventid="1059" points="291" reactiontime="+73" swimtime="00:00:35.71" resultid="18348" heatid="18948" lane="8" entrytime="00:00:35.63" entrycourse="LCM" />
                <RESULT eventid="1067" points="206" reactiontime="+88" swimtime="00:00:49.74" resultid="18349" heatid="18965" lane="6" entrytime="00:00:47.42" entrycourse="LCM" />
                <RESULT eventid="1117" points="263" reactiontime="+80" swimtime="00:00:42.08" resultid="18350" heatid="19027" lane="4" entrytime="00:00:41.47" entrycourse="LCM" />
                <RESULT eventid="1159" points="249" reactiontime="+88" swimtime="00:01:22.19" resultid="18351" heatid="19061" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04003" nation="POL" region="03" clubid="17974" name="UKP Bychawa">
          <ATHLETES>
            <ATHLETE firstname="Alan" lastname="Janik" birthdate="2008-02-19" gender="M" nation="POL" license="104003700016" swrid="5140940" athleteid="18029">
              <RESULTS>
                <RESULT eventid="1079" points="230" reactiontime="+69" swimtime="00:01:20.74" resultid="18030" heatid="18979" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1087" points="246" reactiontime="+56" swimtime="00:02:42.63" resultid="18031" heatid="18987" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="271" reactiontime="+66" swimtime="00:00:34.40" resultid="18032" heatid="19019" lane="6" />
                <RESULT eventid="1145" points="244" reactiontime="+67" swimtime="00:03:02.42" resultid="18033" heatid="19052" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.78" />
                    <SPLIT distance="100" swimtime="00:01:24.32" />
                    <SPLIT distance="150" swimtime="00:02:21.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="271" reactiontime="+68" swimtime="00:01:12.41" resultid="18034" heatid="19067" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amelia" lastname="Prącik" birthdate="2008-04-06" gender="F" nation="POL" license="104003600012" swrid="5335564" athleteid="18022">
              <RESULTS>
                <RESULT eventid="1075" points="256" reactiontime="+75" swimtime="00:01:27.34" resultid="18023" heatid="18975" lane="6" entrytime="00:01:30.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="320" reactiontime="+76" swimtime="00:06:29.06" resultid="18024" heatid="18999" lane="0" entrytime="00:06:35.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.28" />
                    <SPLIT distance="100" swimtime="00:01:28.37" />
                    <SPLIT distance="150" swimtime="00:02:15.66" />
                    <SPLIT distance="200" swimtime="00:03:02.08" />
                    <SPLIT distance="250" swimtime="00:04:01.50" />
                    <SPLIT distance="300" swimtime="00:05:00.43" />
                    <SPLIT distance="350" swimtime="00:05:45.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="300" reactiontime="+78" swimtime="00:05:52.97" resultid="18025" heatid="19005" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.83" />
                    <SPLIT distance="100" swimtime="00:01:20.69" />
                    <SPLIT distance="150" swimtime="00:02:05.26" />
                    <SPLIT distance="200" swimtime="00:02:51.25" />
                    <SPLIT distance="250" swimtime="00:03:36.73" />
                    <SPLIT distance="300" swimtime="00:04:23.88" />
                    <SPLIT distance="350" swimtime="00:05:09.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="314" reactiontime="+60" swimtime="00:03:05.38" resultid="18026" heatid="19049" lane="8" entrytime="00:03:08.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                    <SPLIT distance="100" swimtime="00:01:23.87" />
                    <SPLIT distance="150" swimtime="00:02:22.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1150" points="196" reactiontime="+76" swimtime="00:03:29.46" resultid="18027" heatid="19056" lane="4" entrytime="00:03:18.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.28" />
                    <SPLIT distance="100" swimtime="00:01:39.27" />
                    <SPLIT distance="150" swimtime="00:02:34.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="325" reactiontime="+73" swimtime="00:01:23.66" resultid="18028" heatid="19078" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcel" lastname="Nowak" birthdate="2008-04-18" gender="M" nation="POL" license="104003700020" swrid="5427439" athleteid="17997">
              <RESULTS>
                <RESULT eventid="1063" points="227" reactiontime="+77" swimtime="00:00:34.27" resultid="17998" heatid="18955" lane="7" entrytime="00:00:39.67" entrycourse="LCM" />
                <RESULT eventid="1071" points="150" reactiontime="+79" swimtime="00:00:48.79" resultid="17999" heatid="18970" lane="7" entrytime="00:00:50.04" entrycourse="LCM" />
                <RESULT eventid="1121" points="151" reactiontime="+84" swimtime="00:00:45.01" resultid="18000" heatid="19033" lane="9" />
                <RESULT eventid="1137" points="137" reactiontime="+75" swimtime="00:01:50.14" resultid="18001" heatid="19044" lane="1" entrytime="00:01:50.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="188" reactiontime="+74" swimtime="00:01:21.81" resultid="18002" heatid="19070" lane="9" entrytime="00:01:21.63" entrycourse="LCM" />
                <RESULT eventid="1171" points="135" reactiontime="+79" swimtime="00:01:40.90" resultid="18003" heatid="19083" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Szafran" birthdate="2007-01-13" gender="M" nation="POL" license="104003700017" swrid="5141046" athleteid="18015">
              <RESULTS>
                <RESULT eventid="1063" points="321" reactiontime="+86" swimtime="00:00:30.53" resultid="18016" heatid="18954" lane="8" />
                <RESULT eventid="1087" points="234" reactiontime="+92" swimtime="00:02:45.34" resultid="18017" heatid="18989" lane="0" entrytime="00:02:42.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.30" />
                    <SPLIT distance="100" swimtime="00:01:16.45" />
                    <SPLIT distance="150" swimtime="00:02:00.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="281" reactiontime="+76" swimtime="00:00:33.99" resultid="18018" heatid="19022" lane="8" entrytime="00:00:36.37" entrycourse="LCM" />
                <RESULT eventid="1121" points="268" reactiontime="+90" swimtime="00:00:37.22" resultid="18019" heatid="19035" lane="3" entrytime="00:00:38.08" entrycourse="LCM" />
                <RESULT eventid="1163" points="286" reactiontime="+96" swimtime="00:01:11.12" resultid="18020" heatid="19071" lane="9" entrytime="00:01:16.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="262" reactiontime="+83" swimtime="00:01:21.03" resultid="18021" heatid="19086" lane="8" entrytime="00:01:21.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ernest" lastname="Biernat" birthdate="2009-07-13" gender="M" nation="POL" license="104003700022" swrid="5431064" athleteid="17987">
              <RESULTS>
                <RESULT eventid="1063" status="DNS" swimtime="00:00:00.00" resultid="17988" heatid="18954" lane="6" entrytime="00:00:43.75" entrycourse="LCM" />
                <RESULT eventid="1071" status="DNS" swimtime="00:00:00.00" resultid="17989" heatid="18968" lane="5" />
                <RESULT eventid="1137" status="DNS" swimtime="00:00:00.00" resultid="17990" heatid="19044" lane="9" entrytime="00:02:16.11" entrycourse="LCM" />
                <RESULT eventid="1163" status="DNS" swimtime="00:00:00.00" resultid="17991" heatid="19068" lane="2" entrytime="00:01:43.70" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Erwin" lastname="Rechul" birthdate="2008-07-14" gender="M" nation="POL" license="104003700023" swrid="5431089" athleteid="17992">
              <RESULTS>
                <RESULT eventid="1063" points="83" reactiontime="+92" swimtime="00:00:47.76" resultid="17993" heatid="18953" lane="4" />
                <RESULT eventid="1071" points="80" reactiontime="+87" swimtime="00:01:00.18" resultid="17994" heatid="18969" lane="6" />
                <RESULT eventid="1121" points="102" reactiontime="+73" swimtime="00:00:51.26" resultid="17995" heatid="19032" lane="7" />
                <RESULT eventid="1163" points="89" reactiontime="+87" swimtime="00:01:44.73" resultid="17996" heatid="19067" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alicja" lastname="Nowicka" birthdate="2006-07-29" gender="F" nation="POL" license="104003600003" swrid="5288433" athleteid="17978">
              <RESULTS>
                <RESULT eventid="1059" points="126" reactiontime="+95" swimtime="00:00:47.16" resultid="17979" heatid="18946" lane="3" entrytime="00:00:44.57" entrycourse="LCM" />
                <RESULT eventid="1067" points="170" reactiontime="+90" swimtime="00:00:52.99" resultid="17980" heatid="18964" lane="6" entrytime="00:00:54.98" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Góźdź" birthdate="2006-07-07" gender="M" nation="POL" license="104003700001" swrid="5340916" athleteid="18004">
              <RESULTS>
                <RESULT eventid="1063" points="298" reactiontime="+84" swimtime="00:00:31.30" resultid="18005" heatid="18957" lane="5" entrytime="00:00:33.18" entrycourse="LCM" />
                <RESULT eventid="1071" points="262" reactiontime="+90" swimtime="00:00:40.55" resultid="18006" heatid="18972" lane="8" entrytime="00:00:41.48" entrycourse="LCM" />
                <RESULT eventid="1113" points="233" reactiontime="+85" swimtime="00:00:36.18" resultid="18007" heatid="19019" lane="5" />
                <RESULT eventid="1137" points="233" reactiontime="+84" swimtime="00:01:32.41" resultid="18008" heatid="19045" lane="2" entrytime="00:01:34.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="293" reactiontime="+84" swimtime="00:01:10.55" resultid="18009" heatid="19071" lane="2" entrytime="00:01:14.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Batko" birthdate="2007-07-02" gender="M" nation="POL" license="104003700015" swrid="5353686" athleteid="17981">
              <RESULTS>
                <RESULT eventid="1063" points="283" reactiontime="+79" swimtime="00:00:31.83" resultid="17982" heatid="18958" lane="6" entrytime="00:00:31.88" entrycourse="LCM" />
                <RESULT eventid="1071" status="DNS" swimtime="00:00:00.00" resultid="17983" heatid="18971" lane="1" entrytime="00:00:44.61" entrycourse="LCM" />
                <RESULT eventid="1113" points="175" reactiontime="+86" swimtime="00:00:39.77" resultid="17984" heatid="19021" lane="1" entrytime="00:00:42.60" entrycourse="LCM" />
                <RESULT comment="K4 - Pływak wykonał cykl ruchowy inny niż jeden ruch ramion i jedno kopnięcie nogami (z wyjątkiem ostatniego cyklu przed nawrotem lub zakończeniem wyścigu)" eventid="1137" reactiontime="+85" status="DSQ" swimtime="00:01:38.64" resultid="17985" heatid="19044" lane="6" entrytime="00:01:42.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="189" reactiontime="+86" swimtime="00:01:21.66" resultid="17986" heatid="19071" lane="0" entrytime="00:01:16.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Lipiński" birthdate="2007-10-03" gender="M" nation="POL" license="104003700004" swrid="5335562" athleteid="18042">
              <RESULTS>
                <RESULT eventid="1087" points="402" reactiontime="+71" swimtime="00:02:18.19" resultid="18043" heatid="18990" lane="1" entrytime="00:02:20.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                    <SPLIT distance="100" swimtime="00:01:05.88" />
                    <SPLIT distance="150" swimtime="00:01:41.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="336" reactiontime="+76" swimtime="00:05:50.55" resultid="18044" heatid="19001" lane="8" entrytime="00:05:56.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                    <SPLIT distance="100" swimtime="00:01:10.28" />
                    <SPLIT distance="150" swimtime="00:01:55.93" />
                    <SPLIT distance="200" swimtime="00:02:40.31" />
                    <SPLIT distance="250" swimtime="00:03:33.40" />
                    <SPLIT distance="300" swimtime="00:04:27.55" />
                    <SPLIT distance="350" swimtime="00:05:08.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="395" reactiontime="+72" swimtime="00:04:59.75" resultid="18045" heatid="19010" lane="7" entrytime="00:05:03.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                    <SPLIT distance="100" swimtime="00:01:09.33" />
                    <SPLIT distance="150" swimtime="00:01:46.68" />
                    <SPLIT distance="200" swimtime="00:02:25.10" />
                    <SPLIT distance="250" swimtime="00:03:03.61" />
                    <SPLIT distance="300" swimtime="00:03:42.94" />
                    <SPLIT distance="350" swimtime="00:04:23.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="349" reactiontime="+74" swimtime="00:00:31.63" resultid="18046" heatid="19018" lane="5" />
                <RESULT eventid="1163" points="413" reactiontime="+72" swimtime="00:01:02.96" resultid="18047" heatid="19074" lane="8" entrytime="00:01:02.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="341" reactiontime="+72" swimtime="00:20:45.61" resultid="18048" heatid="19099" lane="3" entrytime="00:20:32.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                    <SPLIT distance="100" swimtime="00:01:12.18" />
                    <SPLIT distance="150" swimtime="00:01:52.31" />
                    <SPLIT distance="200" swimtime="00:02:33.33" />
                    <SPLIT distance="250" swimtime="00:03:14.73" />
                    <SPLIT distance="300" swimtime="00:03:56.48" />
                    <SPLIT distance="350" swimtime="00:04:37.57" />
                    <SPLIT distance="400" swimtime="00:05:19.81" />
                    <SPLIT distance="450" swimtime="00:06:02.17" />
                    <SPLIT distance="500" swimtime="00:06:44.40" />
                    <SPLIT distance="550" swimtime="00:07:26.18" />
                    <SPLIT distance="600" swimtime="00:08:08.22" />
                    <SPLIT distance="650" swimtime="00:08:49.37" />
                    <SPLIT distance="700" swimtime="00:09:32.72" />
                    <SPLIT distance="750" swimtime="00:10:14.88" />
                    <SPLIT distance="800" swimtime="00:10:57.39" />
                    <SPLIT distance="850" swimtime="00:11:41.08" />
                    <SPLIT distance="900" swimtime="00:12:21.07" />
                    <SPLIT distance="950" swimtime="00:13:04.66" />
                    <SPLIT distance="1000" swimtime="00:13:46.07" />
                    <SPLIT distance="1050" swimtime="00:14:29.48" />
                    <SPLIT distance="1100" swimtime="00:15:10.04" />
                    <SPLIT distance="1150" swimtime="00:15:53.22" />
                    <SPLIT distance="1200" swimtime="00:16:36.19" />
                    <SPLIT distance="1250" swimtime="00:17:17.98" />
                    <SPLIT distance="1300" swimtime="00:18:00.68" />
                    <SPLIT distance="1350" swimtime="00:18:42.90" />
                    <SPLIT distance="1400" swimtime="00:19:25.15" />
                    <SPLIT distance="1450" swimtime="00:20:06.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łucja" lastname="Frączek" birthdate="2008-02-29" gender="F" nation="POL" license="104003600005" swrid="5335563" athleteid="18035">
              <RESULTS>
                <RESULT eventid="1083" points="396" reactiontime="+94" swimtime="00:02:33.78" resultid="18036" heatid="18983" lane="0" entrytime="00:02:34.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                    <SPLIT distance="100" swimtime="00:01:16.52" />
                    <SPLIT distance="150" swimtime="00:01:58.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1091" points="432" swimtime="00:02:43.17" resultid="18037" heatid="18993" lane="6" entrytime="00:02:44.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.09" />
                    <SPLIT distance="100" swimtime="00:01:19.77" />
                    <SPLIT distance="150" swimtime="00:02:02.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="376" reactiontime="+93" swimtime="00:05:27.40" resultid="18038" heatid="19005" lane="6" entrytime="00:05:31.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.58" />
                    <SPLIT distance="100" swimtime="00:01:17.63" />
                    <SPLIT distance="150" swimtime="00:01:59.94" />
                    <SPLIT distance="200" swimtime="00:02:42.35" />
                    <SPLIT distance="250" swimtime="00:03:24.74" />
                    <SPLIT distance="300" swimtime="00:04:08.13" />
                    <SPLIT distance="350" swimtime="00:04:50.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="485" reactiontime="+82" swimtime="00:00:34.33" resultid="18039" heatid="19029" lane="0" entrytime="00:00:35.57" entrycourse="LCM" />
                <RESULT eventid="1167" points="424" reactiontime="+89" swimtime="00:01:16.60" resultid="18040" heatid="19081" lane="0" entrytime="00:01:17.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="369" swimtime="00:11:15.46" resultid="18041" heatid="19096" lane="7" entrytime="00:11:28.24" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Teter" birthdate="2009-05-02" gender="M" nation="POL" license="104003700024" swrid="5431096" athleteid="18010">
              <RESULTS>
                <RESULT eventid="1063" points="117" reactiontime="+73" swimtime="00:00:42.75" resultid="18011" heatid="18953" lane="8" />
                <RESULT eventid="1071" points="105" swimtime="00:00:54.88" resultid="18012" heatid="18969" lane="1" />
                <RESULT eventid="1121" points="113" reactiontime="+78" swimtime="00:00:49.62" resultid="18013" heatid="19032" lane="8" />
                <RESULT eventid="1163" points="97" swimtime="00:01:41.93" resultid="18014" heatid="19068" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrianna" lastname="Nowicka" birthdate="2009-10-02" gender="F" nation="POL" license="104003600002" swrid="5340918" athleteid="17975">
              <RESULTS>
                <RESULT eventid="1059" points="177" reactiontime="+92" swimtime="00:00:42.11" resultid="17976" heatid="18945" lane="6" />
                <RESULT eventid="1067" points="102" swimtime="00:01:02.83" resultid="17977" heatid="18964" lane="7" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04214" nation="POL" region="14" clubid="18575" name="Warsaw Masters Team">
          <ATHLETES>
            <ATHLETE firstname="Anna" lastname="Szemberg" birthdate="1949-07-26" gender="F" nation="POL" license="504214600017" swrid="4302692" athleteid="18576">
              <RESULTS>
                <RESULT eventid="1059" points="64" status="EXH" swimtime="00:00:59.07" resultid="18577" heatid="18945" lane="3" />
                <RESULT eventid="1083" points="66" status="EXH" swimtime="00:04:39.07" resultid="18578" heatid="18982" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.31" />
                    <SPLIT distance="100" swimtime="00:02:16.01" />
                    <SPLIT distance="150" swimtime="00:03:29.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="68" status="EXH" swimtime="00:09:38.19" resultid="18579" heatid="19004" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.61" />
                    <SPLIT distance="100" swimtime="00:02:17.30" />
                    <SPLIT distance="150" swimtime="00:03:31.78" />
                    <SPLIT distance="200" swimtime="00:04:44.84" />
                    <SPLIT distance="250" swimtime="00:05:59.24" />
                    <SPLIT distance="300" swimtime="00:07:12.53" />
                    <SPLIT distance="350" swimtime="00:08:26.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="58" status="EXH" swimtime="00:02:13.01" resultid="18580" heatid="19061" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02003" nation="POL" region="03" clubid="18389" name="Uks 51">
          <ATHLETES>
            <ATHLETE firstname="Filip" lastname="Suchański" birthdate="2005-10-06" gender="M" nation="POL" license="102003700025" swrid="4931007" athleteid="18434">
              <RESULTS>
                <RESULT eventid="1095" points="632" reactiontime="+63" swimtime="00:02:10.39" resultid="18435" heatid="18997" lane="4" entrytime="00:02:10.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                    <SPLIT distance="100" swimtime="00:01:03.11" />
                    <SPLIT distance="150" swimtime="00:01:37.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="590" reactiontime="+68" swimtime="00:04:22.36" resultid="18436" heatid="19012" lane="9" entrytime="00:04:26.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.82" />
                    <SPLIT distance="100" swimtime="00:01:00.78" />
                    <SPLIT distance="150" swimtime="00:01:34.23" />
                    <SPLIT distance="200" swimtime="00:02:08.07" />
                    <SPLIT distance="250" swimtime="00:02:41.91" />
                    <SPLIT distance="300" swimtime="00:03:15.47" />
                    <SPLIT distance="350" swimtime="00:03:49.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="495" reactiontime="+70" swimtime="00:02:19.94" resultid="18437" heatid="19059" lane="7" entrytime="00:02:19.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.24" />
                    <SPLIT distance="100" swimtime="00:01:04.12" />
                    <SPLIT distance="150" swimtime="00:01:42.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="605" reactiontime="+66" swimtime="00:01:01.29" resultid="18438" heatid="19088" lane="3" entrytime="00:01:01.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Hapak" birthdate="2009-04-28" gender="F" nation="POL" license="102003600097" swrid="5193103" athleteid="18399">
              <RESULTS>
                <RESULT eventid="1059" points="423" reactiontime="+75" swimtime="00:00:31.51" resultid="18400" heatid="18948" lane="5" entrytime="00:00:32.40" entrycourse="LCM" />
                <RESULT eventid="1117" points="366" reactiontime="+87" swimtime="00:00:37.70" resultid="18401" heatid="19028" lane="7" entrytime="00:00:38.72" entrycourse="LCM" />
                <RESULT eventid="1159" points="380" reactiontime="+86" swimtime="00:01:11.33" resultid="18402" heatid="19063" lane="1" entrytime="00:01:10.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="312" reactiontime="+91" swimtime="00:01:24.83" resultid="18403" heatid="19080" lane="2" entrytime="00:01:23.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Niezgoda" birthdate="2007-01-04" gender="F" nation="POL" license="102003600078" swrid="5148657" athleteid="18390">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="18391" heatid="18950" lane="1" entrytime="00:00:30.09" entrycourse="LCM" />
                <RESULT eventid="1117" status="DNS" swimtime="00:00:00.00" resultid="18392" heatid="19029" lane="9" entrytime="00:00:35.59" entrycourse="LCM" />
                <RESULT eventid="1159" status="DNS" swimtime="00:00:00.00" resultid="18393" heatid="19064" lane="6" entrytime="00:01:07.08" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robert" lastname="Wajler" birthdate="2007-09-18" gender="M" nation="POL" license="102003700074" swrid="5148659" athleteid="18414">
              <RESULTS>
                <RESULT eventid="1063" points="208" reactiontime="+83" swimtime="00:00:35.25" resultid="18415" heatid="18954" lane="7" />
                <RESULT eventid="1079" points="164" swimtime="00:01:30.43" resultid="18416" heatid="18979" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="160" swimtime="00:00:40.94" resultid="18417" heatid="19019" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Ciurska" birthdate="2006-10-20" gender="F" nation="POL" license="102003600030" swrid="5006503" athleteid="18428">
              <RESULTS>
                <RESULT eventid="1091" points="532" reactiontime="+73" swimtime="00:02:32.22" resultid="18429" heatid="18994" lane="8" entrytime="00:02:32.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.62" />
                    <SPLIT distance="100" swimtime="00:01:13.86" />
                    <SPLIT distance="150" swimtime="00:01:53.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="505" reactiontime="+76" swimtime="00:00:33.88" resultid="18430" heatid="19029" lane="2" entrytime="00:00:34.25" entrycourse="LCM" />
                <RESULT eventid="1141" points="455" reactiontime="+89" swimtime="00:02:43.97" resultid="18431" heatid="19049" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                    <SPLIT distance="100" swimtime="00:01:16.64" />
                    <SPLIT distance="150" swimtime="00:02:07.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="506" reactiontime="+80" swimtime="00:01:04.88" resultid="18432" heatid="19065" lane="7" entrytime="00:01:04.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="520" reactiontime="+72" swimtime="00:01:11.56" resultid="18433" heatid="19081" lane="3" entrytime="00:01:11.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jagoda" lastname="Roczon" birthdate="2007-01-10" gender="F" nation="POL" license="102003600066" swrid="5109134" athleteid="18394">
              <RESULTS>
                <RESULT eventid="1059" points="333" reactiontime="+76" swimtime="00:00:34.13" resultid="18395" heatid="18945" lane="7" />
                <RESULT eventid="1083" points="313" reactiontime="+76" swimtime="00:02:46.24" resultid="18396" heatid="18983" lane="9" entrytime="00:02:45.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.49" />
                    <SPLIT distance="100" swimtime="00:01:21.82" />
                    <SPLIT distance="150" swimtime="00:02:05.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="300" reactiontime="+72" swimtime="00:05:53.01" resultid="18397" heatid="19005" lane="2" entrytime="00:05:48.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                    <SPLIT distance="100" swimtime="00:01:23.05" />
                    <SPLIT distance="150" swimtime="00:02:08.50" />
                    <SPLIT distance="200" swimtime="00:02:54.78" />
                    <SPLIT distance="250" swimtime="00:03:40.72" />
                    <SPLIT distance="300" swimtime="00:04:27.11" />
                    <SPLIT distance="350" swimtime="00:05:11.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="317" reactiontime="+71" swimtime="00:01:15.79" resultid="18398" heatid="19060" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Gościński" birthdate="2007-09-23" gender="M" nation="POL" license="102003700062" swrid="5109118" athleteid="18423">
              <RESULTS>
                <RESULT eventid="1087" points="352" reactiontime="+73" swimtime="00:02:24.39" resultid="18424" heatid="18989" lane="5" entrytime="00:02:27.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                    <SPLIT distance="100" swimtime="00:01:09.60" />
                    <SPLIT distance="150" swimtime="00:01:48.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="364" reactiontime="+74" swimtime="00:05:08.16" resultid="18425" heatid="19010" lane="1" entrytime="00:05:06.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                    <SPLIT distance="100" swimtime="00:01:11.36" />
                    <SPLIT distance="150" swimtime="00:01:50.91" />
                    <SPLIT distance="200" swimtime="00:02:30.46" />
                    <SPLIT distance="250" swimtime="00:03:10.37" />
                    <SPLIT distance="300" swimtime="00:03:51.72" />
                    <SPLIT distance="350" swimtime="00:04:30.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="314" reactiontime="+73" swimtime="00:00:32.75" resultid="18426" heatid="19022" lane="6" entrytime="00:00:32.52" entrycourse="LCM" />
                <RESULT eventid="1163" points="385" reactiontime="+72" swimtime="00:01:04.43" resultid="18427" heatid="19073" lane="2" entrytime="00:01:05.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Królik" birthdate="2007-04-18" gender="M" nation="POL" license="102003700069" swrid="5109127" athleteid="18408">
              <RESULTS>
                <RESULT eventid="1063" points="273" swimtime="00:00:32.21" resultid="18409" heatid="18958" lane="9" entrytime="00:00:32.59" entrycourse="LCM" />
                <RESULT eventid="1071" points="299" reactiontime="+74" swimtime="00:00:38.78" resultid="18410" heatid="18972" lane="6" entrytime="00:00:40.59" entrycourse="LCM" />
                <RESULT eventid="1121" points="314" reactiontime="+55" swimtime="00:00:35.29" resultid="18411" heatid="19035" lane="7" entrytime="00:00:39.03" entrycourse="LCM" />
                <RESULT eventid="1137" points="289" reactiontime="+49" swimtime="00:01:26.02" resultid="18412" heatid="19046" lane="8" entrytime="00:01:27.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="312" reactiontime="+63" swimtime="00:03:05.89" resultid="18413" heatid="19093" lane="5" entrytime="00:03:11.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                    <SPLIT distance="100" swimtime="00:01:28.82" />
                    <SPLIT distance="150" swimtime="00:02:17.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Sokół" birthdate="2007-11-28" gender="M" nation="POL" license="102003700133" swrid="5109140" athleteid="18418">
              <RESULTS>
                <RESULT eventid="1063" points="228" reactiontime="+82" swimtime="00:00:34.18" resultid="18419" heatid="18956" lane="7" entrytime="00:00:35.82" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Dybowski" birthdate="2007-02-08" gender="M" nation="POL" license="102003700073" swrid="5109115" athleteid="18439">
              <RESULTS>
                <RESULT eventid="1095" points="417" reactiontime="+79" swimtime="00:02:29.70" resultid="18440" heatid="18997" lane="1" entrytime="00:02:27.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.46" />
                    <SPLIT distance="100" swimtime="00:01:12.24" />
                    <SPLIT distance="150" swimtime="00:01:51.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="393" reactiontime="+71" swimtime="00:00:32.74" resultid="18441" heatid="19036" lane="5" entrytime="00:00:33.12" entrycourse="LCM" />
                <RESULT eventid="1171" points="409" reactiontime="+91" swimtime="00:01:09.81" resultid="18442" heatid="19088" lane="8" entrytime="00:01:08.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02108" nation="POL" region="08" clubid="16851" name="AZS SMS Jarosław">
          <ATHLETES>
            <ATHLETE firstname="Kornel" lastname="Gil Amador" birthdate="2007-05-07" gender="M" nation="POL" license="102108700025" swrid="4905770" athleteid="16852">
              <RESULTS>
                <RESULT eventid="1063" points="388" reactiontime="+71" status="EXH" swimtime="00:00:28.65" resultid="16853" heatid="18960" lane="7" entrytime="00:00:28.62" entrycourse="LCM" />
                <RESULT eventid="1087" points="339" reactiontime="+72" status="EXH" swimtime="00:02:26.26" resultid="16854" heatid="18986" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                    <SPLIT distance="100" swimtime="00:01:08.32" />
                    <SPLIT distance="150" swimtime="00:01:49.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ignacy" lastname="Ożga" birthdate="2008-10-19" gender="M" nation="POL" license="102108700036" swrid="5264265" athleteid="16858">
              <RESULTS>
                <RESULT eventid="1063" points="251" status="EXH" swimtime="00:00:33.12" resultid="16859" heatid="18952" lane="0" />
                <RESULT eventid="1095" points="279" reactiontime="+73" status="EXH" swimtime="00:02:51.15" resultid="16860" heatid="18996" lane="5" entrytime="00:02:50.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                    <SPLIT distance="100" swimtime="00:01:22.51" />
                    <SPLIT distance="150" swimtime="00:02:08.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04114" nation="POL" region="14" clubid="18377" name="UKS 48 Warszawa Śródmieście">
          <ATHLETES>
            <ATHLETE firstname="Bartłomiej" lastname="Gawenda" birthdate="2006-09-13" gender="M" nation="POL" license="104114700086" swrid="5199155" athleteid="18386">
              <RESULTS>
                <RESULT eventid="1163" points="466" reactiontime="+78" status="EXH" swimtime="00:01:00.48" resultid="18387" heatid="19075" lane="6" entrytime="00:00:59.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="487" reactiontime="+83" status="EXH" swimtime="00:18:26.40" resultid="18388" heatid="19100" lane="1" entrytime="00:18:25.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                    <SPLIT distance="100" swimtime="00:01:08.53" />
                    <SPLIT distance="150" swimtime="00:01:45.14" />
                    <SPLIT distance="200" swimtime="00:02:21.80" />
                    <SPLIT distance="250" swimtime="00:02:59.50" />
                    <SPLIT distance="300" swimtime="00:03:36.11" />
                    <SPLIT distance="350" swimtime="00:04:14.31" />
                    <SPLIT distance="400" swimtime="00:04:51.21" />
                    <SPLIT distance="450" swimtime="00:05:29.15" />
                    <SPLIT distance="500" swimtime="00:06:06.00" />
                    <SPLIT distance="550" swimtime="00:06:42.97" />
                    <SPLIT distance="600" swimtime="00:07:22.85" />
                    <SPLIT distance="650" swimtime="00:08:00.29" />
                    <SPLIT distance="700" swimtime="00:08:38.31" />
                    <SPLIT distance="750" swimtime="00:09:15.60" />
                    <SPLIT distance="800" swimtime="00:09:52.42" />
                    <SPLIT distance="850" swimtime="00:10:29.42" />
                    <SPLIT distance="900" swimtime="00:11:06.57" />
                    <SPLIT distance="950" swimtime="00:11:43.49" />
                    <SPLIT distance="1000" swimtime="00:12:20.94" />
                    <SPLIT distance="1050" swimtime="00:12:57.47" />
                    <SPLIT distance="1100" swimtime="00:13:34.95" />
                    <SPLIT distance="1150" swimtime="00:14:12.22" />
                    <SPLIT distance="1200" swimtime="00:14:48.68" />
                    <SPLIT distance="1250" swimtime="00:15:25.17" />
                    <SPLIT distance="1300" swimtime="00:16:01.94" />
                    <SPLIT distance="1350" swimtime="00:16:38.57" />
                    <SPLIT distance="1400" swimtime="00:17:14.72" />
                    <SPLIT distance="1450" swimtime="00:17:51.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mikołaj" lastname="Miłkowski" birthdate="2007-03-24" gender="M" nation="POL" license="104114700075" swrid="4999446" athleteid="18378">
              <RESULTS>
                <RESULT eventid="1063" points="487" reactiontime="+73" status="EXH" swimtime="00:00:26.56" resultid="18379" heatid="18961" lane="3" entrytime="00:00:26.61" entrycourse="LCM" />
                <RESULT eventid="1079" points="510" reactiontime="+75" status="EXH" swimtime="00:01:01.93" resultid="18380" heatid="18981" lane="1" entrytime="00:01:01.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Janusz" lastname="Łazarowicz" birthdate="2007-02-22" gender="M" nation="POL" license="104114700117" swrid="5443958" athleteid="18381">
              <RESULTS>
                <RESULT eventid="1063" points="427" reactiontime="+75" status="EXH" swimtime="00:00:27.75" resultid="18382" heatid="18960" lane="3" entrytime="00:00:28.48" entrycourse="LCM" />
                <RESULT eventid="1095" points="424" reactiontime="+61" status="EXH" swimtime="00:02:28.89" resultid="18383" heatid="18997" lane="8" entrytime="00:02:29.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                    <SPLIT distance="100" swimtime="00:01:12.55" />
                    <SPLIT distance="150" swimtime="00:01:51.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="468" reactiontime="+69" status="EXH" swimtime="00:01:00.42" resultid="18384" heatid="19074" lane="3" entrytime="00:01:01.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="380" reactiontime="+76" status="EXH" swimtime="00:20:01.99" resultid="18385" heatid="19099" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                    <SPLIT distance="100" swimtime="00:01:09.63" />
                    <SPLIT distance="150" swimtime="00:01:48.01" />
                    <SPLIT distance="200" swimtime="00:02:27.32" />
                    <SPLIT distance="250" swimtime="00:03:06.78" />
                    <SPLIT distance="300" swimtime="00:03:46.00" />
                    <SPLIT distance="350" swimtime="00:04:25.32" />
                    <SPLIT distance="400" swimtime="00:05:04.81" />
                    <SPLIT distance="450" swimtime="00:05:44.44" />
                    <SPLIT distance="500" swimtime="00:06:24.06" />
                    <SPLIT distance="550" swimtime="00:07:03.94" />
                    <SPLIT distance="600" swimtime="00:07:44.06" />
                    <SPLIT distance="650" swimtime="00:08:24.50" />
                    <SPLIT distance="700" swimtime="00:09:04.61" />
                    <SPLIT distance="750" swimtime="00:09:44.35" />
                    <SPLIT distance="800" swimtime="00:10:24.42" />
                    <SPLIT distance="850" swimtime="00:11:04.73" />
                    <SPLIT distance="900" swimtime="00:11:44.15" />
                    <SPLIT distance="950" swimtime="00:12:23.49" />
                    <SPLIT distance="1000" swimtime="00:13:03.25" />
                    <SPLIT distance="1050" swimtime="00:13:50.60" />
                    <SPLIT distance="1100" swimtime="00:14:48.42" />
                    <SPLIT distance="1150" swimtime="00:15:26.36" />
                    <SPLIT distance="1200" swimtime="00:16:05.43" />
                    <SPLIT distance="1250" swimtime="00:16:45.78" />
                    <SPLIT distance="1300" swimtime="00:17:25.03" />
                    <SPLIT distance="1350" swimtime="00:18:05.46" />
                    <SPLIT distance="1400" swimtime="00:18:44.68" />
                    <SPLIT distance="1450" swimtime="00:19:23.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01003" nation="POL" region="03" clubid="18543" name="Uks Skarpa Lublin">
          <ATHLETES>
            <ATHLETE firstname="Nadia" lastname="Adamowska" birthdate="2007-12-04" gender="F" nation="POL" license="101003600265" swrid="5109150" athleteid="18568">
              <RESULTS>
                <RESULT eventid="1091" points="445" reactiontime="+63" swimtime="00:02:41.55" resultid="18569" heatid="18993" lane="3" entrytime="00:02:44.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.73" />
                    <SPLIT distance="100" swimtime="00:01:18.52" />
                    <SPLIT distance="150" swimtime="00:02:00.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="470" reactiontime="+63" swimtime="00:00:34.69" resultid="18570" heatid="19029" lane="6" entrytime="00:00:34.18" entrycourse="LCM" />
                <RESULT eventid="1167" points="435" reactiontime="+64" swimtime="00:01:15.98" resultid="18571" heatid="19081" lane="7" entrytime="00:01:14.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karol" lastname="Bronisz" birthdate="2007-10-11" gender="M" nation="POL" license="101003700236" swrid="5255418" athleteid="18548">
              <RESULTS>
                <RESULT eventid="1063" points="352" reactiontime="+48" swimtime="00:00:29.60" resultid="18549" heatid="18960" lane="0" entrytime="00:00:29.01" entrycourse="LCM" />
                <RESULT eventid="1087" points="373" reactiontime="+73" swimtime="00:02:21.68" resultid="18550" heatid="18990" lane="7" entrytime="00:02:17.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                    <SPLIT distance="100" swimtime="00:01:09.19" />
                    <SPLIT distance="150" swimtime="00:01:46.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="392" reactiontime="+72" swimtime="00:05:00.51" resultid="18551" heatid="19010" lane="2" entrytime="00:05:02.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="100" swimtime="00:01:09.66" />
                    <SPLIT distance="150" swimtime="00:01:48.43" />
                    <SPLIT distance="200" swimtime="00:02:27.63" />
                    <SPLIT distance="250" swimtime="00:03:07.19" />
                    <SPLIT distance="300" swimtime="00:03:46.22" />
                    <SPLIT distance="350" swimtime="00:04:25.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="383" reactiontime="+72" swimtime="00:01:04.57" resultid="18552" heatid="19073" lane="7" entrytime="00:01:05.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Jakubiak" birthdate="2007-05-21" gender="M" nation="POL" license="101003700244" swrid="5255458" athleteid="18553">
              <RESULTS>
                <RESULT eventid="1063" points="248" reactiontime="+68" swimtime="00:00:33.25" resultid="18554" heatid="18958" lane="8" entrytime="00:00:32.56" entrycourse="LCM" />
                <RESULT eventid="1087" points="257" reactiontime="+61" swimtime="00:02:40.34" resultid="18555" heatid="18989" lane="8" entrytime="00:02:40.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.05" />
                    <SPLIT distance="100" swimtime="00:01:16.12" />
                    <SPLIT distance="150" swimtime="00:01:58.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="251" reactiontime="+68" swimtime="00:00:35.28" resultid="18556" heatid="19022" lane="7" entrytime="00:00:35.59" entrycourse="LCM" />
                <RESULT eventid="1163" points="277" reactiontime="+72" swimtime="00:01:11.93" resultid="18557" heatid="19072" lane="1" entrytime="00:01:11.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Bartoś" birthdate="2007-09-30" gender="F" nation="POL" license="101003600232" swrid="5255357" athleteid="18544">
              <RESULTS>
                <RESULT eventid="1059" points="437" reactiontime="+77" swimtime="00:00:31.18" resultid="18545" heatid="18949" lane="1" entrytime="00:00:31.40" entrycourse="LCM" />
                <RESULT eventid="1117" points="466" reactiontime="+67" swimtime="00:00:34.80" resultid="18546" heatid="19029" lane="8" entrytime="00:00:35.27" entrycourse="LCM" />
                <RESULT eventid="1159" points="414" reactiontime="+78" swimtime="00:01:09.36" resultid="18547" heatid="19063" lane="6" entrytime="00:01:10.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paula" lastname="Brzyszko" birthdate="2007-03-23" gender="F" nation="POL" license="101003600237" swrid="5255351" athleteid="18565">
              <RESULTS>
                <RESULT eventid="1067" points="529" reactiontime="+78" swimtime="00:00:36.33" resultid="18566" heatid="18966" lane="4" entrytime="00:00:36.48" entrycourse="LCM" />
                <RESULT eventid="1133" points="485" swimtime="00:01:21.61" resultid="18567" heatid="19041" lane="0" entrytime="00:01:20.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Rybczyński" birthdate="2008-05-09" gender="M" nation="POL" license="101003700256" swrid="5113670" athleteid="18563">
              <RESULTS>
                <RESULT eventid="1063" points="398" reactiontime="+59" swimtime="00:00:28.42" resultid="18564" heatid="18960" lane="6" entrytime="00:00:28.55" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Winiarczyk" birthdate="2007-03-23" gender="M" nation="POL" license="101003700261" swrid="5280817" athleteid="18558">
              <RESULTS>
                <RESULT eventid="1063" points="246" swimtime="00:00:33.35" resultid="18559" heatid="18957" lane="3" entrytime="00:00:33.41" entrycourse="LCM" />
                <RESULT eventid="1071" points="208" swimtime="00:00:43.76" resultid="18560" heatid="18971" lane="7" entrytime="00:00:44.19" entrycourse="LCM" />
                <RESULT eventid="1137" points="218" reactiontime="+99" swimtime="00:01:34.38" resultid="18561" heatid="19045" lane="7" entrytime="00:01:35.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="260" swimtime="00:01:13.43" resultid="18562" heatid="19072" lane="9" entrytime="00:01:12.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01403" nation="POL" region="03" clubid="16907" name="KS ,,OLIMPIA&apos;&apos; Lublin">
          <ATHLETES>
            <ATHLETE firstname="Nicholai" lastname="Wysmulski" birthdate="2006-09-09" gender="M" nation="POL" license="101403700100" swrid="5019843" athleteid="16954">
              <RESULTS>
                <RESULT eventid="1063" points="443" reactiontime="+56" swimtime="00:00:27.42" resultid="16955" heatid="18960" lane="2" entrytime="00:00:28.57" entrycourse="LCM" />
                <RESULT eventid="1113" points="433" reactiontime="+57" swimtime="00:00:29.42" resultid="16956" heatid="19023" lane="2" entrytime="00:00:30.43" entrycourse="LCM" />
                <RESULT eventid="1137" points="380" reactiontime="+75" swimtime="00:01:18.52" resultid="16957" heatid="19042" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Iga" lastname="Rumińska" birthdate="2007-09-05" gender="F" nation="POL" license="101403600173" swrid="5109135" athleteid="17001">
              <RESULTS>
                <RESULT eventid="1067" points="393" reactiontime="+74" swimtime="00:00:40.13" resultid="17002" heatid="18966" lane="8" entrytime="00:00:42.65" entrycourse="LCM" />
                <RESULT eventid="1083" points="389" reactiontime="+80" swimtime="00:02:34.68" resultid="17003" heatid="18983" lane="2" entrytime="00:02:32.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                    <SPLIT distance="100" swimtime="00:01:16.05" />
                    <SPLIT distance="150" swimtime="00:01:56.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="336" reactiontime="+80" swimtime="00:01:32.17" resultid="17004" heatid="19040" lane="1" entrytime="00:01:32.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="433" reactiontime="+76" swimtime="00:01:08.32" resultid="17005" heatid="19063" lane="5" entrytime="00:01:08.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Daniel" birthdate="2006-08-31" gender="M" nation="POL" license="101403700084" swrid="4936956" athleteid="17016">
              <RESULTS>
                <RESULT eventid="1071" points="312" reactiontime="+67" swimtime="00:00:38.24" resultid="17017" heatid="18973" lane="2" entrytime="00:00:37.42" entrycourse="LCM" />
                <RESULT eventid="1137" points="327" reactiontime="+68" swimtime="00:01:22.50" resultid="17018" heatid="19046" lane="6" entrytime="00:01:23.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="340" reactiontime="+68" swimtime="00:01:07.17" resultid="17019" heatid="19073" lane="9" entrytime="00:01:07.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patrycja" lastname="Ciećko" birthdate="2005-07-08" gender="F" nation="POL" license="101403600210" swrid="4996867" athleteid="16924">
              <RESULTS>
                <RESULT eventid="1059" points="431" reactiontime="+58" swimtime="00:00:31.33" resultid="16925" heatid="18949" lane="2" entrytime="00:00:31.06" entrycourse="LCM" />
                <RESULT eventid="1117" points="481" reactiontime="+81" swimtime="00:00:34.42" resultid="16926" heatid="19029" lane="7" entrytime="00:00:34.58" entrycourse="LCM" />
                <RESULT eventid="1159" points="404" reactiontime="+78" swimtime="00:01:09.93" resultid="16927" heatid="19063" lane="0" entrytime="00:01:12.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="430" reactiontime="+80" swimtime="00:01:16.25" resultid="16928" heatid="19081" lane="1" entrytime="00:01:15.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Stempurski" birthdate="2004-09-30" gender="M" nation="POL" license="101403700153" swrid="5233337" athleteid="16968">
              <RESULTS>
                <RESULT eventid="1063" points="488" reactiontime="+70" swimtime="00:00:26.55" resultid="16969" heatid="18961" lane="5" entrytime="00:00:26.59" entrycourse="LCM" />
                <RESULT eventid="1095" points="459" reactiontime="+66" swimtime="00:02:25.04" resultid="16970" heatid="18997" lane="7" entrytime="00:02:25.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                    <SPLIT distance="100" swimtime="00:01:10.86" />
                    <SPLIT distance="150" swimtime="00:01:48.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="494" reactiontime="+64" swimtime="00:00:28.16" resultid="16971" heatid="19024" lane="2" entrytime="00:00:28.13" entrycourse="LCM" />
                <RESULT eventid="1121" points="455" reactiontime="+70" swimtime="00:00:31.19" resultid="16972" heatid="19033" lane="0" />
                <RESULT eventid="1163" points="530" reactiontime="+70" swimtime="00:00:57.94" resultid="16973" heatid="19076" lane="8" entrytime="00:00:57.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="428" reactiontime="+62" swimtime="00:01:08.78" resultid="16974" heatid="19083" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Zuzaniuk" birthdate="2004-07-06" gender="M" nation="POL" license="101403700068" swrid="4744904" athleteid="17011">
              <RESULTS>
                <RESULT eventid="1071" points="551" reactiontime="+66" swimtime="00:00:31.64" resultid="17012" heatid="18974" lane="1" entrytime="00:00:32.48" entrycourse="LCM" />
                <RESULT eventid="1103" points="560" reactiontime="+66" swimtime="00:04:55.77" resultid="17013" heatid="19001" lane="5" entrytime="00:04:52.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.10" />
                    <SPLIT distance="100" swimtime="00:01:06.08" />
                    <SPLIT distance="150" swimtime="00:01:44.37" />
                    <SPLIT distance="200" swimtime="00:02:21.64" />
                    <SPLIT distance="250" swimtime="00:03:03.85" />
                    <SPLIT distance="300" swimtime="00:03:44.91" />
                    <SPLIT distance="350" swimtime="00:04:20.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="527" reactiontime="+68" swimtime="00:02:21.08" resultid="17014" heatid="19054" lane="6" entrytime="00:02:17.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.45" />
                    <SPLIT distance="100" swimtime="00:01:06.21" />
                    <SPLIT distance="150" swimtime="00:01:47.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="513" reactiontime="+65" swimtime="00:00:58.57" resultid="17015" heatid="19076" lane="6" entrytime="00:00:57.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Panasiuk" birthdate="2005-03-28" gender="F" nation="POL" license="101403600208" swrid="4917601" athleteid="17036">
              <RESULTS>
                <RESULT eventid="1075" points="433" reactiontime="+84" swimtime="00:01:13.28" resultid="17037" heatid="18976" lane="1" entrytime="00:01:16.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="483" reactiontime="+82" swimtime="00:02:23.96" resultid="17038" heatid="18982" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                    <SPLIT distance="100" swimtime="00:01:10.73" />
                    <SPLIT distance="150" swimtime="00:01:48.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="423" reactiontime="+80" swimtime="00:00:32.53" resultid="17039" heatid="19016" lane="8" entrytime="00:00:33.44" entrycourse="LCM" />
                <RESULT eventid="1117" points="436" reactiontime="+78" swimtime="00:00:35.58" resultid="17040" heatid="19028" lane="4" entrytime="00:00:35.89" entrycourse="LCM" />
                <RESULT eventid="1159" points="472" reactiontime="+84" swimtime="00:01:06.40" resultid="17041" heatid="19064" lane="2" entrytime="00:01:07.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Kawecki" birthdate="2008-07-14" gender="M" nation="POL" license="101403700205" swrid="5453704" athleteid="16944">
              <RESULTS>
                <RESULT eventid="1063" points="188" reactiontime="+81" swimtime="00:00:36.48" resultid="16945" heatid="18952" lane="4" />
                <RESULT eventid="1121" points="157" reactiontime="+73" swimtime="00:00:44.42" resultid="16946" heatid="19031" lane="2" />
                <RESULT eventid="1163" points="215" reactiontime="+93" swimtime="00:01:18.23" resultid="16947" heatid="19069" lane="3" entrytime="00:01:24.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="190" reactiontime="+81" swimtime="00:01:30.13" resultid="16948" heatid="19084" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pola" lastname="Kędzior" birthdate="2007-01-10" gender="F" nation="POL" license="101403600137" swrid="4621831" athleteid="17071">
              <RESULTS>
                <RESULT eventid="1099" points="565" reactiontime="+74" swimtime="00:05:22.19" resultid="17072" heatid="18999" lane="2" entrytime="00:05:23.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.03" />
                    <SPLIT distance="100" swimtime="00:01:12.00" />
                    <SPLIT distance="150" swimtime="00:01:54.42" />
                    <SPLIT distance="200" swimtime="00:02:35.49" />
                    <SPLIT distance="250" swimtime="00:03:22.50" />
                    <SPLIT distance="300" swimtime="00:04:08.25" />
                    <SPLIT distance="350" swimtime="00:04:45.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="566" reactiontime="+54" swimtime="00:02:32.39" resultid="17073" heatid="19050" lane="8" entrytime="00:02:33.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.61" />
                    <SPLIT distance="100" swimtime="00:01:12.60" />
                    <SPLIT distance="150" swimtime="00:01:58.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1150" points="507" reactiontime="+79" swimtime="00:02:32.75" resultid="17074" heatid="19057" lane="2" entrytime="00:02:36.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.69" />
                    <SPLIT distance="100" swimtime="00:01:13.69" />
                    <SPLIT distance="150" swimtime="00:01:53.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="511" reactiontime="+73" swimtime="00:02:54.00" resultid="17075" heatid="19089" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.52" />
                    <SPLIT distance="100" swimtime="00:01:24.84" />
                    <SPLIT distance="150" swimtime="00:02:10.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksander" lastname="Ciepałowicz" birthdate="2008-02-27" gender="M" nation="POL" license="101403700116" swrid="5098720" athleteid="16958">
              <RESULTS>
                <RESULT eventid="1063" points="295" reactiontime="+86" swimtime="00:00:31.41" resultid="16959" heatid="18959" lane="1" entrytime="00:00:31.02" entrycourse="LCM" />
                <RESULT eventid="1087" points="284" reactiontime="+77" swimtime="00:02:35.10" resultid="16960" heatid="18989" lane="7" entrytime="00:02:38.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                    <SPLIT distance="100" swimtime="00:01:14.70" />
                    <SPLIT distance="150" swimtime="00:01:56.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1137" points="247" reactiontime="+73" swimtime="00:01:30.63" resultid="16961" heatid="19046" lane="0" entrytime="00:01:31.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="325" reactiontime="+70" swimtime="00:01:08.19" resultid="16962" heatid="19072" lane="3" entrytime="00:01:10.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ernest" lastname="Szychiewicz" birthdate="2004-04-16" gender="M" nation="POL" license="101403700193" swrid="5204715" athleteid="16981">
              <RESULTS>
                <RESULT eventid="1063" points="506" reactiontime="+70" swimtime="00:00:26.24" resultid="16982" heatid="18952" lane="3" />
                <RESULT eventid="1079" points="493" reactiontime="+77" swimtime="00:01:02.65" resultid="16983" heatid="18981" lane="7" entrytime="00:01:01.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1087" points="498" reactiontime="+74" swimtime="00:02:08.66" resultid="16984" heatid="18991" lane="8" entrytime="00:02:03.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.33" />
                    <SPLIT distance="100" swimtime="00:01:01.91" />
                    <SPLIT distance="150" swimtime="00:01:35.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="553" reactiontime="+75" swimtime="00:04:28.02" resultid="16985" heatid="19011" lane="2" entrytime="00:04:29.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                    <SPLIT distance="100" swimtime="00:01:03.45" />
                    <SPLIT distance="150" swimtime="00:01:37.01" />
                    <SPLIT distance="200" swimtime="00:02:11.34" />
                    <SPLIT distance="250" swimtime="00:02:45.76" />
                    <SPLIT distance="300" swimtime="00:03:20.18" />
                    <SPLIT distance="350" swimtime="00:03:54.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="445" reactiontime="+70" swimtime="00:00:29.15" resultid="16986" heatid="19024" lane="8" entrytime="00:00:28.54" entrycourse="LCM" />
                <RESULT eventid="1155" points="487" reactiontime="+76" swimtime="00:02:20.71" resultid="16987" heatid="19059" lane="3" entrytime="00:02:16.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.15" />
                    <SPLIT distance="100" swimtime="00:01:05.63" />
                    <SPLIT distance="150" swimtime="00:01:42.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="487" reactiontime="+74" swimtime="00:00:59.59" resultid="16988" heatid="19076" lane="2" entrytime="00:00:57.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tymon" lastname="Mrówczyński" birthdate="2008-11-14" gender="M" nation="POL" license="101403700198" swrid="5453740" athleteid="16963">
              <RESULTS>
                <RESULT eventid="1063" points="213" reactiontime="+68" swimtime="00:00:34.97" resultid="16964" heatid="18955" lane="4" entrytime="00:00:37.66" entrycourse="LCM" />
                <RESULT eventid="1071" points="171" reactiontime="+93" swimtime="00:00:46.68" resultid="16965" heatid="18969" lane="8" />
                <RESULT comment="K4 - Pływak wykonał cykl ruchowy inny niż jeden ruch ramion i jedno kopnięcie nogami (z wyjątkiem ostatniego cyklu przed nawrotem lub zakończeniem wyścigu)" eventid="1137" reactiontime="+82" status="DSQ" swimtime="00:01:43.81" resultid="16966" heatid="19042" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.45" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej, a przed sygnałem startu" eventid="1163" reactiontime="+61" status="DSQ" swimtime="00:01:19.73" resultid="16967" heatid="19069" lane="1" entrytime="00:01:27.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amelia" lastname="Grabowska" birthdate="2007-01-29" gender="F" nation="POL" license="101403600140" swrid="5109080" athleteid="17042">
              <RESULTS>
                <RESULT eventid="1075" points="409" reactiontime="+72" swimtime="00:01:14.72" resultid="17043" heatid="18976" lane="6" entrytime="00:01:13.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="411" reactiontime="+74" swimtime="00:05:17.93" resultid="17044" heatid="19005" lane="5" entrytime="00:05:20.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.37" />
                    <SPLIT distance="100" swimtime="00:01:11.93" />
                    <SPLIT distance="150" swimtime="00:01:51.96" />
                    <SPLIT distance="200" swimtime="00:02:32.60" />
                    <SPLIT distance="250" swimtime="00:03:13.87" />
                    <SPLIT distance="300" swimtime="00:03:55.02" />
                    <SPLIT distance="350" swimtime="00:04:36.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="423" reactiontime="+71" swimtime="00:00:32.53" resultid="17045" heatid="19015" lane="4" entrytime="00:00:35.08" entrycourse="LCM" />
                <RESULT eventid="1167" points="463" reactiontime="+74" swimtime="00:01:14.38" resultid="17046" heatid="19079" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="366" reactiontime="+74" swimtime="00:11:17.62" resultid="17047" heatid="19095" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.51" />
                    <SPLIT distance="100" swimtime="00:01:17.59" />
                    <SPLIT distance="150" swimtime="00:02:00.12" />
                    <SPLIT distance="200" swimtime="00:02:42.90" />
                    <SPLIT distance="250" swimtime="00:03:25.90" />
                    <SPLIT distance="300" swimtime="00:04:08.52" />
                    <SPLIT distance="350" swimtime="00:04:51.66" />
                    <SPLIT distance="400" swimtime="00:05:34.82" />
                    <SPLIT distance="450" swimtime="00:06:18.71" />
                    <SPLIT distance="500" swimtime="00:07:01.81" />
                    <SPLIT distance="550" swimtime="00:07:45.57" />
                    <SPLIT distance="600" swimtime="00:08:28.94" />
                    <SPLIT distance="650" swimtime="00:09:12.54" />
                    <SPLIT distance="700" swimtime="00:09:55.01" />
                    <SPLIT distance="750" swimtime="00:10:37.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emil" lastname="Zieliński" birthdate="2006-02-13" gender="M" nation="POL" license="101403700192" swrid="4901077" athleteid="16975">
              <RESULTS>
                <RESULT eventid="1063" points="485" reactiontime="+69" swimtime="00:00:26.60" resultid="16976" heatid="18961" lane="7" entrytime="00:00:26.77" entrycourse="LCM" />
                <RESULT eventid="1071" points="418" reactiontime="+72" swimtime="00:00:34.70" resultid="16977" heatid="18973" lane="5" entrytime="00:00:35.30" entrycourse="LCM" />
                <RESULT eventid="1121" points="431" reactiontime="+70" swimtime="00:00:31.76" resultid="16978" heatid="19037" lane="8" entrytime="00:00:31.41" entrycourse="LCM" />
                <RESULT eventid="1137" points="332" reactiontime="+74" swimtime="00:01:22.13" resultid="16979" heatid="19043" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="441" reactiontime="+73" swimtime="00:01:01.62" resultid="16980" heatid="19074" lane="4" entrytime="00:01:00.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Magdalena" lastname="Mituła" birthdate="2004-09-21" gender="F" nation="POL" license="101403600105" swrid="4892154" athleteid="16929">
              <RESULTS>
                <RESULT eventid="1059" points="459" reactiontime="+63" swimtime="00:00:30.67" resultid="16930" heatid="18950" lane="0" entrytime="00:00:30.19" entrycourse="LCM" />
                <RESULT eventid="1083" points="431" reactiontime="+67" swimtime="00:02:29.49" resultid="16931" heatid="18984" lane="0" entrytime="00:02:27.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                    <SPLIT distance="100" swimtime="00:01:12.93" />
                    <SPLIT distance="150" swimtime="00:01:51.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="401" reactiontime="+67" swimtime="00:05:20.41" resultid="16932" heatid="19006" lane="0" entrytime="00:05:17.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                    <SPLIT distance="100" swimtime="00:01:15.40" />
                    <SPLIT distance="150" swimtime="00:01:56.58" />
                    <SPLIT distance="200" swimtime="00:02:37.62" />
                    <SPLIT distance="250" swimtime="00:03:18.87" />
                    <SPLIT distance="300" swimtime="00:04:00.48" />
                    <SPLIT distance="350" swimtime="00:04:41.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="436" reactiontime="+67" swimtime="00:01:08.18" resultid="16933" heatid="19064" lane="7" entrytime="00:01:07.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Szemro" birthdate="2008-06-20" gender="M" nation="POL" license="101403700180" swrid="5387648" athleteid="17006">
              <RESULTS>
                <RESULT eventid="1071" points="157" reactiontime="+75" swimtime="00:00:48.01" resultid="17007" heatid="18970" lane="6" entrytime="00:00:49.28" entrycourse="LCM" />
                <RESULT eventid="1087" points="210" reactiontime="+78" swimtime="00:02:51.38" resultid="17008" heatid="18988" lane="5" entrytime="00:02:50.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                    <SPLIT distance="100" swimtime="00:01:22.68" />
                    <SPLIT distance="150" swimtime="00:02:08.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="178" reactiontime="+88" swimtime="00:00:42.65" resultid="17009" heatid="19031" lane="4" />
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej, a przed sygnałem startu" eventid="1137" reactiontime="+58" status="DSQ" swimtime="00:01:44.36" resultid="17010" heatid="19044" lane="2" entrytime="00:01:42.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emilia" lastname="Nowoświatłowska" birthdate="2007-09-16" gender="F" nation="POL" license="101403600181" swrid="5387647" athleteid="16920">
              <RESULTS>
                <RESULT eventid="1059" points="446" reactiontime="+75" swimtime="00:00:30.98" resultid="16921" heatid="18949" lane="5" entrytime="00:00:30.53" entrycourse="LCM" />
                <RESULT eventid="1108" points="320" reactiontime="+76" swimtime="00:00:35.68" resultid="16922" heatid="19015" lane="5" entrytime="00:00:35.25" entrycourse="LCM" />
                <RESULT eventid="1159" points="479" reactiontime="+69" swimtime="00:01:06.08" resultid="16923" heatid="19064" lane="5" entrytime="00:01:06.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonina" lastname="Siek" birthdate="2008-02-14" gender="F" nation="POL" license="101403600160" swrid="5285778" athleteid="16994">
              <RESULTS>
                <RESULT eventid="1067" points="314" swimtime="00:00:43.25" resultid="16995" heatid="18966" lane="9" entrytime="00:00:43.90" entrycourse="LCM" />
                <RESULT eventid="1075" points="359" swimtime="00:01:17.99" resultid="16996" heatid="18976" lane="8" entrytime="00:01:17.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="425" reactiontime="+63" swimtime="00:05:14.50" resultid="16997" heatid="19005" lane="4" entrytime="00:05:19.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                    <SPLIT distance="100" swimtime="00:01:13.37" />
                    <SPLIT distance="150" swimtime="00:01:54.10" />
                    <SPLIT distance="200" swimtime="00:02:35.10" />
                    <SPLIT distance="250" swimtime="00:03:16.05" />
                    <SPLIT distance="300" swimtime="00:03:56.24" />
                    <SPLIT distance="350" swimtime="00:04:35.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="331" swimtime="00:00:35.31" resultid="16998" heatid="19016" lane="9" entrytime="00:00:34.78" entrycourse="LCM" />
                <RESULT eventid="1175" points="361" reactiontime="+73" swimtime="00:03:15.36" resultid="16999" heatid="19090" lane="3" entrytime="00:03:18.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.87" />
                    <SPLIT distance="100" swimtime="00:01:32.53" />
                    <SPLIT distance="150" swimtime="00:02:23.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="415" swimtime="00:10:49.75" resultid="17000" heatid="19096" lane="5" entrytime="00:10:55.47" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Danilewicz" birthdate="2007-08-10" gender="F" nation="POL" license="101403600156" swrid="5109112" athleteid="17025">
              <RESULTS>
                <RESULT eventid="1075" points="499" reactiontime="+72" swimtime="00:01:09.93" resultid="17026" heatid="18975" lane="5" entrytime="00:01:23.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1091" points="512" reactiontime="+73" swimtime="00:02:34.18" resultid="17027" heatid="18993" lane="4" entrytime="00:02:37.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.56" />
                    <SPLIT distance="100" swimtime="00:01:16.60" />
                    <SPLIT distance="150" swimtime="00:01:56.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="521" reactiontime="+62" swimtime="00:00:30.36" resultid="17028" heatid="19017" lane="1" entrytime="00:00:30.53" entrycourse="LCM" />
                <RESULT eventid="1117" points="579" reactiontime="+74" swimtime="00:00:32.37" resultid="17029" heatid="19030" lane="0" entrytime="00:00:32.75" entrycourse="LCM" />
                <RESULT eventid="1167" points="568" reactiontime="+71" swimtime="00:01:09.51" resultid="17030" heatid="19082" lane="9" entrytime="00:01:09.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julianna" lastname="Wyrwas" birthdate="2008-07-12" gender="F" nation="POL" license="101403600179" swrid="5148618" athleteid="16914">
              <RESULTS>
                <RESULT eventid="1059" points="489" reactiontime="+60" swimtime="00:00:30.03" resultid="16915" heatid="18950" lane="8" entrytime="00:00:30.14" entrycourse="LCM" />
                <RESULT eventid="1083" points="419" reactiontime="+61" swimtime="00:02:30.88" resultid="16916" heatid="18983" lane="5" entrytime="00:02:29.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.99" />
                    <SPLIT distance="100" swimtime="00:01:16.78" />
                    <SPLIT distance="150" swimtime="00:01:56.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="415" reactiontime="+77" swimtime="00:00:36.16" resultid="16917" heatid="19028" lane="5" entrytime="00:00:36.12" entrycourse="LCM" />
                <RESULT eventid="1159" points="482" reactiontime="+76" swimtime="00:01:05.91" resultid="16918" heatid="19064" lane="4" entrytime="00:01:06.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="386" reactiontime="+77" swimtime="00:01:19.01" resultid="16919" heatid="19078" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwia" lastname="Grączak" birthdate="2008-06-18" gender="F" nation="POL" license="101403600157" swrid="5158155" athleteid="17065">
              <RESULTS>
                <RESULT eventid="1091" points="556" reactiontime="+91" swimtime="00:02:29.98" resultid="17066" heatid="18994" lane="0" entrytime="00:02:32.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                    <SPLIT distance="100" swimtime="00:01:12.91" />
                    <SPLIT distance="150" swimtime="00:01:52.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="534" reactiontime="+87" swimtime="00:00:33.24" resultid="17067" heatid="19030" lane="9" entrytime="00:00:32.81" entrycourse="LCM" />
                <RESULT eventid="1141" points="488" reactiontime="+81" swimtime="00:02:40.10" resultid="17068" heatid="19049" lane="4" entrytime="00:02:39.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.91" />
                    <SPLIT distance="100" swimtime="00:01:14.96" />
                    <SPLIT distance="150" swimtime="00:02:02.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1150" points="412" reactiontime="+99" swimtime="00:02:43.67" resultid="17069" heatid="19057" lane="1" entrytime="00:02:47.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.13" />
                    <SPLIT distance="100" swimtime="00:01:16.50" />
                    <SPLIT distance="150" swimtime="00:02:00.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="545" reactiontime="+81" swimtime="00:01:10.44" resultid="17070" heatid="19081" lane="5" entrytime="00:01:10.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rozalia" lastname="Turska" birthdate="2007-11-03" gender="F" nation="POL" license="101403600161" swrid="5045346" athleteid="17031">
              <RESULTS>
                <RESULT eventid="1075" points="345" reactiontime="+70" swimtime="00:01:19.05" resultid="17032" heatid="18976" lane="9" entrytime="00:01:21.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="384" swimtime="00:00:33.59" resultid="17033" heatid="19016" lane="0" entrytime="00:00:34.39" entrycourse="LCM" />
                <RESULT eventid="1133" points="359" reactiontime="+59" swimtime="00:01:30.20" resultid="17034" heatid="19040" lane="8" entrytime="00:01:33.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.25" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="M5 - Pływak nie przeniósł ramion do przodu nad lustrem wody" eventid="1150" reactiontime="+67" status="DSQ" swimtime="00:03:13.08" resultid="17035" heatid="19056" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.80" />
                    <SPLIT distance="100" swimtime="00:01:27.76" />
                    <SPLIT distance="150" swimtime="00:02:16.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kamila" lastname="Bielak" birthdate="2008-01-02" gender="F" nation="POL" license="101403600162" swrid="5109074" athleteid="16989">
              <RESULTS>
                <RESULT eventid="1067" points="495" reactiontime="+55" swimtime="00:00:37.16" resultid="16990" heatid="18967" lane="0" entrytime="00:00:36.27" entrycourse="LCM" />
                <RESULT eventid="1083" points="421" reactiontime="+72" swimtime="00:02:30.68" resultid="16991" heatid="18983" lane="6" entrytime="00:02:32.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.10" />
                    <SPLIT distance="100" swimtime="00:01:14.49" />
                    <SPLIT distance="150" swimtime="00:01:53.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="474" reactiontime="+74" swimtime="00:01:22.24" resultid="16992" heatid="19041" lane="7" entrytime="00:01:19.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="458" reactiontime="+73" swimtime="00:03:00.35" resultid="16993" heatid="19091" lane="9" entrytime="00:02:58.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.94" />
                    <SPLIT distance="100" swimtime="00:01:27.57" />
                    <SPLIT distance="150" swimtime="00:02:14.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Dragan" birthdate="2004-07-16" gender="F" nation="POL" license="101403600131" swrid="4744917" athleteid="17054">
              <RESULTS>
                <RESULT eventid="1083" points="636" reactiontime="+80" swimtime="00:02:11.31" resultid="17055" heatid="18985" lane="2" entrytime="00:02:12.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.28" />
                    <SPLIT distance="100" swimtime="00:01:03.85" />
                    <SPLIT distance="150" swimtime="00:01:38.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="622" reactiontime="+85" swimtime="00:05:11.95" resultid="17056" heatid="18999" lane="3" entrytime="00:05:11.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.35" />
                    <SPLIT distance="100" swimtime="00:01:14.13" />
                    <SPLIT distance="150" swimtime="00:01:54.48" />
                    <SPLIT distance="200" swimtime="00:02:34.69" />
                    <SPLIT distance="250" swimtime="00:03:19.51" />
                    <SPLIT distance="300" swimtime="00:04:03.65" />
                    <SPLIT distance="350" swimtime="00:04:38.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="600" reactiontime="+83" swimtime="00:02:29.52" resultid="17057" heatid="19050" lane="2" entrytime="00:02:28.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                    <SPLIT distance="100" swimtime="00:01:12.50" />
                    <SPLIT distance="150" swimtime="00:01:56.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="586" reactiontime="+75" swimtime="00:01:01.78" resultid="17058" heatid="19065" lane="4" entrytime="00:01:02.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Serga" birthdate="2003-06-14" gender="M" nation="POL" license="101403700172" swrid="5345125" athleteid="17020">
              <RESULTS>
                <RESULT eventid="1071" points="572" reactiontime="+66" swimtime="00:00:31.25" resultid="17021" heatid="18974" lane="6" entrytime="00:00:31.11" entrycourse="LCM" />
                <RESULT eventid="1113" points="533" reactiontime="+67" swimtime="00:00:27.46" resultid="17022" heatid="19024" lane="5" entrytime="00:00:27.64" entrycourse="LCM" />
                <RESULT eventid="1137" points="548" reactiontime="+67" swimtime="00:01:09.49" resultid="17023" heatid="19047" lane="3" entrytime="00:01:09.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="539" reactiontime="+72" swimtime="00:02:34.96" resultid="17024" heatid="19094" lane="5" entrytime="00:02:33.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.88" />
                    <SPLIT distance="100" swimtime="00:01:12.98" />
                    <SPLIT distance="150" swimtime="00:01:54.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwier" lastname="Ponieważ" birthdate="2007-02-03" gender="M" nation="POL" license="101403700096" swrid="5098718" athleteid="17059">
              <RESULTS>
                <RESULT eventid="1087" points="522" reactiontime="+74" swimtime="00:02:06.67" resultid="17060" heatid="18991" lane="9" entrytime="00:02:05.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.75" />
                    <SPLIT distance="100" swimtime="00:01:02.54" />
                    <SPLIT distance="150" swimtime="00:01:35.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6365" points="517" reactiontime="+77" swimtime="00:09:23.28" resultid="17061" heatid="19003" lane="9" entrytime="00:09:45.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.55" />
                    <SPLIT distance="100" swimtime="00:01:06.21" />
                    <SPLIT distance="150" swimtime="00:01:41.36" />
                    <SPLIT distance="200" swimtime="00:02:17.11" />
                    <SPLIT distance="250" swimtime="00:02:53.42" />
                    <SPLIT distance="300" swimtime="00:03:29.24" />
                    <SPLIT distance="350" swimtime="00:04:05.06" />
                    <SPLIT distance="400" swimtime="00:04:42.02" />
                    <SPLIT distance="450" swimtime="00:05:17.89" />
                    <SPLIT distance="500" swimtime="00:05:54.00" />
                    <SPLIT distance="550" swimtime="00:06:29.92" />
                    <SPLIT distance="600" swimtime="00:07:05.22" />
                    <SPLIT distance="650" swimtime="00:07:40.47" />
                    <SPLIT distance="700" swimtime="00:08:15.07" />
                    <SPLIT distance="750" swimtime="00:08:49.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="568" reactiontime="+77" swimtime="00:04:25.64" resultid="17062" heatid="19011" lane="6" entrytime="00:04:28.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.58" />
                    <SPLIT distance="100" swimtime="00:01:04.20" />
                    <SPLIT distance="150" swimtime="00:01:38.00" />
                    <SPLIT distance="200" swimtime="00:02:11.58" />
                    <SPLIT distance="250" swimtime="00:02:45.51" />
                    <SPLIT distance="300" swimtime="00:03:20.37" />
                    <SPLIT distance="350" swimtime="00:03:54.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="370" reactiontime="+82" swimtime="00:01:05.31" resultid="17063" heatid="19076" lane="0" entrytime="00:00:58.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="558" reactiontime="+84" swimtime="00:17:37.38" resultid="17064" heatid="19100" lane="2" entrytime="00:18:13.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                    <SPLIT distance="100" swimtime="00:01:08.83" />
                    <SPLIT distance="150" swimtime="00:01:43.81" />
                    <SPLIT distance="200" swimtime="00:02:19.44" />
                    <SPLIT distance="250" swimtime="00:02:55.05" />
                    <SPLIT distance="300" swimtime="00:03:30.58" />
                    <SPLIT distance="350" swimtime="00:04:06.42" />
                    <SPLIT distance="400" swimtime="00:04:41.86" />
                    <SPLIT distance="450" swimtime="00:05:18.33" />
                    <SPLIT distance="500" swimtime="00:05:54.03" />
                    <SPLIT distance="550" swimtime="00:06:29.95" />
                    <SPLIT distance="600" swimtime="00:07:06.14" />
                    <SPLIT distance="650" swimtime="00:07:42.77" />
                    <SPLIT distance="700" swimtime="00:08:18.31" />
                    <SPLIT distance="750" swimtime="00:08:54.25" />
                    <SPLIT distance="800" swimtime="00:09:29.94" />
                    <SPLIT distance="850" swimtime="00:10:05.73" />
                    <SPLIT distance="900" swimtime="00:10:41.58" />
                    <SPLIT distance="950" swimtime="00:11:16.76" />
                    <SPLIT distance="1000" swimtime="00:11:50.78" />
                    <SPLIT distance="1050" swimtime="00:12:25.32" />
                    <SPLIT distance="1100" swimtime="00:13:00.30" />
                    <SPLIT distance="1150" swimtime="00:13:36.14" />
                    <SPLIT distance="1200" swimtime="00:14:11.99" />
                    <SPLIT distance="1250" swimtime="00:14:47.26" />
                    <SPLIT distance="1300" swimtime="00:15:21.97" />
                    <SPLIT distance="1350" swimtime="00:15:57.13" />
                    <SPLIT distance="1400" swimtime="00:16:31.32" />
                    <SPLIT distance="1450" swimtime="00:17:05.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miłosz" lastname="Tama-Poniatowski" birthdate="2007-04-09" gender="M" nation="POL" license="101403700169" swrid="5323850" athleteid="16949">
              <RESULTS>
                <RESULT eventid="1063" points="354" reactiontime="+72" swimtime="00:00:29.54" resultid="16950" heatid="18959" lane="8" entrytime="00:00:31.05" entrycourse="LCM" />
                <RESULT eventid="1071" points="327" reactiontime="+66" swimtime="00:00:37.63" resultid="16951" heatid="18973" lane="0" entrytime="00:00:37.89" entrycourse="LCM" />
                <RESULT eventid="1113" points="276" reactiontime="+69" swimtime="00:00:34.20" resultid="16952" heatid="19019" lane="4" />
                <RESULT eventid="1121" points="281" reactiontime="+72" swimtime="00:00:36.63" resultid="16953" heatid="19032" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Klaudia" lastname="Kazanowska" birthdate="2008-03-05" gender="F" nation="POL" license="101403600202" swrid="5193104" athleteid="16908">
              <RESULTS>
                <RESULT eventid="1059" points="505" swimtime="00:00:29.71" resultid="16909" heatid="18950" lane="2" entrytime="00:00:29.65" entrycourse="LCM" />
                <RESULT eventid="1083" points="465" reactiontime="+75" swimtime="00:02:25.81" resultid="16910" heatid="18984" lane="9" entrytime="00:02:27.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                    <SPLIT distance="100" swimtime="00:01:10.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="456" reactiontime="+73" swimtime="00:00:35.05" resultid="16911" heatid="19029" lane="1" entrytime="00:00:35.16" entrycourse="LCM" />
                <RESULT eventid="1159" points="504" reactiontime="+75" swimtime="00:01:04.95" resultid="16912" heatid="19064" lane="3" entrytime="00:01:06.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="426" reactiontime="+80" swimtime="00:01:16.46" resultid="16913" heatid="19080" lane="4" entrytime="00:01:21.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Kozak" birthdate="2006-11-13" gender="M" nation="POL" license="101403700120" swrid="5109083" athleteid="17048">
              <RESULTS>
                <RESULT eventid="1079" points="390" reactiontime="+69" swimtime="00:01:07.71" resultid="17049" heatid="18980" lane="2" entrytime="00:01:06.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6365" points="417" reactiontime="+68" swimtime="00:10:04.91" resultid="17050" heatid="19002" lane="4" entrytime="00:09:45.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                    <SPLIT distance="100" swimtime="00:01:09.51" />
                    <SPLIT distance="150" swimtime="00:01:46.03" />
                    <SPLIT distance="200" swimtime="00:02:22.34" />
                    <SPLIT distance="250" swimtime="00:02:59.21" />
                    <SPLIT distance="300" swimtime="00:03:37.19" />
                    <SPLIT distance="350" swimtime="00:04:15.63" />
                    <SPLIT distance="400" swimtime="00:04:55.08" />
                    <SPLIT distance="450" swimtime="00:05:34.52" />
                    <SPLIT distance="500" swimtime="00:06:13.44" />
                    <SPLIT distance="550" swimtime="00:06:53.18" />
                    <SPLIT distance="600" swimtime="00:07:32.04" />
                    <SPLIT distance="650" swimtime="00:08:10.83" />
                    <SPLIT distance="700" swimtime="00:08:49.43" />
                    <SPLIT distance="750" swimtime="00:09:28.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="494" reactiontime="+62" swimtime="00:04:38.35" resultid="17051" heatid="19011" lane="8" entrytime="00:04:37.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.73" />
                    <SPLIT distance="100" swimtime="00:01:05.51" />
                    <SPLIT distance="150" swimtime="00:01:40.78" />
                    <SPLIT distance="200" swimtime="00:02:16.11" />
                    <SPLIT distance="250" swimtime="00:02:51.68" />
                    <SPLIT distance="300" swimtime="00:03:27.63" />
                    <SPLIT distance="350" swimtime="00:04:03.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="399" reactiontime="+60" swimtime="00:02:30.36" resultid="17052" heatid="19059" lane="8" entrytime="00:02:28.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                    <SPLIT distance="100" swimtime="00:01:11.47" />
                    <SPLIT distance="150" swimtime="00:01:51.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="425" reactiontime="+68" swimtime="00:19:17.83" resultid="17053" heatid="19100" lane="7" entrytime="00:18:20.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                    <SPLIT distance="100" swimtime="00:01:09.68" />
                    <SPLIT distance="150" swimtime="00:01:47.05" />
                    <SPLIT distance="200" swimtime="00:02:24.83" />
                    <SPLIT distance="250" swimtime="00:03:02.89" />
                    <SPLIT distance="300" swimtime="00:03:41.63" />
                    <SPLIT distance="350" swimtime="00:04:20.15" />
                    <SPLIT distance="400" swimtime="00:04:59.06" />
                    <SPLIT distance="450" swimtime="00:05:37.89" />
                    <SPLIT distance="500" swimtime="00:06:16.87" />
                    <SPLIT distance="550" swimtime="00:06:56.32" />
                    <SPLIT distance="600" swimtime="00:07:35.86" />
                    <SPLIT distance="650" swimtime="00:08:15.27" />
                    <SPLIT distance="700" swimtime="00:08:54.47" />
                    <SPLIT distance="750" swimtime="00:09:33.59" />
                    <SPLIT distance="800" swimtime="00:10:12.51" />
                    <SPLIT distance="850" swimtime="00:10:51.41" />
                    <SPLIT distance="900" swimtime="00:11:30.47" />
                    <SPLIT distance="950" swimtime="00:12:09.18" />
                    <SPLIT distance="1000" swimtime="00:12:48.33" />
                    <SPLIT distance="1050" swimtime="00:13:27.75" />
                    <SPLIT distance="1100" swimtime="00:14:07.32" />
                    <SPLIT distance="1150" swimtime="00:14:46.34" />
                    <SPLIT distance="1200" swimtime="00:15:26.18" />
                    <SPLIT distance="1250" swimtime="00:16:05.48" />
                    <SPLIT distance="1300" swimtime="00:16:44.59" />
                    <SPLIT distance="1350" swimtime="00:17:23.37" />
                    <SPLIT distance="1400" swimtime="00:18:02.33" />
                    <SPLIT distance="1450" swimtime="00:18:40.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02203" nation="POL" region="03" clubid="17154" name="KS AZS AWF Biała Podlaska">
          <ATHLETES>
            <ATHLETE firstname="Piotr" lastname="Jędrzejczyk" birthdate="2007-03-20" gender="M" nation="POL" license="102203700117" swrid="5399698" athleteid="17194">
              <RESULTS>
                <RESULT eventid="1087" points="165" reactiontime="+95" swimtime="00:03:05.82" resultid="17195" heatid="18986" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.80" />
                    <SPLIT distance="100" swimtime="00:01:24.10" />
                    <SPLIT distance="150" swimtime="00:02:14.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="184" swimtime="00:00:36.71" resultid="17196" heatid="18952" lane="5" />
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej, a przed sygnałem startu" eventid="1113" reactiontime="+75" status="DSQ" swimtime="00:00:46.25" resultid="17197" heatid="19020" lane="7" />
                <RESULT eventid="1121" points="165" reactiontime="+91" swimtime="00:00:43.70" resultid="17198" heatid="19032" lane="4" />
                <RESULT eventid="1163" points="187" reactiontime="+82" swimtime="00:01:21.89" resultid="17199" heatid="19067" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.29" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej, a przed sygnałem startu" eventid="1171" reactiontime="+91" status="DSQ" swimtime="00:01:36.99" resultid="17200" heatid="19083" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kornelia" lastname="Siennicka" birthdate="2005-04-25" gender="F" nation="POL" license="102203600122" swrid="4552475" athleteid="17168">
              <RESULTS>
                <RESULT eventid="1108" points="209" reactiontime="+89" swimtime="00:00:41.11" resultid="17169" heatid="19013" lane="3" />
                <RESULT eventid="1159" points="286" reactiontime="+87" swimtime="00:01:18.48" resultid="17170" heatid="19061" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1059" points="325" swimtime="00:00:34.40" resultid="17171" heatid="18946" lane="2" />
                <RESULT eventid="1083" points="238" swimtime="00:03:02.24" resultid="17172" heatid="18982" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                    <SPLIT distance="100" swimtime="00:01:22.86" />
                    <SPLIT distance="150" swimtime="00:02:12.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="275" swimtime="00:00:41.46" resultid="17173" heatid="19026" lane="5" />
                <RESULT eventid="1167" points="245" reactiontime="+99" swimtime="00:01:31.97" resultid="17174" heatid="19079" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Dragan" birthdate="2008-01-04" gender="F" nation="POL" license="102203600108" swrid="5085637" athleteid="17155">
              <RESULTS>
                <RESULT eventid="1108" points="133" reactiontime="+88" swimtime="00:00:47.80" resultid="17156" heatid="19014" lane="8" />
                <RESULT eventid="1159" points="220" reactiontime="+82" swimtime="00:01:25.59" resultid="17157" heatid="19060" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1059" points="280" reactiontime="+88" swimtime="00:00:36.16" resultid="17158" heatid="18946" lane="8" />
                <RESULT eventid="1067" points="228" reactiontime="+89" swimtime="00:00:48.08" resultid="17159" heatid="18963" lane="5" />
                <RESULT eventid="1133" points="245" swimtime="00:01:42.38" resultid="17160" heatid="19039" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="244" swimtime="00:03:42.47" resultid="17161" heatid="19090" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.69" />
                    <SPLIT distance="100" swimtime="00:01:46.26" />
                    <SPLIT distance="150" swimtime="00:02:44.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Borsuk" birthdate="2002-05-04" gender="M" nation="POL" license="102203700033" swrid="4945690" athleteid="17207">
              <RESULTS>
                <RESULT eventid="1063" points="587" reactiontime="+67" swimtime="00:00:24.96" resultid="17208" heatid="18962" lane="2" entrytime="00:00:25.17" entrycourse="LCM" />
                <RESULT eventid="1079" points="429" reactiontime="+69" swimtime="00:01:05.59" resultid="17209" heatid="18980" lane="3" entrytime="00:01:05.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="558" reactiontime="+71" swimtime="00:00:27.05" resultid="17210" heatid="19025" lane="7" entrytime="00:00:26.89" entrycourse="LCM" />
                <RESULT eventid="1121" points="494" reactiontime="+67" swimtime="00:00:30.34" resultid="17211" heatid="19037" lane="2" entrytime="00:00:30.24" entrycourse="LCM" />
                <RESULT eventid="1163" points="592" reactiontime="+71" swimtime="00:00:55.86" resultid="17212" heatid="19077" lane="1" entrytime="00:00:55.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Makaruk" birthdate="2003-02-09" gender="M" nation="POL" license="102203700038" swrid="5033819" athleteid="17187">
              <RESULTS>
                <RESULT eventid="1087" points="462" reactiontime="+89" swimtime="00:02:11.87" resultid="17188" heatid="18986" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.23" />
                    <SPLIT distance="100" swimtime="00:01:02.96" />
                    <SPLIT distance="150" swimtime="00:01:37.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="504" reactiontime="+83" swimtime="00:00:26.26" resultid="17189" heatid="18962" lane="9" entrytime="00:00:26.36" entrycourse="LCM" />
                <RESULT eventid="1113" points="420" reactiontime="+86" swimtime="00:00:29.72" resultid="17190" heatid="19023" lane="5" entrytime="00:00:29.60" entrycourse="LCM" />
                <RESULT eventid="1121" points="518" reactiontime="+69" swimtime="00:00:29.87" resultid="17191" heatid="19037" lane="3" entrytime="00:00:30.09" entrycourse="LCM" />
                <RESULT eventid="1163" points="521" reactiontime="+92" swimtime="00:00:58.28" resultid="17192" heatid="19076" lane="1" entrytime="00:00:57.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="444" reactiontime="+75" swimtime="00:01:07.93" resultid="17193" heatid="19088" lane="7" entrytime="00:01:06.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Godlewski" birthdate="2009-01-25" gender="M" nation="POL" license="102203700110" swrid="5140959" athleteid="17201">
              <RESULTS>
                <RESULT eventid="1063" points="286" reactiontime="+73" swimtime="00:00:31.73" resultid="17202" heatid="18953" lane="6" />
                <RESULT eventid="1071" points="242" reactiontime="+84" swimtime="00:00:41.61" resultid="17203" heatid="18969" lane="7" />
                <RESULT eventid="1113" points="162" reactiontime="+61" swimtime="00:00:40.81" resultid="17204" heatid="19020" lane="2" />
                <RESULT eventid="1137" points="249" reactiontime="+86" swimtime="00:01:30.37" resultid="17205" heatid="19042" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="264" reactiontime="+78" swimtime="00:01:13.04" resultid="17206" heatid="19072" lane="0" entrytime="00:01:12.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maksymilian" lastname="Mich" birthdate="2006-06-28" gender="M" nation="POL" license="102203700060" swrid="5033812" athleteid="17182">
              <RESULTS>
                <RESULT eventid="1087" points="445" reactiontime="+69" swimtime="00:02:13.51" resultid="17183" heatid="18990" lane="2" entrytime="00:02:15.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                    <SPLIT distance="100" swimtime="00:01:02.63" />
                    <SPLIT distance="150" swimtime="00:01:38.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="520" reactiontime="+79" swimtime="00:00:26.00" resultid="17184" heatid="18961" lane="4" entrytime="00:00:26.38" entrycourse="LCM" />
                <RESULT eventid="1113" points="439" reactiontime="+82" swimtime="00:00:29.29" resultid="17185" heatid="19024" lane="9" entrytime="00:00:29.50" entrycourse="LCM" />
                <RESULT eventid="1163" points="516" reactiontime="+83" swimtime="00:00:58.46" resultid="17186" heatid="19075" lane="5" entrytime="00:00:58.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Zieliński" birthdate="2009-04-16" gender="M" nation="POL" license="102203700116" swrid="5399667" athleteid="17175">
              <RESULTS>
                <RESULT eventid="1087" points="172" reactiontime="+89" swimtime="00:03:03.06" resultid="17176" heatid="18987" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.74" />
                    <SPLIT distance="100" swimtime="00:01:25.56" />
                    <SPLIT distance="150" swimtime="00:02:15.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="239" reactiontime="+81" swimtime="00:00:33.66" resultid="17177" heatid="18952" lane="7" />
                <RESULT eventid="1137" points="208" reactiontime="+75" swimtime="00:01:35.87" resultid="17178" heatid="19043" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="231" reactiontime="+86" swimtime="00:00:39.08" resultid="17179" heatid="19033" lane="1" />
                <RESULT eventid="1163" points="218" reactiontime="+95" swimtime="00:01:17.87" resultid="17180" heatid="19070" lane="6" entrytime="00:01:17.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="208" reactiontime="+84" swimtime="00:01:27.42" resultid="17181" heatid="19085" lane="4" entrytime="00:01:27.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwia" lastname="Silipicka" birthdate="2002-10-24" gender="F" nation="POL" license="102203600034" swrid="4900055" athleteid="17162">
              <RESULTS>
                <RESULT eventid="1108" points="415" reactiontime="+70" swimtime="00:00:32.73" resultid="17163" heatid="19016" lane="3" entrytime="00:00:32.38" entrycourse="LCM" />
                <RESULT eventid="1159" points="433" reactiontime="+66" swimtime="00:01:08.30" resultid="17164" heatid="19064" lane="8" entrytime="00:01:07.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1059" points="477" reactiontime="+68" swimtime="00:00:30.29" resultid="17165" heatid="18950" lane="7" entrytime="00:00:29.88" entrycourse="LCM" />
                <RESULT eventid="1075" points="373" reactiontime="+83" swimtime="00:01:17.04" resultid="17166" heatid="18976" lane="0" entrytime="00:01:17.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="448" reactiontime="+85" swimtime="00:00:35.26" resultid="17167" heatid="19028" lane="3" entrytime="00:00:36.24" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01103" nation="POL" region="03" clubid="17582" name="MTP ,,Lublinianka&apos;&apos;">
          <ATHLETES>
            <ATHLETE firstname="Jakub" lastname="Kulbieda" birthdate="2005-10-07" gender="M" nation="POL" license="101103700170" swrid="5087791" athleteid="17649">
              <RESULTS>
                <RESULT eventid="1063" points="332" reactiontime="+67" swimtime="00:00:30.18" resultid="17650" heatid="18959" lane="3" entrytime="00:00:30.22" entrycourse="LCM" />
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej, a przed sygnałem startu" eventid="1071" reactiontime="+47" status="DSQ" swimtime="00:00:41.63" resultid="17651" heatid="18972" lane="1" entrytime="00:00:41.21" entrycourse="LCM" />
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej, a przed sygnałem startu" eventid="1121" reactiontime="+44" status="DSQ" swimtime="00:00:33.99" resultid="17652" heatid="19036" lane="7" entrytime="00:00:33.71" entrycourse="LCM" />
                <RESULT eventid="1171" points="322" reactiontime="+75" swimtime="00:01:15.62" resultid="17654" heatid="19087" lane="9" entrytime="00:01:14.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emilia" lastname="Adamek" birthdate="2008-08-27" gender="F" nation="POL" license="101103600182" swrid="5105309" athleteid="17728">
              <RESULTS>
                <RESULT eventid="1075" points="274" reactiontime="+73" swimtime="00:01:25.40" resultid="17729" heatid="18975" lane="3" entrytime="00:01:25.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" status="DNS" swimtime="00:00:00.00" resultid="17730" heatid="18998" lane="6" />
                <RESULT eventid="1125" points="396" reactiontime="+71" swimtime="00:05:21.89" resultid="17731" heatid="19005" lane="3" entrytime="00:05:26.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.21" />
                    <SPLIT distance="100" swimtime="00:01:16.38" />
                    <SPLIT distance="150" swimtime="00:01:57.26" />
                    <SPLIT distance="200" swimtime="00:02:37.96" />
                    <SPLIT distance="250" swimtime="00:03:19.36" />
                    <SPLIT distance="300" swimtime="00:04:00.81" />
                    <SPLIT distance="350" swimtime="00:04:42.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="330" reactiontime="+72" swimtime="00:03:02.50" resultid="17732" heatid="19049" lane="7" entrytime="00:03:03.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.57" />
                    <SPLIT distance="100" swimtime="00:01:26.42" />
                    <SPLIT distance="150" swimtime="00:02:22.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="316" reactiontime="+81" swimtime="00:01:24.45" resultid="17733" heatid="19080" lane="3" entrytime="00:01:21.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="385" swimtime="00:11:06.17" resultid="17734" heatid="19096" lane="6" entrytime="00:11:12.16" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Krukowski" birthdate="2008-11-18" gender="M" nation="POL" license="101103700231" swrid="5431080" athleteid="17659">
              <RESULTS>
                <RESULT eventid="1063" points="230" reactiontime="+64" swimtime="00:00:34.09" resultid="17660" heatid="18956" lane="6" entrytime="00:00:35.59" entrycourse="LCM" />
                <RESULT eventid="1087" points="186" reactiontime="+79" swimtime="00:02:58.59" resultid="17661" heatid="18988" lane="1" entrytime="00:03:00.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.57" />
                    <SPLIT distance="100" swimtime="00:01:23.15" />
                    <SPLIT distance="150" swimtime="00:02:13.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="149" reactiontime="+84" swimtime="00:00:42.00" resultid="17662" heatid="19018" lane="3" />
                <RESULT eventid="1121" points="164" reactiontime="+68" swimtime="00:00:43.81" resultid="17663" heatid="19032" lane="0" />
                <RESULT eventid="1163" points="211" reactiontime="+80" swimtime="00:01:18.71" resultid="17664" heatid="19068" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="141" reactiontime="+73" swimtime="00:01:39.48" resultid="17665" heatid="19083" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Kiełbasa" birthdate="2008-04-16" gender="M" nation="POL" license="101103700247" athleteid="17758">
              <RESULTS>
                <RESULT eventid="1121" points="85" reactiontime="+73" swimtime="00:00:54.40" resultid="17759" heatid="19031" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Zielińska" birthdate="2007-07-19" gender="F" nation="POL" license="101103600172" swrid="4879723" athleteid="17701">
              <RESULTS>
                <RESULT eventid="1067" points="527" reactiontime="+58" swimtime="00:00:36.39" resultid="17702" heatid="18967" lane="9" entrytime="00:00:36.30" entrycourse="LCM" />
                <RESULT eventid="1099" points="419" reactiontime="+74" swimtime="00:05:55.82" resultid="17703" heatid="18999" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                    <SPLIT distance="100" swimtime="00:01:17.46" />
                    <SPLIT distance="150" swimtime="00:02:06.12" />
                    <SPLIT distance="200" swimtime="00:02:53.68" />
                    <SPLIT distance="250" swimtime="00:03:41.03" />
                    <SPLIT distance="300" swimtime="00:04:29.63" />
                    <SPLIT distance="350" swimtime="00:05:13.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="422" reactiontime="+73" swimtime="00:05:15.12" resultid="17704" heatid="19006" lane="1" entrytime="00:05:11.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                    <SPLIT distance="100" swimtime="00:01:13.44" />
                    <SPLIT distance="150" swimtime="00:01:53.85" />
                    <SPLIT distance="200" swimtime="00:02:34.42" />
                    <SPLIT distance="250" swimtime="00:03:14.56" />
                    <SPLIT distance="300" swimtime="00:03:54.62" />
                    <SPLIT distance="350" swimtime="00:04:34.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="509" reactiontime="+72" swimtime="00:01:20.28" resultid="17705" heatid="19041" lane="6" entrytime="00:01:18.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="439" reactiontime="+72" swimtime="00:01:08.03" resultid="17706" heatid="19060" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="514" reactiontime="+80" swimtime="00:02:53.65" resultid="17707" heatid="19091" lane="6" entrytime="00:02:49.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                    <SPLIT distance="100" swimtime="00:01:24.97" />
                    <SPLIT distance="150" swimtime="00:02:10.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zofia" lastname="Wożakowska" birthdate="2007-11-20" gender="F" nation="POL" license="101103600171" swrid="5006494" athleteid="17694">
              <RESULTS>
                <RESULT eventid="1067" points="453" reactiontime="+70" swimtime="00:00:38.27" resultid="17695" heatid="18966" lane="3" entrytime="00:00:38.46" entrycourse="LCM" />
                <RESULT eventid="1083" points="466" swimtime="00:02:25.69" resultid="17696" heatid="18984" lane="8" entrytime="00:02:25.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                    <SPLIT distance="100" swimtime="00:01:09.82" />
                    <SPLIT distance="150" swimtime="00:01:47.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" status="DNS" swimtime="00:00:00.00" resultid="17697" heatid="19006" lane="8" entrytime="00:05:11.80" entrycourse="LCM" />
                <RESULT eventid="1133" status="DNS" swimtime="00:00:00.00" resultid="17698" heatid="19040" lane="5" entrytime="00:01:23.12" entrycourse="LCM" />
                <RESULT eventid="1175" status="DNS" swimtime="00:00:00.00" resultid="17699" heatid="19091" lane="0" entrytime="00:02:57.76" entrycourse="LCM" />
                <RESULT eventid="1183" status="DNS" swimtime="00:00:00.00" resultid="17700" heatid="19096" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonina" lastname="Jadach" birthdate="2007-09-02" gender="F" nation="POL" license="101103600213" swrid="5331782" athleteid="17595">
              <RESULTS>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej, a przed sygnałem startu" eventid="1059" reactiontime="+47" status="DSQ" swimtime="00:00:36.26" resultid="17596" heatid="18947" lane="4" entrytime="00:00:36.60" entrycourse="LCM" />
                <RESULT eventid="1067" points="191" reactiontime="+65" swimtime="00:00:51.03" resultid="17597" heatid="18965" lane="9" entrytime="00:00:52.12" entrycourse="LCM" />
                <RESULT eventid="1133" status="DNS" swimtime="00:00:00.00" resultid="17598" heatid="19039" lane="2" />
                <RESULT eventid="1159" points="254" reactiontime="+78" swimtime="00:01:21.63" resultid="17599" heatid="19062" lane="7" entrytime="00:01:21.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Mitrus" birthdate="2006-04-01" gender="F" nation="POL" license="101103600157" swrid="5019836" athleteid="17586">
              <RESULTS>
                <RESULT eventid="1059" points="446" reactiontime="+66" swimtime="00:00:30.98" resultid="17587" heatid="18949" lane="6" entrytime="00:00:31.01" entrycourse="LCM" />
                <RESULT eventid="1067" points="379" reactiontime="+70" swimtime="00:00:40.62" resultid="17588" heatid="18966" lane="7" entrytime="00:00:39.68" entrycourse="LCM" />
                <RESULT eventid="1108" points="365" reactiontime="+66" swimtime="00:00:34.18" resultid="17589" heatid="19016" lane="1" entrytime="00:00:33.05" entrycourse="LCM" />
                <RESULT comment="K11 - Pływak wykonał nierównoczesne lub naprzemienne ruchy nóg" eventid="1133" reactiontime="+66" status="DSQ" swimtime="00:00:00.00" resultid="17590" heatid="19040" lane="6" entrytime="00:01:27.14" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sebastian" lastname="Sak" birthdate="2008-11-14" gender="M" nation="POL" license="101103700196" swrid="4135746" athleteid="17647">
              <RESULTS>
                <RESULT eventid="1063" points="129" swimtime="00:00:41.37" resultid="17648" heatid="18955" lane="9" entrytime="00:00:40.48" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zofia" lastname="Górna" birthdate="2009-12-10" gender="F" nation="POL" license="101103600218" swrid="5286978" athleteid="17742">
              <RESULTS>
                <RESULT eventid="1091" points="276" reactiontime="+80" swimtime="00:03:09.23" resultid="17743" heatid="18993" lane="8" entrytime="00:03:06.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.31" />
                    <SPLIT distance="100" swimtime="00:01:32.08" />
                    <SPLIT distance="150" swimtime="00:02:22.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="185" swimtime="00:00:42.84" resultid="17744" heatid="19014" lane="0" />
                <RESULT eventid="1117" points="335" reactiontime="+76" swimtime="00:00:38.83" resultid="17745" heatid="19028" lane="2" entrytime="00:00:37.81" entrycourse="LCM" />
                <RESULT eventid="1167" points="340" reactiontime="+65" swimtime="00:01:22.42" resultid="17746" heatid="19080" lane="7" entrytime="00:01:25.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Krusiński" birthdate="2008-02-22" gender="M" nation="POL" license="101103700197" swrid="4133263" athleteid="17655">
              <RESULTS>
                <RESULT eventid="1063" points="159" reactiontime="+70" swimtime="00:00:38.59" resultid="17656" heatid="18955" lane="5" entrytime="00:00:38.47" entrycourse="LCM" />
                <RESULT eventid="1121" status="DNS" swimtime="00:00:00.00" resultid="17657" heatid="19034" lane="5" entrytime="00:00:43.93" entrycourse="LCM" />
                <RESULT eventid="1163" status="DNS" swimtime="00:00:00.00" resultid="17658" heatid="19067" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Bożek" birthdate="2005-07-24" gender="M" nation="POL" license="101103700242" swrid="4917582" athleteid="17619">
              <RESULTS>
                <RESULT eventid="1063" points="415" reactiontime="+81" swimtime="00:00:28.03" resultid="17620" heatid="18960" lane="4" entrytime="00:00:27.83" entrycourse="LCM" />
                <RESULT eventid="1121" points="417" reactiontime="+57" swimtime="00:00:32.10" resultid="17621" heatid="19037" lane="0" entrytime="00:00:32.17" entrycourse="LCM" />
                <RESULT eventid="1171" points="371" reactiontime="+57" swimtime="00:01:12.14" resultid="17623" heatid="19087" lane="5" entrytime="00:01:11.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Sawczuk" birthdate="2009-06-24" gender="F" nation="POL" license="101103600250" athleteid="18617">
              <RESULTS>
                <RESULT eventid="1117" status="DNS" swimtime="00:00:00.00" resultid="18618" heatid="19026" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hanna" lastname="Fus" birthdate="2009-08-11" gender="F" nation="POL" license="101103600207" swrid="4135757" athleteid="17606">
              <RESULTS>
                <RESULT eventid="1059" points="361" reactiontime="+71" swimtime="00:00:33.23" resultid="17607" heatid="18948" lane="3" entrytime="00:00:32.94" entrycourse="LCM" />
                <RESULT eventid="1067" points="298" reactiontime="+72" swimtime="00:00:43.99" resultid="17608" heatid="18965" lane="4" entrytime="00:00:44.01" entrycourse="LCM" />
                <RESULT eventid="1125" points="235" reactiontime="+76" swimtime="00:06:22.70" resultid="17609" heatid="19005" lane="7" entrytime="00:06:14.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                    <SPLIT distance="100" swimtime="00:01:29.65" />
                    <SPLIT distance="150" swimtime="00:02:19.42" />
                    <SPLIT distance="200" swimtime="00:03:10.11" />
                    <SPLIT distance="250" swimtime="00:04:00.11" />
                    <SPLIT distance="300" swimtime="00:04:50.48" />
                    <SPLIT distance="350" swimtime="00:05:41.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="256" reactiontime="+73" swimtime="00:01:40.99" resultid="17610" heatid="19039" lane="4" entrytime="00:01:43.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="310" reactiontime="+59" swimtime="00:01:16.34" resultid="17611" heatid="19063" lane="8" entrytime="00:01:12.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cezary" lastname="Rudawski" birthdate="2009-08-07" gender="M" nation="POL" license="101103700206" swrid="4622966" athleteid="17747">
              <RESULTS>
                <RESULT eventid="1095" points="319" reactiontime="+75" swimtime="00:02:43.64" resultid="17748" heatid="18996" lane="4" entrytime="00:02:43.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                    <SPLIT distance="100" swimtime="00:01:19.27" />
                    <SPLIT distance="150" swimtime="00:02:02.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6365" points="288" reactiontime="+76" swimtime="00:11:24.08" resultid="17749" heatid="19002" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.15" />
                    <SPLIT distance="100" swimtime="00:01:21.46" />
                    <SPLIT distance="150" swimtime="00:02:05.94" />
                    <SPLIT distance="200" swimtime="00:02:50.52" />
                    <SPLIT distance="250" swimtime="00:03:34.43" />
                    <SPLIT distance="300" swimtime="00:04:18.48" />
                    <SPLIT distance="350" swimtime="00:05:00.69" />
                    <SPLIT distance="400" swimtime="00:05:43.16" />
                    <SPLIT distance="450" swimtime="00:06:25.68" />
                    <SPLIT distance="500" swimtime="00:07:08.67" />
                    <SPLIT distance="550" swimtime="00:07:51.37" />
                    <SPLIT distance="600" swimtime="00:08:34.62" />
                    <SPLIT distance="650" swimtime="00:09:17.59" />
                    <SPLIT distance="700" swimtime="00:10:01.56" />
                    <SPLIT distance="750" swimtime="00:10:44.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="347" reactiontime="+65" swimtime="00:00:34.14" resultid="17750" heatid="19036" lane="0" entrytime="00:00:34.35" entrycourse="LCM" />
                <RESULT eventid="1145" points="282" reactiontime="+70" swimtime="00:02:53.79" resultid="17751" heatid="19053" lane="2" entrytime="00:02:51.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.03" />
                    <SPLIT distance="100" swimtime="00:01:23.03" />
                    <SPLIT distance="150" swimtime="00:02:14.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="328" reactiontime="+66" swimtime="00:01:15.16" resultid="17752" heatid="19086" lane="4" entrytime="00:01:15.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="308" reactiontime="+74" swimtime="00:03:06.61" resultid="17753" heatid="19092" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.56" />
                    <SPLIT distance="100" swimtime="00:01:28.90" />
                    <SPLIT distance="150" swimtime="00:02:19.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Pogoda" birthdate="2006-05-22" gender="F" nation="POL" license="101103600274" swrid="5461056" athleteid="17592">
              <RESULTS>
                <RESULT eventid="1059" points="281" reactiontime="+67" swimtime="00:00:36.13" resultid="17593" heatid="18948" lane="0" entrytime="00:00:35.84" entrycourse="LCM" />
                <RESULT eventid="1159" points="256" reactiontime="+75" swimtime="00:01:21.37" resultid="17594" heatid="19060" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksander" lastname="Stępniak" birthdate="2006-12-16" gender="M" nation="POL" license="101103700188" swrid="4133531" athleteid="17680">
              <RESULTS>
                <RESULT eventid="1063" points="348" reactiontime="+70" swimtime="00:00:29.70" resultid="17681" heatid="18959" lane="4" entrytime="00:00:29.96" entrycourse="LCM" />
                <RESULT eventid="1087" points="334" reactiontime="+73" swimtime="00:02:26.94" resultid="17682" heatid="18989" lane="4" entrytime="00:02:27.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.53" />
                    <SPLIT distance="100" swimtime="00:01:08.01" />
                    <SPLIT distance="150" swimtime="00:01:48.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="323" reactiontime="+53" swimtime="00:00:32.43" resultid="17683" heatid="19022" lane="2" entrytime="00:00:32.77" entrycourse="LCM" />
                <RESULT eventid="1145" points="299" reactiontime="+78" swimtime="00:02:50.35" resultid="17684" heatid="19053" lane="7" entrytime="00:02:52.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                    <SPLIT distance="100" swimtime="00:01:18.71" />
                    <SPLIT distance="150" swimtime="00:02:11.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="352" reactiontime="+76" swimtime="00:01:06.43" resultid="17685" heatid="19073" lane="1" entrytime="00:01:06.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="242" reactiontime="+84" swimtime="00:01:23.17" resultid="17686" heatid="19086" lane="0" entrytime="00:01:22.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Furmańczuk" birthdate="2009-02-04" gender="M" nation="POL" license="101103700257" athleteid="17762">
              <RESULTS>
                <RESULT eventid="1121" points="97" reactiontime="+87" swimtime="00:00:52.23" resultid="17763" heatid="19032" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrian" lastname="Dziewulski" birthdate="2006-08-22" gender="M" nation="POL" license="101103700158" swrid="5019837" athleteid="17629">
              <RESULTS>
                <RESULT eventid="1063" points="313" reactiontime="+66" swimtime="00:00:30.77" resultid="17630" heatid="18959" lane="0" entrytime="00:00:31.14" entrycourse="LCM" />
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej, a przed sygnałem startu" eventid="1071" status="DSQ" swimtime="00:00:39.39" resultid="17631" heatid="18972" lane="3" entrytime="00:00:40.15" entrycourse="LCM" />
                <RESULT eventid="1137" points="280" reactiontime="+77" swimtime="00:01:26.93" resultid="17632" heatid="19043" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksander" lastname="Dąbek" birthdate="2008-08-11" gender="M" nation="POL" license="101103700193" swrid="5173023" athleteid="17721">
              <RESULTS>
                <RESULT eventid="1071" points="265" swimtime="00:00:40.37" resultid="17722" heatid="18972" lane="2" entrytime="00:00:40.80" entrycourse="LCM" />
                <RESULT eventid="1103" points="274" reactiontime="+63" swimtime="00:06:15.37" resultid="17723" heatid="19000" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.25" />
                    <SPLIT distance="100" swimtime="00:01:31.45" />
                    <SPLIT distance="150" swimtime="00:02:20.00" />
                    <SPLIT distance="200" swimtime="00:03:06.34" />
                    <SPLIT distance="250" swimtime="00:03:58.39" />
                    <SPLIT distance="300" swimtime="00:04:49.70" />
                    <SPLIT distance="350" swimtime="00:05:33.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="259" reactiontime="+47" swimtime="00:00:34.92" resultid="17724" heatid="19022" lane="1" entrytime="00:00:35.86" entrycourse="LCM" />
                <RESULT eventid="1137" points="255" reactiontime="+47" swimtime="00:01:29.61" resultid="17725" heatid="19042" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="232" reactiontime="+66" swimtime="00:01:24.35" resultid="17726" heatid="19086" lane="1" entrytime="00:01:21.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="292" reactiontime="+64" swimtime="00:03:10.01" resultid="17727" heatid="19093" lane="2" entrytime="00:03:19.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.85" />
                    <SPLIT distance="100" swimtime="00:01:33.49" />
                    <SPLIT distance="150" swimtime="00:02:22.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kinga" lastname="Gąsior" birthdate="2008-10-02" gender="F" nation="POL" license="101103600183" swrid="5109078" athleteid="17687">
              <RESULTS>
                <RESULT eventid="1067" points="350" reactiontime="+46" swimtime="00:00:41.68" resultid="17688" heatid="18966" lane="2" entrytime="00:00:39.56" entrycourse="LCM" />
                <RESULT eventid="1091" points="330" reactiontime="+68" swimtime="00:02:58.41" resultid="17689" heatid="18993" lane="2" entrytime="00:02:52.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.82" />
                    <SPLIT distance="100" swimtime="00:01:27.55" />
                    <SPLIT distance="150" swimtime="00:02:13.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="351" reactiontime="+68" swimtime="00:00:38.22" resultid="17690" heatid="19028" lane="6" entrytime="00:00:37.07" entrycourse="LCM" />
                <RESULT eventid="1133" points="327" reactiontime="+68" swimtime="00:01:33.08" resultid="17691" heatid="19040" lane="2" entrytime="00:01:29.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" status="DNS" swimtime="00:00:00.00" resultid="17692" heatid="19080" lane="5" entrytime="00:01:21.50" entrycourse="LCM" />
                <RESULT eventid="1175" points="346" reactiontime="+51" swimtime="00:03:18.12" resultid="17693" heatid="19090" lane="5" entrytime="00:03:11.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.95" />
                    <SPLIT distance="100" swimtime="00:01:36.06" />
                    <SPLIT distance="150" swimtime="00:02:29.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Weronika" lastname="Baranowska" birthdate="2009-04-28" gender="F" nation="POL" license="101103600219" swrid="5288415" athleteid="17715">
              <RESULTS>
                <RESULT eventid="1067" points="289" reactiontime="+73" swimtime="00:00:44.43" resultid="17716" heatid="18964" lane="1" />
                <RESULT eventid="1083" points="284" reactiontime="+87" swimtime="00:02:51.79" resultid="17717" heatid="18982" lane="4" entrytime="00:02:53.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                    <SPLIT distance="100" swimtime="00:01:24.69" />
                    <SPLIT distance="150" swimtime="00:02:11.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="287" swimtime="00:00:37.01" resultid="17718" heatid="19015" lane="2" entrytime="00:00:37.89" entrycourse="LCM" />
                <RESULT eventid="1141" points="284" reactiontime="+76" swimtime="00:03:11.67" resultid="17719" heatid="19049" lane="1" entrytime="00:03:05.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.58" />
                    <SPLIT distance="100" swimtime="00:01:32.61" />
                    <SPLIT distance="150" swimtime="00:02:30.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="292" reactiontime="+68" swimtime="00:12:09.97" resultid="17720" heatid="19095" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.20" />
                    <SPLIT distance="100" swimtime="00:01:24.47" />
                    <SPLIT distance="150" swimtime="00:02:12.29" />
                    <SPLIT distance="200" swimtime="00:02:59.27" />
                    <SPLIT distance="250" swimtime="00:03:46.27" />
                    <SPLIT distance="300" swimtime="00:04:32.94" />
                    <SPLIT distance="350" swimtime="00:05:20.93" />
                    <SPLIT distance="400" swimtime="00:06:07.55" />
                    <SPLIT distance="450" swimtime="00:06:55.08" />
                    <SPLIT distance="500" swimtime="00:07:42.83" />
                    <SPLIT distance="550" swimtime="00:08:28.94" />
                    <SPLIT distance="600" swimtime="00:09:15.22" />
                    <SPLIT distance="650" swimtime="00:10:00.26" />
                    <SPLIT distance="700" swimtime="00:10:45.61" />
                    <SPLIT distance="750" swimtime="00:11:29.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Wołoszko" birthdate="2008-12-30" gender="M" nation="POL" license="101103700194" swrid="5225183" athleteid="17666">
              <RESULTS>
                <RESULT eventid="1063" points="221" reactiontime="+79" swimtime="00:00:34.58" resultid="17667" heatid="18957" lane="6" entrytime="00:00:33.61" entrycourse="LCM" />
                <RESULT eventid="1087" points="204" reactiontime="+79" swimtime="00:02:53.26" resultid="17668" heatid="18988" lane="3" entrytime="00:02:52.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.10" />
                    <SPLIT distance="100" swimtime="00:01:24.29" />
                    <SPLIT distance="150" swimtime="00:02:09.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="234" reactiontime="+76" swimtime="00:05:57.06" resultid="17669" heatid="19010" lane="9" entrytime="00:06:41.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.84" />
                    <SPLIT distance="100" swimtime="00:01:22.56" />
                    <SPLIT distance="150" swimtime="00:02:08.93" />
                    <SPLIT distance="200" swimtime="00:02:57.12" />
                    <SPLIT distance="250" swimtime="00:03:43.71" />
                    <SPLIT distance="300" swimtime="00:04:32.66" />
                    <SPLIT distance="350" swimtime="00:05:18.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="132" reactiontime="+90" swimtime="00:00:47.09" resultid="17670" heatid="19034" lane="4" entrytime="00:00:43.54" entrycourse="LCM" />
                <RESULT eventid="1163" points="233" reactiontime="+89" swimtime="00:01:16.21" resultid="17671" heatid="19071" lane="8" entrytime="00:01:16.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="117" reactiontime="+99" swimtime="00:01:45.75" resultid="17672" heatid="19084" lane="5" entrytime="00:01:50.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Kamola" birthdate="2008-08-22" gender="M" nation="POL" license="101103700195" swrid="4135743" athleteid="17673">
              <RESULTS>
                <RESULT eventid="1113" points="226" reactiontime="+72" swimtime="00:00:36.51" resultid="17676" heatid="19021" lane="4" entrytime="00:00:37.00" entrycourse="LCM" />
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej, a przed sygnałem startu" eventid="1137" reactiontime="+56" status="DSQ" swimtime="00:01:37.84" resultid="17677" heatid="19045" lane="6" entrytime="00:01:34.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="256" reactiontime="+60" swimtime="00:01:13.87" resultid="17678" heatid="19071" lane="5" entrytime="00:01:14.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="199" reactiontime="+72" swimtime="00:01:28.69" resultid="17679" heatid="19084" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Michałek" birthdate="2006-02-13" gender="M" nation="POL" license="101103700169" swrid="4917589" athleteid="17735">
              <RESULTS>
                <RESULT eventid="1079" points="414" reactiontime="+73" swimtime="00:01:06.37" resultid="17736" heatid="18980" lane="5" entrytime="00:01:04.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="411" reactiontime="+78" swimtime="00:05:27.92" resultid="17737" heatid="19000" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                    <SPLIT distance="100" swimtime="00:01:11.39" />
                    <SPLIT distance="150" swimtime="00:01:53.15" />
                    <SPLIT distance="200" swimtime="00:02:34.29" />
                    <SPLIT distance="250" swimtime="00:03:24.78" />
                    <SPLIT distance="300" swimtime="00:04:14.81" />
                    <SPLIT distance="350" swimtime="00:04:52.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="511" reactiontime="+72" swimtime="00:00:27.84" resultid="17738" heatid="19024" lane="6" entrytime="00:00:27.92" entrycourse="LCM" />
                <RESULT eventid="1145" points="425" reactiontime="+77" swimtime="00:02:31.54" resultid="17739" heatid="19054" lane="0" entrytime="00:02:27.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.58" />
                    <SPLIT distance="100" swimtime="00:01:09.24" />
                    <SPLIT distance="150" swimtime="00:01:57.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="498" reactiontime="+72" swimtime="00:00:59.15" resultid="17740" heatid="19076" lane="9" entrytime="00:00:58.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" status="DNS" swimtime="00:00:00.00" resultid="17741" heatid="19100" lane="8" entrytime="00:18:29.06" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kalina" lastname="Jakubiak" birthdate="2009-04-23" gender="F" nation="POL" license="101103600214" swrid="5339634" athleteid="17708">
              <RESULTS>
                <RESULT eventid="1067" points="321" reactiontime="+67" swimtime="00:00:42.92" resultid="17709" heatid="18964" lane="2" />
                <RESULT eventid="1099" points="348" reactiontime="+82" swimtime="00:06:18.51" resultid="17710" heatid="18998" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.25" />
                    <SPLIT distance="100" swimtime="00:01:24.88" />
                    <SPLIT distance="150" swimtime="00:02:15.58" />
                    <SPLIT distance="200" swimtime="00:03:02.82" />
                    <SPLIT distance="250" swimtime="00:03:55.51" />
                    <SPLIT distance="300" swimtime="00:04:49.46" />
                    <SPLIT distance="350" swimtime="00:05:35.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="392" reactiontime="+88" swimtime="00:00:36.86" resultid="17711" heatid="19026" lane="3" />
                <RESULT eventid="1141" points="339" reactiontime="+97" swimtime="00:03:00.87" resultid="17712" heatid="19049" lane="2" entrytime="00:03:00.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.11" />
                    <SPLIT distance="100" swimtime="00:01:24.95" />
                    <SPLIT distance="150" swimtime="00:02:18.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="338" reactiontime="+88" swimtime="00:01:22.58" resultid="17713" heatid="19080" lane="6" entrytime="00:01:23.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="315" swimtime="00:03:24.35" resultid="17714" heatid="19090" lane="2" entrytime="00:03:20.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.10" />
                    <SPLIT distance="100" swimtime="00:01:40.39" />
                    <SPLIT distance="150" swimtime="00:02:34.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Weronika" lastname="Drozd" birthdate="2005-11-16" gender="F" nation="POL" license="101103600243" swrid="5455430" athleteid="17583">
              <RESULTS>
                <RESULT eventid="1059" points="276" reactiontime="+68" swimtime="00:00:36.35" resultid="17584" heatid="18947" lane="8" entrytime="00:00:38.38" entrycourse="LCM" />
                <RESULT eventid="1117" points="178" reactiontime="+70" swimtime="00:00:47.96" resultid="17585" heatid="19027" lane="8" entrytime="00:00:47.36" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martyna" lastname="Mazurek" birthdate="2009-08-11" gender="F" nation="POL" license="101103600209" swrid="5287010" athleteid="17612">
              <RESULTS>
                <RESULT eventid="1059" points="235" swimtime="00:00:38.35" resultid="17613" heatid="18947" lane="2" entrytime="00:00:37.48" entrycourse="LCM" />
                <RESULT eventid="1067" points="169" reactiontime="+69" swimtime="00:00:53.17" resultid="17614" heatid="18964" lane="4" entrytime="00:00:52.89" entrycourse="LCM" />
                <RESULT eventid="1108" points="122" reactiontime="+59" swimtime="00:00:49.15" resultid="17615" heatid="19014" lane="4" entrytime="00:00:46.76" entrycourse="LCM" />
                <RESULT eventid="1141" points="201" swimtime="00:03:35.30" resultid="17616" heatid="19048" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.28" />
                    <SPLIT distance="100" swimtime="00:01:43.50" />
                    <SPLIT distance="150" swimtime="00:02:46.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="197" swimtime="00:01:28.82" resultid="17617" heatid="19062" lane="8" entrytime="00:01:25.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="203" reactiontime="+92" swimtime="00:01:37.85" resultid="17618" heatid="19079" lane="5" entrytime="00:01:37.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Czech" birthdate="2003-03-14" gender="M" nation="POL" license="101103700228" swrid="5431067" athleteid="17624">
              <RESULTS>
                <RESULT eventid="1063" points="235" reactiontime="+76" swimtime="00:00:33.84" resultid="17625" heatid="18956" lane="4" entrytime="00:00:34.54" entrycourse="LCM" />
                <RESULT eventid="1071" points="194" reactiontime="+82" swimtime="00:00:44.75" resultid="17626" heatid="18971" lane="5" entrytime="00:00:42.95" entrycourse="LCM" />
                <RESULT eventid="1137" status="DNS" swimtime="00:00:00.00" resultid="17627" heatid="19045" lane="8" entrytime="00:01:36.72" entrycourse="LCM" />
                <RESULT eventid="1163" status="DNS" swimtime="00:00:00.00" resultid="17628" heatid="19070" lane="1" entrytime="00:01:17.56" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Konrad" lastname="Gordziejko" birthdate="2006-10-28" gender="M" nation="POL" license="101103700198" swrid="5043779" athleteid="17633">
              <RESULTS>
                <RESULT eventid="1063" points="422" reactiontime="+61" swimtime="00:00:27.86" resultid="17634" heatid="18959" lane="5" entrytime="00:00:30.21" entrycourse="LCM" />
                <RESULT eventid="6365" points="438" reactiontime="+70" swimtime="00:09:55.05" resultid="17635" heatid="19003" lane="0" entrytime="00:09:39.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                    <SPLIT distance="100" swimtime="00:01:07.46" />
                    <SPLIT distance="150" swimtime="00:01:44.57" />
                    <SPLIT distance="200" swimtime="00:02:21.06" />
                    <SPLIT distance="250" swimtime="00:02:57.82" />
                    <SPLIT distance="300" swimtime="00:03:35.79" />
                    <SPLIT distance="350" swimtime="00:04:12.65" />
                    <SPLIT distance="400" swimtime="00:04:50.89" />
                    <SPLIT distance="450" swimtime="00:05:28.48" />
                    <SPLIT distance="500" swimtime="00:06:07.47" />
                    <SPLIT distance="550" swimtime="00:06:46.62" />
                    <SPLIT distance="600" swimtime="00:07:24.03" />
                    <SPLIT distance="650" swimtime="00:08:02.66" />
                    <SPLIT distance="700" swimtime="00:08:41.49" />
                    <SPLIT distance="750" swimtime="00:09:18.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="453" reactiontime="+69" swimtime="00:04:46.34" resultid="17636" heatid="19011" lane="0" entrytime="00:04:38.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                    <SPLIT distance="100" swimtime="00:01:07.02" />
                    <SPLIT distance="150" swimtime="00:01:43.15" />
                    <SPLIT distance="200" swimtime="00:02:20.53" />
                    <SPLIT distance="250" swimtime="00:02:56.76" />
                    <SPLIT distance="300" swimtime="00:03:34.61" />
                    <SPLIT distance="350" swimtime="00:04:11.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="398" reactiontime="+76" swimtime="00:00:32.61" resultid="17637" heatid="19036" lane="4" entrytime="00:00:33.02" entrycourse="LCM" />
                <RESULT eventid="1163" points="478" reactiontime="+45" swimtime="00:00:59.98" resultid="17638" heatid="19075" lane="8" entrytime="00:00:59.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" status="DNS" swimtime="00:00:00.00" resultid="17639" heatid="19087" lane="3" entrytime="00:01:11.81" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antoni" lastname="Bajek" birthdate="2009-08-25" gender="M" nation="POL" license="101103700256" athleteid="17754">
              <RESULTS>
                <RESULT eventid="1121" status="DNS" swimtime="00:00:00.00" resultid="17755" heatid="19032" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alicja" lastname="Piasecka" birthdate="2008-02-04" gender="F" nation="POL" license="101103600201" swrid="4880035" athleteid="17600">
              <RESULTS>
                <RESULT eventid="1059" points="344" reactiontime="+70" swimtime="00:00:33.78" resultid="17601" heatid="18948" lane="6" entrytime="00:00:33.41" entrycourse="LCM" />
                <RESULT eventid="1083" points="305" reactiontime="+58" swimtime="00:02:47.75" resultid="17602" heatid="18982" lane="5" entrytime="00:02:55.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                    <SPLIT distance="100" swimtime="00:01:22.56" />
                    <SPLIT distance="150" swimtime="00:02:07.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="276" reactiontime="+71" swimtime="00:00:41.42" resultid="17603" heatid="19028" lane="1" entrytime="00:00:39.88" entrycourse="LCM" />
                <RESULT eventid="1159" points="330" reactiontime="+73" swimtime="00:01:14.76" resultid="17604" heatid="19062" lane="6" entrytime="00:01:19.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="224" reactiontime="+76" swimtime="00:01:34.76" resultid="17605" heatid="19080" lane="9" entrytime="00:01:33.60" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Pietrow" birthdate="2009-06-30" gender="M" nation="POL" license="101103700255" athleteid="17760">
              <RESULTS>
                <RESULT eventid="1121" status="DNS" swimtime="00:00:00.00" resultid="17761" heatid="19031" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Gordziejko" birthdate="2010-07-14" gender="F" nation="POL" license="101103600236" athleteid="19102">
              <RESULTS>
                <RESULT eventid="1059" points="272" reactiontime="+73" status="EXH" swimtime="00:00:36.51" resultid="19103" heatid="18945" lane="8" />
                <RESULT eventid="1067" status="DNS" swimtime="00:00:00.00" resultid="19104" heatid="18963" lane="6" />
                <RESULT eventid="1133" status="DNS" swimtime="00:00:00.00" resultid="19105" heatid="19038" lane="6" />
                <RESULT eventid="1159" status="DNS" swimtime="00:00:00.00" resultid="19106" heatid="19060" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maksym" lastname="Kapuśniak" birthdate="2006-12-19" gender="M" nation="POL" license="101103700168" swrid="4879704" athleteid="17640">
              <RESULTS>
                <RESULT eventid="1063" points="539" reactiontime="+62" swimtime="00:00:25.69" resultid="17641" heatid="18962" lane="1" entrytime="00:00:25.64" entrycourse="LCM" />
                <RESULT eventid="1071" points="520" reactiontime="+71" swimtime="00:00:32.27" resultid="17642" heatid="18974" lane="7" entrytime="00:00:31.92" entrycourse="LCM" />
                <RESULT eventid="1137" points="484" reactiontime="+69" swimtime="00:01:12.44" resultid="17643" heatid="19047" lane="6" entrytime="00:01:10.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="425" reactiontime="+76" swimtime="00:02:31.52" resultid="17644" heatid="19054" lane="9" entrytime="00:02:31.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                    <SPLIT distance="100" swimtime="00:01:12.69" />
                    <SPLIT distance="150" swimtime="00:01:57.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="554" reactiontime="+71" swimtime="00:00:57.10" resultid="17645" heatid="19076" lane="7" entrytime="00:00:57.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="462" reactiontime="+73" swimtime="00:02:43.06" resultid="17646" heatid="19094" lane="6" entrytime="00:02:42.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.54" />
                    <SPLIT distance="100" swimtime="00:01:20.14" />
                    <SPLIT distance="150" swimtime="00:02:04.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="08314" nation="POL" region="14" clubid="18446" name="UKS Delfin Garwolin">
          <ATHLETES>
            <ATHLETE firstname="Alicja" lastname="Więckowska" birthdate="2003-02-10" gender="F" nation="POL" license="108314600059" swrid="5056729" athleteid="18453">
              <RESULTS>
                <RESULT eventid="1125" points="531" reactiontime="+80" status="EXH" swimtime="00:04:51.98" resultid="18454" heatid="19006" lane="7" entrytime="00:04:58.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                    <SPLIT distance="100" swimtime="00:01:08.29" />
                    <SPLIT distance="150" swimtime="00:01:45.35" />
                    <SPLIT distance="200" swimtime="00:02:22.78" />
                    <SPLIT distance="250" swimtime="00:03:00.69" />
                    <SPLIT distance="300" swimtime="00:03:38.32" />
                    <SPLIT distance="350" swimtime="00:04:16.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6361" points="525" status="EXH" swimtime="00:19:00.38" resultid="18455" heatid="19055" lane="5" entrytime="00:19:13.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                    <SPLIT distance="100" swimtime="00:01:10.11" />
                    <SPLIT distance="150" swimtime="00:01:47.53" />
                    <SPLIT distance="200" swimtime="00:02:24.81" />
                    <SPLIT distance="250" swimtime="00:03:02.57" />
                    <SPLIT distance="300" swimtime="00:03:40.19" />
                    <SPLIT distance="350" swimtime="00:04:18.17" />
                    <SPLIT distance="400" swimtime="00:04:56.03" />
                    <SPLIT distance="450" swimtime="00:05:34.09" />
                    <SPLIT distance="500" swimtime="00:06:12.33" />
                    <SPLIT distance="550" swimtime="00:06:50.64" />
                    <SPLIT distance="600" swimtime="00:07:28.99" />
                    <SPLIT distance="650" swimtime="00:08:07.39" />
                    <SPLIT distance="700" swimtime="00:08:45.42" />
                    <SPLIT distance="750" swimtime="00:09:23.56" />
                    <SPLIT distance="800" swimtime="00:10:01.94" />
                    <SPLIT distance="850" swimtime="00:10:40.57" />
                    <SPLIT distance="900" swimtime="00:11:18.89" />
                    <SPLIT distance="950" swimtime="00:11:57.72" />
                    <SPLIT distance="1000" swimtime="00:12:36.24" />
                    <SPLIT distance="1050" swimtime="00:13:15.12" />
                    <SPLIT distance="1100" swimtime="00:13:54.17" />
                    <SPLIT distance="1150" swimtime="00:14:33.10" />
                    <SPLIT distance="1200" swimtime="00:15:12.15" />
                    <SPLIT distance="1250" swimtime="00:15:50.96" />
                    <SPLIT distance="1300" swimtime="00:16:29.42" />
                    <SPLIT distance="1350" swimtime="00:17:08.19" />
                    <SPLIT distance="1400" swimtime="00:17:46.86" />
                    <SPLIT distance="1450" swimtime="00:18:25.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="537" status="EXH" swimtime="00:09:56.40" resultid="18456" heatid="19097" lane="8" entrytime="00:10:09.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.14" />
                    <SPLIT distance="100" swimtime="00:01:09.94" />
                    <SPLIT distance="150" swimtime="00:01:47.58" />
                    <SPLIT distance="200" swimtime="00:02:25.11" />
                    <SPLIT distance="250" swimtime="00:03:02.65" />
                    <SPLIT distance="300" swimtime="00:03:40.55" />
                    <SPLIT distance="350" swimtime="00:04:18.37" />
                    <SPLIT distance="400" swimtime="00:04:56.12" />
                    <SPLIT distance="450" swimtime="00:05:33.93" />
                    <SPLIT distance="500" swimtime="00:06:11.95" />
                    <SPLIT distance="550" swimtime="00:06:49.82" />
                    <SPLIT distance="600" swimtime="00:07:27.65" />
                    <SPLIT distance="650" swimtime="00:08:05.60" />
                    <SPLIT distance="700" swimtime="00:08:43.49" />
                    <SPLIT distance="750" swimtime="00:09:20.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Sitnik" birthdate="2003-10-07" gender="M" nation="POL" license="108314700020" swrid="5120231" athleteid="18447">
              <RESULTS>
                <RESULT eventid="1063" points="500" reactiontime="+70" status="EXH" swimtime="00:00:26.33" resultid="18448" heatid="18962" lane="8" entrytime="00:00:25.73" entrycourse="LCM" />
                <RESULT eventid="1079" points="434" reactiontime="+79" status="EXH" swimtime="00:01:05.36" resultid="18449" heatid="18978" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="524" reactiontime="+68" status="EXH" swimtime="00:00:27.62" resultid="18450" heatid="19024" lane="4" entrytime="00:00:27.55" entrycourse="LCM" />
                <RESULT eventid="1145" points="415" reactiontime="+74" status="EXH" swimtime="00:02:32.73" resultid="18451" heatid="19053" lane="3" entrytime="00:02:39.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.23" />
                    <SPLIT distance="100" swimtime="00:01:11.57" />
                    <SPLIT distance="150" swimtime="00:01:58.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="483" reactiontime="+68" status="EXH" swimtime="00:00:59.76" resultid="18452" heatid="19075" lane="2" entrytime="00:00:59.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04503" nation="POL" region="03" clubid="16864" name="Bialski Klub Zimowego Pływania Arua-Aqua">
          <ATHLETES>
            <ATHLETE firstname="Ewelina" lastname="Cuch" birthdate="1979-02-05" gender="F" nation="POL" license="504593600001" athleteid="16865">
              <RESULTS>
                <RESULT eventid="1067" points="291" reactiontime="+85" status="EXH" swimtime="00:00:44.35" resultid="16866" heatid="18964" lane="8" />
                <RESULT eventid="1083" points="260" reactiontime="+85" status="EXH" swimtime="00:02:56.90" resultid="16867" heatid="18982" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                    <SPLIT distance="100" swimtime="00:01:20.26" />
                    <SPLIT distance="150" swimtime="00:02:06.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="273" reactiontime="+86" status="EXH" swimtime="00:00:37.62" resultid="16868" heatid="19014" lane="6" />
                <RESULT eventid="1133" points="265" reactiontime="+69" status="EXH" swimtime="00:01:39.78" resultid="16869" heatid="19039" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="267" reactiontime="+92" status="EXH" swimtime="00:01:20.21" resultid="16870" heatid="19060" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="240" reactiontime="+88" status="EXH" swimtime="00:03:43.57" resultid="16871" heatid="19089" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.66" />
                    <SPLIT distance="100" swimtime="00:01:47.00" />
                    <SPLIT distance="150" swimtime="00:02:46.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00908" nation="POL" region="08" clubid="17913" name="SP Motyl MOSiR Stalowa Wola">
          <ATHLETES>
            <ATHLETE firstname="Adam" lastname="Procnal" birthdate="2004-08-03" gender="M" nation="POL" license="100908700307" swrid="5020343" athleteid="17914">
              <RESULTS>
                <RESULT eventid="1079" points="543" reactiontime="+68" status="EXH" swimtime="00:01:00.65" resultid="17915" heatid="18981" lane="2" entrytime="00:01:00.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="535" reactiontime="+68" status="EXH" swimtime="00:05:00.35" resultid="17916" heatid="19001" lane="3" entrytime="00:05:03.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.08" />
                    <SPLIT distance="100" swimtime="00:01:04.66" />
                    <SPLIT distance="150" swimtime="00:01:44.57" />
                    <SPLIT distance="200" swimtime="00:02:24.48" />
                    <SPLIT distance="250" swimtime="00:03:07.57" />
                    <SPLIT distance="300" swimtime="00:03:51.34" />
                    <SPLIT distance="350" swimtime="00:04:26.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="567" reactiontime="+71" status="EXH" swimtime="00:04:25.78" resultid="17917" heatid="19011" lane="4" entrytime="00:04:26.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.40" />
                    <SPLIT distance="100" swimtime="00:01:02.52" />
                    <SPLIT distance="150" swimtime="00:01:36.41" />
                    <SPLIT distance="200" swimtime="00:02:10.31" />
                    <SPLIT distance="250" swimtime="00:02:44.68" />
                    <SPLIT distance="300" swimtime="00:03:19.30" />
                    <SPLIT distance="350" swimtime="00:03:53.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="540" reactiontime="+69" status="EXH" swimtime="00:02:19.93" resultid="17918" heatid="19054" lane="1" entrytime="00:02:20.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.07" />
                    <SPLIT distance="100" swimtime="00:01:07.04" />
                    <SPLIT distance="150" swimtime="00:01:47.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="512" reactiontime="+74" status="EXH" swimtime="00:02:18.41" resultid="17919" heatid="19059" lane="6" entrytime="00:02:16.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.38" />
                    <SPLIT distance="100" swimtime="00:01:05.92" />
                    <SPLIT distance="150" swimtime="00:01:42.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="467" reactiontime="+65" status="EXH" swimtime="00:01:06.83" resultid="17920" heatid="19088" lane="1" entrytime="00:01:07.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="09514" nation="POL" region="14" clubid="17963" name="UKP ,,Polonia Warszawa&apos;&apos;">
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Guliński" birthdate="2004-08-19" gender="M" nation="POL" license="109514700258" swrid="5034149" athleteid="17972">
              <RESULTS>
                <RESULT eventid="1155" points="624" reactiontime="+72" status="EXH" swimtime="00:02:09.52" resultid="17973" heatid="19059" lane="5" entrytime="00:02:12.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.29" />
                    <SPLIT distance="100" swimtime="00:01:01.03" />
                    <SPLIT distance="150" swimtime="00:01:35.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Bolek" birthdate="2005-07-02" gender="M" nation="POL" license="109514700030" swrid="5004416" athleteid="17968">
              <RESULTS>
                <RESULT eventid="1095" points="526" reactiontime="+58" status="EXH" swimtime="00:02:18.57" resultid="17969" heatid="18997" lane="2" entrytime="00:02:24.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.06" />
                    <SPLIT distance="100" swimtime="00:01:07.04" />
                    <SPLIT distance="150" swimtime="00:01:43.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="631" reactiontime="+71" status="EXH" swimtime="00:04:16.50" resultid="17970" heatid="19012" lane="2" entrytime="00:04:14.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.71" />
                    <SPLIT distance="100" swimtime="00:01:00.02" />
                    <SPLIT distance="150" swimtime="00:01:32.58" />
                    <SPLIT distance="200" swimtime="00:02:05.24" />
                    <SPLIT distance="250" swimtime="00:02:37.92" />
                    <SPLIT distance="300" swimtime="00:03:10.82" />
                    <SPLIT distance="350" swimtime="00:03:44.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="659" reactiontime="+74" status="EXH" swimtime="00:16:40.82" resultid="17971" heatid="19100" lane="3" entrytime="00:16:52.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.57" />
                    <SPLIT distance="100" swimtime="00:01:02.32" />
                    <SPLIT distance="150" swimtime="00:01:35.34" />
                    <SPLIT distance="200" swimtime="00:02:08.36" />
                    <SPLIT distance="250" swimtime="00:02:41.80" />
                    <SPLIT distance="300" swimtime="00:03:15.43" />
                    <SPLIT distance="350" swimtime="00:03:48.73" />
                    <SPLIT distance="400" swimtime="00:04:22.37" />
                    <SPLIT distance="450" swimtime="00:04:55.71" />
                    <SPLIT distance="500" swimtime="00:05:28.94" />
                    <SPLIT distance="550" swimtime="00:06:02.41" />
                    <SPLIT distance="600" swimtime="00:06:35.72" />
                    <SPLIT distance="650" swimtime="00:07:09.58" />
                    <SPLIT distance="700" swimtime="00:07:43.45" />
                    <SPLIT distance="750" swimtime="00:08:17.10" />
                    <SPLIT distance="800" swimtime="00:08:50.71" />
                    <SPLIT distance="850" swimtime="00:09:24.34" />
                    <SPLIT distance="900" swimtime="00:09:57.79" />
                    <SPLIT distance="950" swimtime="00:10:31.29" />
                    <SPLIT distance="1000" swimtime="00:11:05.15" />
                    <SPLIT distance="1050" swimtime="00:11:38.89" />
                    <SPLIT distance="1100" swimtime="00:12:13.03" />
                    <SPLIT distance="1150" swimtime="00:12:46.47" />
                    <SPLIT distance="1200" swimtime="00:13:20.11" />
                    <SPLIT distance="1250" swimtime="00:13:53.76" />
                    <SPLIT distance="1300" swimtime="00:14:27.84" />
                    <SPLIT distance="1350" swimtime="00:15:01.74" />
                    <SPLIT distance="1400" swimtime="00:15:35.46" />
                    <SPLIT distance="1450" swimtime="00:16:08.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matylda" lastname="Romaniuk" birthdate="2004-05-08" gender="F" nation="POL" license="109514600253" swrid="5083139" athleteid="17964">
              <RESULTS>
                <RESULT eventid="1091" points="538" reactiontime="+75" status="EXH" swimtime="00:02:31.60" resultid="17965" heatid="18992" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                    <SPLIT distance="100" swimtime="00:01:13.64" />
                    <SPLIT distance="150" swimtime="00:01:53.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="575" reactiontime="+73" status="EXH" swimtime="00:04:44.29" resultid="17966" heatid="19006" lane="4" entrytime="00:04:46.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.26" />
                    <SPLIT distance="100" swimtime="00:01:08.26" />
                    <SPLIT distance="150" swimtime="00:01:44.94" />
                    <SPLIT distance="200" swimtime="00:02:21.32" />
                    <SPLIT distance="250" swimtime="00:02:57.49" />
                    <SPLIT distance="300" swimtime="00:03:33.75" />
                    <SPLIT distance="350" swimtime="00:04:09.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="524" reactiontime="+70" status="EXH" swimtime="00:01:11.39" resultid="17967" heatid="19079" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01803" nation="POL" region="03" clubid="18364" name="UKS ,,Wodnik Krasnystaw&apos;&apos;">
          <ATHLETES>
            <ATHLETE firstname="Fabian" lastname="Wiśniewski" birthdate="2009-08-30" gender="M" nation="POL" license="101803700038" swrid="4996311" athleteid="18371">
              <RESULTS>
                <RESULT eventid="1071" points="175" swimtime="00:00:46.38" resultid="18372" heatid="18971" lane="9" entrytime="00:00:45.11" entrycourse="LCM" />
                <RESULT eventid="1095" points="197" reactiontime="+57" swimtime="00:03:12.05" resultid="18373" heatid="18995" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.86" />
                    <SPLIT distance="100" swimtime="00:01:35.82" />
                    <SPLIT distance="150" swimtime="00:02:25.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="106" swimtime="00:00:46.99" resultid="18374" heatid="19019" lane="0" />
                <RESULT eventid="1137" points="183" swimtime="00:01:40.06" resultid="18375" heatid="19045" lane="0" entrytime="00:01:37.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="214" swimtime="00:03:30.62" resultid="18376" heatid="19093" lane="0" entrytime="00:03:26.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.18" />
                    <SPLIT distance="100" swimtime="00:01:43.70" />
                    <SPLIT distance="150" swimtime="00:02:38.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martyna" lastname="Lewandowska" birthdate="2007-04-15" gender="F" nation="POL" license="101803600035" swrid="4620536" athleteid="18365">
              <RESULTS>
                <RESULT eventid="1059" points="389" swimtime="00:00:32.42" resultid="18366" heatid="18949" lane="0" entrytime="00:00:31.56" entrycourse="LCM" />
                <RESULT eventid="1083" points="363" reactiontime="+88" swimtime="00:02:38.30" resultid="18367" heatid="18983" lane="7" entrytime="00:02:33.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                    <SPLIT distance="100" swimtime="00:01:16.82" />
                    <SPLIT distance="150" swimtime="00:01:58.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="331" reactiontime="+85" swimtime="00:00:35.30" resultid="18368" heatid="19015" lane="3" entrytime="00:00:35.48" entrycourse="LCM" />
                <RESULT eventid="1117" points="319" reactiontime="+68" swimtime="00:00:39.47" resultid="18369" heatid="19026" lane="6" />
                <RESULT eventid="1159" points="383" reactiontime="+87" swimtime="00:01:11.15" resultid="18370" heatid="19063" lane="3" entrytime="00:01:09.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Stawska" birthdate="2005-04-09" gender="F" nation="POL" license="101803600023" swrid="4837460" athleteid="17907">
              <RESULTS>
                <RESULT eventid="1091" points="586" reactiontime="+79" swimtime="00:02:27.34" resultid="17908" heatid="18994" lane="2" entrytime="00:02:29.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                    <SPLIT distance="100" swimtime="00:01:12.71" />
                    <SPLIT distance="150" swimtime="00:01:51.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="555" reactiontime="+79" swimtime="00:00:32.82" resultid="17909" heatid="19029" lane="4" entrytime="00:00:32.86" entrycourse="LCM" />
                <RESULT eventid="1141" points="517" reactiontime="+69" swimtime="00:02:37.13" resultid="17910" heatid="19050" lane="0" entrytime="00:02:33.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                    <SPLIT distance="100" swimtime="00:01:12.84" />
                    <SPLIT distance="150" swimtime="00:02:00.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="554" reactiontime="+76" swimtime="00:01:10.06" resultid="17911" heatid="19082" lane="8" entrytime="00:01:09.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="519" reactiontime="+80" swimtime="00:10:02.93" resultid="17912" heatid="19097" lane="1" entrytime="00:10:05.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                    <SPLIT distance="100" swimtime="00:01:11.85" />
                    <SPLIT distance="150" swimtime="00:01:49.95" />
                    <SPLIT distance="200" swimtime="00:02:28.12" />
                    <SPLIT distance="250" swimtime="00:03:06.15" />
                    <SPLIT distance="300" swimtime="00:03:44.56" />
                    <SPLIT distance="350" swimtime="00:04:22.82" />
                    <SPLIT distance="400" swimtime="00:05:01.23" />
                    <SPLIT distance="450" swimtime="00:05:39.25" />
                    <SPLIT distance="500" swimtime="00:06:17.75" />
                    <SPLIT distance="550" swimtime="00:06:56.15" />
                    <SPLIT distance="600" swimtime="00:07:34.48" />
                    <SPLIT distance="650" swimtime="00:08:12.68" />
                    <SPLIT distance="700" swimtime="00:08:50.59" />
                    <SPLIT distance="750" swimtime="00:09:27.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00103" nation="POL" region="03" clubid="18049" name="UKP Fala Kraśnik">
          <ATHLETES>
            <ATHLETE firstname="Dawid" lastname="Dzięgielewski" birthdate="2007-05-16" gender="M" nation="POL" license="100103700168" swrid="5148639" athleteid="18068">
              <RESULTS>
                <RESULT eventid="1071" points="402" reactiontime="+81" swimtime="00:00:35.15" resultid="18069" heatid="18973" lane="4" entrytime="00:00:35.22" entrycourse="LCM" />
                <RESULT eventid="1103" points="385" reactiontime="+87" swimtime="00:05:35.03" resultid="18070" heatid="19001" lane="7" entrytime="00:05:35.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                    <SPLIT distance="100" swimtime="00:01:15.47" />
                    <SPLIT distance="150" swimtime="00:02:00.86" />
                    <SPLIT distance="200" swimtime="00:02:44.79" />
                    <SPLIT distance="250" swimtime="00:03:30.42" />
                    <SPLIT distance="300" swimtime="00:04:15.69" />
                    <SPLIT distance="350" swimtime="00:04:56.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="303" reactiontime="+84" swimtime="00:00:33.15" resultid="18071" heatid="19020" lane="9" />
                <RESULT eventid="1137" points="385" reactiontime="+87" swimtime="00:01:18.18" resultid="18072" heatid="19047" lane="9" entrytime="00:01:17.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="380" reactiontime="+87" swimtime="00:02:54.05" resultid="18073" heatid="19094" lane="1" entrytime="00:02:49.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.61" />
                    <SPLIT distance="100" swimtime="00:01:22.48" />
                    <SPLIT distance="150" swimtime="00:02:08.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Wójcik" birthdate="2006-10-09" gender="M" nation="POL" license="100103700159" swrid="5164072" athleteid="18080">
              <RESULTS>
                <RESULT eventid="1079" points="488" reactiontime="+69" swimtime="00:01:02.84" resultid="18081" heatid="18980" lane="4" entrytime="00:01:03.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6365" points="548" reactiontime="+69" swimtime="00:09:12.26" resultid="18082" heatid="19003" lane="1" entrytime="00:09:16.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.04" />
                    <SPLIT distance="100" swimtime="00:01:02.86" />
                    <SPLIT distance="150" swimtime="00:01:36.60" />
                    <SPLIT distance="200" swimtime="00:02:10.89" />
                    <SPLIT distance="250" swimtime="00:02:45.36" />
                    <SPLIT distance="300" swimtime="00:03:19.90" />
                    <SPLIT distance="350" swimtime="00:03:54.85" />
                    <SPLIT distance="400" swimtime="00:04:30.37" />
                    <SPLIT distance="450" swimtime="00:05:05.85" />
                    <SPLIT distance="500" swimtime="00:05:40.99" />
                    <SPLIT distance="550" swimtime="00:06:16.19" />
                    <SPLIT distance="600" swimtime="00:06:51.10" />
                    <SPLIT distance="650" swimtime="00:07:26.81" />
                    <SPLIT distance="700" swimtime="00:08:02.05" />
                    <SPLIT distance="750" swimtime="00:08:37.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="547" reactiontime="+66" swimtime="00:04:29.03" resultid="18083" heatid="19011" lane="3" entrytime="00:04:28.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.82" />
                    <SPLIT distance="100" swimtime="00:01:03.18" />
                    <SPLIT distance="150" swimtime="00:01:37.21" />
                    <SPLIT distance="200" swimtime="00:02:11.81" />
                    <SPLIT distance="250" swimtime="00:02:46.84" />
                    <SPLIT distance="300" swimtime="00:03:21.60" />
                    <SPLIT distance="350" swimtime="00:03:55.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="489" reactiontime="+67" swimtime="00:00:28.25" resultid="18084" heatid="19024" lane="1" entrytime="00:00:28.42" entrycourse="LCM" />
                <RESULT eventid="1155" points="446" reactiontime="+74" swimtime="00:02:24.84" resultid="18085" heatid="19059" lane="1" entrytime="00:02:26.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                    <SPLIT distance="100" swimtime="00:01:08.59" />
                    <SPLIT distance="150" swimtime="00:01:46.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="557" reactiontime="+70" swimtime="00:17:38.03" resultid="18086" heatid="19100" lane="6" entrytime="00:17:34.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.49" />
                    <SPLIT distance="100" swimtime="00:01:03.99" />
                    <SPLIT distance="150" swimtime="00:01:38.71" />
                    <SPLIT distance="200" swimtime="00:02:13.39" />
                    <SPLIT distance="250" swimtime="00:02:48.22" />
                    <SPLIT distance="300" swimtime="00:03:23.42" />
                    <SPLIT distance="350" swimtime="00:03:58.94" />
                    <SPLIT distance="400" swimtime="00:04:34.57" />
                    <SPLIT distance="450" swimtime="00:05:09.99" />
                    <SPLIT distance="500" swimtime="00:05:45.30" />
                    <SPLIT distance="550" swimtime="00:06:20.49" />
                    <SPLIT distance="600" swimtime="00:06:55.92" />
                    <SPLIT distance="650" swimtime="00:07:31.61" />
                    <SPLIT distance="700" swimtime="00:08:07.31" />
                    <SPLIT distance="750" swimtime="00:08:43.15" />
                    <SPLIT distance="800" swimtime="00:09:18.75" />
                    <SPLIT distance="850" swimtime="00:09:54.55" />
                    <SPLIT distance="900" swimtime="00:10:30.48" />
                    <SPLIT distance="950" swimtime="00:11:06.42" />
                    <SPLIT distance="1000" swimtime="00:11:42.35" />
                    <SPLIT distance="1050" swimtime="00:12:18.48" />
                    <SPLIT distance="1100" swimtime="00:12:54.63" />
                    <SPLIT distance="1150" swimtime="00:13:30.82" />
                    <SPLIT distance="1200" swimtime="00:14:06.64" />
                    <SPLIT distance="1250" swimtime="00:14:42.79" />
                    <SPLIT distance="1300" swimtime="00:15:18.81" />
                    <SPLIT distance="1350" swimtime="00:15:54.78" />
                    <SPLIT distance="1400" swimtime="00:16:30.69" />
                    <SPLIT distance="1450" swimtime="00:17:05.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Surowiec" birthdate="2007-01-17" gender="F" nation="POL" license="100103600169" swrid="5148647" athleteid="18050">
              <RESULTS>
                <RESULT eventid="1059" points="453" reactiontime="+76" swimtime="00:00:30.80" resultid="18051" heatid="18945" lane="4" />
                <RESULT eventid="1091" points="510" reactiontime="+71" swimtime="00:02:34.32" resultid="18052" heatid="18994" lane="9" entrytime="00:02:33.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                    <SPLIT distance="100" swimtime="00:01:14.87" />
                    <SPLIT distance="150" swimtime="00:01:55.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="531" reactiontime="+68" swimtime="00:00:33.30" resultid="18053" heatid="19029" lane="5" entrytime="00:00:32.95" entrycourse="LCM" />
                <RESULT eventid="1133" points="455" reactiontime="+76" swimtime="00:01:23.36" resultid="18054" heatid="19038" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="500" reactiontime="+69" swimtime="00:01:12.52" resultid="18055" heatid="19081" lane="4" entrytime="00:01:10.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Sosnówka" birthdate="2007-08-20" gender="F" nation="POL" license="100103600167" swrid="5109105" athleteid="18074">
              <RESULTS>
                <RESULT eventid="1075" points="451" reactiontime="+80" swimtime="00:01:12.32" resultid="18075" heatid="18976" lane="4" entrytime="00:01:12.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="416" reactiontime="+80" swimtime="00:05:56.70" resultid="18076" heatid="18999" lane="1" entrytime="00:05:48.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.97" />
                    <SPLIT distance="100" swimtime="00:01:14.91" />
                    <SPLIT distance="150" swimtime="00:02:03.74" />
                    <SPLIT distance="200" swimtime="00:02:49.25" />
                    <SPLIT distance="250" swimtime="00:03:41.72" />
                    <SPLIT distance="300" swimtime="00:04:34.89" />
                    <SPLIT distance="350" swimtime="00:05:16.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="459" reactiontime="+78" swimtime="00:00:31.67" resultid="18077" heatid="19016" lane="5" entrytime="00:00:32.10" entrycourse="LCM" />
                <RESULT eventid="1150" points="371" reactiontime="+80" swimtime="00:02:49.44" resultid="18078" heatid="19057" lane="7" entrytime="00:02:46.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                    <SPLIT distance="100" swimtime="00:01:20.11" />
                    <SPLIT distance="150" swimtime="00:02:05.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="409" reactiontime="+80" swimtime="00:10:52.70" resultid="18079" heatid="19096" lane="3" entrytime="00:10:59.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                    <SPLIT distance="100" swimtime="00:01:15.54" />
                    <SPLIT distance="150" swimtime="00:01:57.22" />
                    <SPLIT distance="200" swimtime="00:02:38.60" />
                    <SPLIT distance="250" swimtime="00:03:19.06" />
                    <SPLIT distance="300" swimtime="00:04:00.52" />
                    <SPLIT distance="350" swimtime="00:04:41.24" />
                    <SPLIT distance="400" swimtime="00:05:22.89" />
                    <SPLIT distance="450" swimtime="00:06:03.74" />
                    <SPLIT distance="500" swimtime="00:06:44.49" />
                    <SPLIT distance="550" swimtime="00:07:27.57" />
                    <SPLIT distance="600" swimtime="00:08:10.49" />
                    <SPLIT distance="650" swimtime="00:08:52.92" />
                    <SPLIT distance="700" swimtime="00:09:35.16" />
                    <SPLIT distance="750" swimtime="00:10:14.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwia" lastname="Sosnówka" birthdate="2005-07-08" gender="F" nation="POL" license="100103600137" swrid="4971988" athleteid="18062">
              <RESULTS>
                <RESULT eventid="1067" points="365" reactiontime="+71" swimtime="00:00:41.12" resultid="18063" heatid="18963" lane="4" />
                <RESULT eventid="1075" points="412" reactiontime="+73" swimtime="00:01:14.50" resultid="18064" heatid="18976" lane="3" entrytime="00:01:13.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="378" reactiontime="+75" swimtime="00:00:33.77" resultid="18065" heatid="19014" lane="7" />
                <RESULT eventid="1133" points="405" reactiontime="+71" swimtime="00:01:26.62" resultid="18066" heatid="19038" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1150" points="433" reactiontime="+73" swimtime="00:02:40.94" resultid="18067" heatid="19057" lane="6" entrytime="00:02:36.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                    <SPLIT distance="100" swimtime="00:01:17.50" />
                    <SPLIT distance="150" swimtime="00:01:58.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Borsuk" birthdate="2003-12-19" gender="M" nation="POL" license="100103700122" swrid="4744848" athleteid="17893">
              <RESULTS>
                <RESULT eventid="1095" points="487" reactiontime="+69" swimtime="00:02:22.22" resultid="17894" heatid="18997" lane="3" entrytime="00:02:20.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                    <SPLIT distance="100" swimtime="00:01:08.51" />
                    <SPLIT distance="150" swimtime="00:01:45.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6365" points="526" reactiontime="+70" swimtime="00:09:19.76" resultid="17895" heatid="19003" lane="8" entrytime="00:09:20.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.64" />
                    <SPLIT distance="100" swimtime="00:01:03.86" />
                    <SPLIT distance="150" swimtime="00:01:38.34" />
                    <SPLIT distance="200" swimtime="00:02:13.84" />
                    <SPLIT distance="250" swimtime="00:02:48.85" />
                    <SPLIT distance="300" swimtime="00:03:24.01" />
                    <SPLIT distance="350" swimtime="00:03:58.82" />
                    <SPLIT distance="400" swimtime="00:04:34.26" />
                    <SPLIT distance="450" swimtime="00:05:09.65" />
                    <SPLIT distance="500" swimtime="00:05:46.74" />
                    <SPLIT distance="550" swimtime="00:06:22.67" />
                    <SPLIT distance="600" swimtime="00:06:58.67" />
                    <SPLIT distance="650" swimtime="00:07:35.14" />
                    <SPLIT distance="700" swimtime="00:08:10.89" />
                    <SPLIT distance="750" swimtime="00:08:45.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="395" reactiontime="+74" swimtime="00:04:59.85" resultid="17896" heatid="19011" lane="7" entrytime="00:04:31.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                    <SPLIT distance="100" swimtime="00:01:08.40" />
                    <SPLIT distance="150" swimtime="00:01:47.50" />
                    <SPLIT distance="200" swimtime="00:02:26.55" />
                    <SPLIT distance="250" swimtime="00:03:05.14" />
                    <SPLIT distance="300" swimtime="00:03:44.08" />
                    <SPLIT distance="350" swimtime="00:04:22.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="515" reactiontime="+71" swimtime="00:00:29.94" resultid="17897" heatid="19037" lane="5" entrytime="00:00:29.58" entrycourse="LCM" />
                <RESULT eventid="1171" points="509" reactiontime="+69" swimtime="00:01:04.93" resultid="17898" heatid="19088" lane="2" entrytime="00:01:05.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Błażej" lastname="Paszkowski" birthdate="2006-06-07" gender="M" nation="POL" license="100103700153" swrid="5108762" athleteid="17899">
              <RESULTS>
                <RESULT eventid="1095" points="640" reactiontime="+70" swimtime="00:02:09.87" resultid="17901" heatid="18997" lane="5" entrytime="00:02:11.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.67" />
                    <SPLIT distance="100" swimtime="00:01:03.65" />
                    <SPLIT distance="150" swimtime="00:01:37.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6365" points="598" reactiontime="+73" swimtime="00:08:56.36" resultid="17902" heatid="19003" lane="2" entrytime="00:09:07.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.13" />
                    <SPLIT distance="100" swimtime="00:01:02.95" />
                    <SPLIT distance="150" swimtime="00:01:36.47" />
                    <SPLIT distance="200" swimtime="00:02:10.40" />
                    <SPLIT distance="250" swimtime="00:02:44.57" />
                    <SPLIT distance="300" swimtime="00:03:18.10" />
                    <SPLIT distance="350" swimtime="00:03:50.89" />
                    <SPLIT distance="400" swimtime="00:04:24.86" />
                    <SPLIT distance="450" swimtime="00:04:58.29" />
                    <SPLIT distance="500" swimtime="00:05:32.37" />
                    <SPLIT distance="550" swimtime="00:06:06.33" />
                    <SPLIT distance="600" swimtime="00:06:40.85" />
                    <SPLIT distance="650" swimtime="00:07:14.67" />
                    <SPLIT distance="700" swimtime="00:07:48.81" />
                    <SPLIT distance="750" swimtime="00:08:22.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="551" reactiontime="+70" swimtime="00:00:27.15" resultid="17903" heatid="19025" lane="1" entrytime="00:00:26.96" entrycourse="LCM" />
                <RESULT eventid="1145" points="547" reactiontime="+73" swimtime="00:02:19.38" resultid="17905" heatid="19054" lane="7" entrytime="00:02:19.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.05" />
                    <SPLIT distance="100" swimtime="00:01:04.47" />
                    <SPLIT distance="150" swimtime="00:01:48.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="659" reactiontime="+68" swimtime="00:00:59.58" resultid="17906" heatid="19088" lane="5" entrytime="00:01:00.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Bucoń" birthdate="2007-01-31" gender="M" nation="POL" license="100103700155" swrid="4971980" athleteid="18087">
              <RESULTS>
                <RESULT eventid="1095" points="450" reactiontime="+69" swimtime="00:02:26.00" resultid="18088" heatid="18997" lane="6" entrytime="00:02:23.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                    <SPLIT distance="100" swimtime="00:01:10.40" />
                    <SPLIT distance="150" swimtime="00:01:48.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6365" points="450" reactiontime="+78" swimtime="00:09:49.67" resultid="18089" heatid="19002" lane="5" entrytime="00:09:50.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                    <SPLIT distance="100" swimtime="00:01:08.70" />
                    <SPLIT distance="150" swimtime="00:01:46.28" />
                    <SPLIT distance="200" swimtime="00:02:22.88" />
                    <SPLIT distance="250" swimtime="00:02:59.94" />
                    <SPLIT distance="300" swimtime="00:03:37.37" />
                    <SPLIT distance="350" swimtime="00:04:15.60" />
                    <SPLIT distance="400" swimtime="00:04:53.88" />
                    <SPLIT distance="450" swimtime="00:05:30.96" />
                    <SPLIT distance="500" swimtime="00:06:08.76" />
                    <SPLIT distance="550" swimtime="00:06:46.13" />
                    <SPLIT distance="600" swimtime="00:07:23.74" />
                    <SPLIT distance="650" swimtime="00:08:01.07" />
                    <SPLIT distance="700" swimtime="00:08:38.52" />
                    <SPLIT distance="750" swimtime="00:09:15.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1129" points="450" reactiontime="+69" swimtime="00:04:47.06" resultid="18090" heatid="19011" lane="9" entrytime="00:04:41.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.78" />
                    <SPLIT distance="100" swimtime="00:01:05.21" />
                    <SPLIT distance="150" swimtime="00:01:41.18" />
                    <SPLIT distance="200" swimtime="00:02:17.61" />
                    <SPLIT distance="250" swimtime="00:02:54.76" />
                    <SPLIT distance="300" swimtime="00:03:32.13" />
                    <SPLIT distance="350" swimtime="00:04:10.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="441" reactiontime="+68" swimtime="00:00:31.53" resultid="18091" heatid="19037" lane="1" entrytime="00:00:31.09" entrycourse="LCM" />
                <RESULT eventid="1163" points="402" reactiontime="+78" swimtime="00:01:03.53" resultid="18092" heatid="19074" lane="7" entrytime="00:01:02.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="457" reactiontime="+77" swimtime="00:18:50.65" resultid="18093" heatid="19100" lane="0" entrytime="00:18:30.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.52" />
                    <SPLIT distance="100" swimtime="00:01:10.75" />
                    <SPLIT distance="150" swimtime="00:01:48.38" />
                    <SPLIT distance="200" swimtime="00:02:26.32" />
                    <SPLIT distance="250" swimtime="00:03:04.21" />
                    <SPLIT distance="300" swimtime="00:03:42.05" />
                    <SPLIT distance="350" swimtime="00:04:20.03" />
                    <SPLIT distance="400" swimtime="00:04:58.26" />
                    <SPLIT distance="450" swimtime="00:05:36.71" />
                    <SPLIT distance="500" swimtime="00:06:14.67" />
                    <SPLIT distance="550" swimtime="00:06:52.95" />
                    <SPLIT distance="600" swimtime="00:07:31.05" />
                    <SPLIT distance="650" swimtime="00:08:09.52" />
                    <SPLIT distance="700" swimtime="00:08:47.89" />
                    <SPLIT distance="750" swimtime="00:09:26.42" />
                    <SPLIT distance="800" swimtime="00:10:05.04" />
                    <SPLIT distance="850" swimtime="00:10:42.24" />
                    <SPLIT distance="900" swimtime="00:11:20.11" />
                    <SPLIT distance="950" swimtime="00:11:58.51" />
                    <SPLIT distance="1000" swimtime="00:12:36.76" />
                    <SPLIT distance="1050" swimtime="00:13:15.44" />
                    <SPLIT distance="1100" swimtime="00:13:53.47" />
                    <SPLIT distance="1150" swimtime="00:14:31.09" />
                    <SPLIT distance="1200" swimtime="00:15:09.13" />
                    <SPLIT distance="1250" swimtime="00:15:46.78" />
                    <SPLIT distance="1300" swimtime="00:16:24.78" />
                    <SPLIT distance="1350" swimtime="00:17:02.30" />
                    <SPLIT distance="1400" swimtime="00:17:39.04" />
                    <SPLIT distance="1450" swimtime="00:18:15.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amelia" lastname="Wysocka" birthdate="2007-08-11" gender="F" nation="POL" license="100103600154" swrid="5109107" athleteid="18056">
              <RESULTS>
                <RESULT eventid="1059" points="676" reactiontime="+77" swimtime="00:00:26.96" resultid="18057" heatid="18951" lane="5" entrytime="00:00:26.91" entrycourse="LCM" />
                <RESULT eventid="1067" points="588" reactiontime="+58" swimtime="00:00:35.08" resultid="18058" heatid="18967" lane="2" entrytime="00:00:35.39" entrycourse="LCM" />
                <RESULT eventid="1108" points="601" reactiontime="+72" swimtime="00:00:28.94" resultid="18059" heatid="19017" lane="5" entrytime="00:00:28.65" entrycourse="LCM" />
                <RESULT eventid="1159" points="677" reactiontime="+73" swimtime="00:00:58.88" resultid="18060" heatid="19066" lane="6" entrytime="00:00:58.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="535" reactiontime="+76" swimtime="00:09:56.97" resultid="18061" heatid="19097" lane="2" entrytime="00:09:51.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                    <SPLIT distance="100" swimtime="00:01:08.47" />
                    <SPLIT distance="150" swimtime="00:01:46.48" />
                    <SPLIT distance="200" swimtime="00:02:23.85" />
                    <SPLIT distance="250" swimtime="00:03:01.84" />
                    <SPLIT distance="300" swimtime="00:03:39.85" />
                    <SPLIT distance="350" swimtime="00:04:18.37" />
                    <SPLIT distance="400" swimtime="00:04:56.11" />
                    <SPLIT distance="450" swimtime="00:05:34.02" />
                    <SPLIT distance="500" swimtime="00:06:12.09" />
                    <SPLIT distance="550" swimtime="00:06:50.49" />
                    <SPLIT distance="600" swimtime="00:07:28.36" />
                    <SPLIT distance="650" swimtime="00:08:05.65" />
                    <SPLIT distance="700" swimtime="00:08:43.90" />
                    <SPLIT distance="750" swimtime="00:09:21.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>

<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Warminsko-Mazurski Okregowy Zwiazek Plywacki" version="Build 29894">
    <CONTACT name="GeoLogix AG" street="Muristrasse 60" city="Bern" zip="3006" country="CH" phone="+41 31 356 80 56" fax="+41 31 356 80 81" email="info@splash-software.ch" internet="http://www.splash-software.ch" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Olsztyn" name="Letnie Mistrzostwa Polski w Pływaniu w kategorii Masters" name.en="Letnie Mistrzostwa Polski w Plywaniu Masters" course="LCM" deadline="2014-06-18" nation="POL" organizer="Masters Olsztyn" result.url="http://www.megatiming.pl" timing="AUTOMATIC">
      <AGEDATE value="2014-06-25" type="YEAR" />
      <POOL name="OSIR Aquasfera Olsztyn" lanemax="9" />
      <POINTTABLE pointtableid="3007" name="FINA Point Scoring" version="2014" />
      <CONTACT email="elachodyna@poczta.fm" name="Elżbieta Chodyna" phone="600215732" />
      <FEES>
        <FEE currency="PLN" type="ATHLETE" value="10000" />
        <FEE currency="PLN" type="LATEENTRY.INDIVIDUAL" value="15000" />
      </FEES>
      <SESSIONS>
        <SESSION date="2014-06-27" daytime="16:00" number="1" warmupfrom="14:45">
          <EVENTS>
            <EVENT eventid="98777" daytime="16:00" gender="F" number="1" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="98779" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103609" />
                    <RANKING order="2" place="2" resultid="102996" />
                    <RANKING order="3" place="3" resultid="102413" />
                    <RANKING order="4" place="4" resultid="100310" />
                    <RANKING order="5" place="-1" resultid="101719" />
                    <RANKING order="6" place="-1" resultid="103057" />
                    <RANKING order="7" place="-1" resultid="103469" />
                    <RANKING order="8" place="-1" resultid="103475" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98780" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103142" />
                    <RANKING order="2" place="2" resultid="101137" />
                    <RANKING order="3" place="3" resultid="102284" />
                    <RANKING order="4" place="4" resultid="103137" />
                    <RANKING order="5" place="5" resultid="102171" />
                    <RANKING order="6" place="6" resultid="103004" />
                    <RANKING order="7" place="7" resultid="101165" />
                    <RANKING order="8" place="8" resultid="103026" />
                    <RANKING order="9" place="9" resultid="101623" />
                    <RANKING order="10" place="10" resultid="101845" />
                    <RANKING order="11" place="11" resultid="102388" />
                    <RANKING order="12" place="12" resultid="100431" />
                    <RANKING order="13" place="-1" resultid="101224" />
                    <RANKING order="14" place="-1" resultid="101345" />
                    <RANKING order="15" place="-1" resultid="101616" />
                    <RANKING order="16" place="-1" resultid="102909" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98782" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102290" />
                    <RANKING order="2" place="2" resultid="103518" />
                    <RANKING order="3" place="3" resultid="101849" />
                    <RANKING order="4" place="4" resultid="100579" />
                    <RANKING order="5" place="-1" resultid="102954" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98783" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100178" />
                    <RANKING order="2" place="2" resultid="105049" />
                    <RANKING order="3" place="3" resultid="100172" />
                    <RANKING order="4" place="4" resultid="101685" />
                    <RANKING order="5" place="5" resultid="100879" />
                    <RANKING order="6" place="6" resultid="102796" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98781" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102053" />
                    <RANKING order="2" place="2" resultid="103330" />
                    <RANKING order="3" place="3" resultid="101798" />
                    <RANKING order="4" place="4" resultid="101356" />
                    <RANKING order="5" place="5" resultid="103130" />
                    <RANKING order="6" place="6" resultid="103124" />
                    <RANKING order="7" place="7" resultid="100232" />
                    <RANKING order="8" place="8" resultid="103342" />
                    <RANKING order="9" place="-1" resultid="100113" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98785" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103119" />
                    <RANKING order="2" place="2" resultid="103347" />
                    <RANKING order="3" place="3" resultid="100726" />
                    <RANKING order="4" place="4" resultid="105013" />
                    <RANKING order="5" place="5" resultid="103426" />
                    <RANKING order="6" place="6" resultid="100814" />
                    <RANKING order="7" place="7" resultid="101071" />
                    <RANKING order="8" place="8" resultid="105030" />
                    <RANKING order="9" place="9" resultid="100871" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98784" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101269" />
                    <RANKING order="2" place="2" resultid="100629" />
                    <RANKING order="3" place="3" resultid="102456" />
                    <RANKING order="4" place="4" resultid="103099" />
                    <RANKING order="5" place="5" resultid="100587" />
                    <RANKING order="6" place="6" resultid="103094" />
                    <RANKING order="7" place="7" resultid="102834" />
                    <RANKING order="8" place="8" resultid="103461" />
                    <RANKING order="9" place="9" resultid="102727" />
                    <RANKING order="10" place="10" resultid="103111" />
                    <RANKING order="11" place="-1" resultid="101309" />
                    <RANKING order="12" place="-1" resultid="102754" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98787" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103087" />
                    <RANKING order="2" place="2" resultid="102540" />
                    <RANKING order="3" place="3" resultid="103337" />
                    <RANKING order="4" place="4" resultid="102719" />
                    <RANKING order="5" place="5" resultid="105020" />
                    <RANKING order="6" place="6" resultid="103082" />
                    <RANKING order="7" place="7" resultid="100934" />
                    <RANKING order="8" place="8" resultid="102787" />
                    <RANKING order="9" place="9" resultid="102778" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98786" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102533" />
                    <RANKING order="2" place="2" resultid="100669" />
                    <RANKING order="3" place="3" resultid="100951" />
                    <RANKING order="4" place="4" resultid="102461" />
                    <RANKING order="5" place="5" resultid="101433" />
                    <RANKING order="6" place="6" resultid="100443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98789" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101567" />
                    <RANKING order="2" place="2" resultid="101493" />
                    <RANKING order="3" place="3" resultid="101283" />
                    <RANKING order="4" place="4" resultid="101452" />
                    <RANKING order="5" place="5" resultid="101838" />
                    <RANKING order="6" place="6" resultid="103381" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98788" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100685" />
                    <RANKING order="2" place="2" resultid="102740" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98791" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103077" />
                    <RANKING order="2" place="2" resultid="100463" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98793" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="98792" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="98795" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105113" daytime="16:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105114" daytime="16:03" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105115" daytime="16:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105116" daytime="16:07" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="105117" daytime="16:09" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="105118" daytime="16:11" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="105119" daytime="16:13" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="105120" daytime="16:15" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="105121" daytime="16:17" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="98798" daytime="16:20" gender="M" number="2" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99677" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100898" />
                    <RANKING order="2" place="2" resultid="103042" />
                    <RANKING order="3" place="3" resultid="102409" />
                    <RANKING order="4" place="4" resultid="103028" />
                    <RANKING order="5" place="5" resultid="101045" />
                    <RANKING order="6" place="6" resultid="102418" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99678" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102275" />
                    <RANKING order="2" place="2" resultid="105108" />
                    <RANKING order="3" place="3" resultid="101150" />
                    <RANKING order="4" place="4" resultid="101725" />
                    <RANKING order="5" place="5" resultid="100157" />
                    <RANKING order="6" place="6" resultid="101855" />
                    <RANKING order="7" place="7" resultid="103366" />
                    <RANKING order="8" place="8" resultid="100317" />
                    <RANKING order="9" place="9" resultid="100295" />
                    <RANKING order="10" place="10" resultid="101821" />
                    <RANKING order="11" place="11" resultid="101315" />
                    <RANKING order="12" place="12" resultid="101300" />
                    <RANKING order="13" place="13" resultid="101102" />
                    <RANKING order="14" place="14" resultid="101318" />
                    <RANKING order="15" place="-1" resultid="100663" />
                    <RANKING order="16" place="-1" resultid="101207" />
                    <RANKING order="17" place="-1" resultid="101228" />
                    <RANKING order="18" place="-1" resultid="101760" />
                    <RANKING order="19" place="-1" resultid="102484" />
                    <RANKING order="20" place="-1" resultid="102862" />
                    <RANKING order="21" place="-1" resultid="103007" />
                    <RANKING order="22" place="-1" resultid="103437" />
                    <RANKING order="23" place="-1" resultid="105105" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99679" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101766" />
                    <RANKING order="2" place="2" resultid="103317" />
                    <RANKING order="3" place="3" resultid="100424" />
                    <RANKING order="4" place="4" resultid="102987" />
                    <RANKING order="5" place="5" resultid="100277" />
                    <RANKING order="6" place="6" resultid="102813" />
                    <RANKING order="7" place="7" resultid="102180" />
                    <RANKING order="8" place="8" resultid="102367" />
                    <RANKING order="9" place="9" resultid="102891" />
                    <RANKING order="10" place="10" resultid="102474" />
                    <RANKING order="11" place="11" resultid="102206" />
                    <RANKING order="12" place="12" resultid="101049" />
                    <RANKING order="13" place="13" resultid="100152" />
                    <RANKING order="14" place="14" resultid="104372" />
                    <RANKING order="15" place="15" resultid="101649" />
                    <RANKING order="16" place="16" resultid="102886" />
                    <RANKING order="17" place="17" resultid="102212" />
                    <RANKING order="18" place="18" resultid="100304" />
                    <RANKING order="19" place="19" resultid="101249" />
                    <RANKING order="20" place="-1" resultid="105111" />
                    <RANKING order="21" place="-1" resultid="100324" />
                    <RANKING order="22" place="-1" resultid="101220" />
                    <RANKING order="23" place="-1" resultid="101792" />
                    <RANKING order="24" place="-1" resultid="103451" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99680" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102153" />
                    <RANKING order="2" place="2" resultid="100751" />
                    <RANKING order="3" place="3" resultid="102880" />
                    <RANKING order="4" place="4" resultid="100831" />
                    <RANKING order="5" place="5" resultid="103047" />
                    <RANKING order="6" place="6" resultid="101919" />
                    <RANKING order="7" place="7" resultid="101132" />
                    <RANKING order="8" place="8" resultid="102471" />
                    <RANKING order="9" place="9" resultid="101253" />
                    <RANKING order="10" place="10" resultid="100412" />
                    <RANKING order="11" place="11" resultid="102098" />
                    <RANKING order="12" place="12" resultid="102579" />
                    <RANKING order="13" place="13" resultid="103446" />
                    <RANKING order="14" place="14" resultid="100291" />
                    <RANKING order="15" place="15" resultid="102477" />
                    <RANKING order="16" place="16" resultid="101598" />
                    <RANKING order="17" place="17" resultid="102491" />
                    <RANKING order="18" place="18" resultid="100219" />
                    <RANKING order="19" place="19" resultid="100805" />
                    <RANKING order="20" place="20" resultid="101712" />
                    <RANKING order="21" place="21" resultid="100104" />
                    <RANKING order="22" place="22" resultid="101066" />
                    <RANKING order="23" place="23" resultid="102252" />
                    <RANKING order="24" place="-1" resultid="102913" />
                    <RANKING order="25" place="-1" resultid="101264" />
                    <RANKING order="26" place="-1" resultid="101674" />
                    <RANKING order="27" place="-1" resultid="102962" />
                    <RANKING order="28" place="-1" resultid="103256" />
                    <RANKING order="29" place="-1" resultid="103262" />
                    <RANKING order="30" place="-1" resultid="100205" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99681" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101351" />
                    <RANKING order="2" place="2" resultid="100760" />
                    <RANKING order="3" place="3" resultid="101401" />
                    <RANKING order="4" place="4" resultid="103510" />
                    <RANKING order="5" place="5" resultid="101186" />
                    <RANKING order="6" place="6" resultid="103251" />
                    <RANKING order="7" place="7" resultid="101211" />
                    <RANKING order="8" place="8" resultid="100210" />
                    <RANKING order="9" place="9" resultid="105072" />
                    <RANKING order="10" place="10" resultid="102510" />
                    <RANKING order="11" place="11" resultid="100241" />
                    <RANKING order="12" place="12" resultid="103590" />
                    <RANKING order="13" place="13" resultid="100199" />
                    <RANKING order="14" place="14" resultid="100778" />
                    <RANKING order="15" place="15" resultid="102481" />
                    <RANKING order="16" place="16" resultid="102270" />
                    <RANKING order="17" place="17" resultid="103582" />
                    <RANKING order="18" place="18" resultid="100975" />
                    <RANKING order="19" place="-1" resultid="100958" />
                    <RANKING order="20" place="-1" resultid="101203" />
                    <RANKING order="21" place="-1" resultid="101928" />
                    <RANKING order="22" place="-1" resultid="101941" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99682" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="104999" />
                    <RANKING order="2" place="2" resultid="101829" />
                    <RANKING order="3" place="3" resultid="100477" />
                    <RANKING order="4" place="4" resultid="104972" />
                    <RANKING order="5" place="5" resultid="101750" />
                    <RANKING order="6" place="6" resultid="104964" />
                    <RANKING order="7" place="7" resultid="101558" />
                    <RANKING order="8" place="8" resultid="101036" />
                    <RANKING order="9" place="9" resultid="100823" />
                    <RANKING order="10" place="10" resultid="100458" />
                    <RANKING order="11" place="11" resultid="103240" />
                    <RANKING order="12" place="12" resultid="101696" />
                    <RANKING order="13" place="13" resultid="103233" />
                    <RANKING order="14" place="14" resultid="100452" />
                    <RANKING order="15" place="15" resultid="101418" />
                    <RANKING order="16" place="16" resultid="103573" />
                    <RANKING order="17" place="17" resultid="102850" />
                    <RANKING order="18" place="18" resultid="105078" />
                    <RANKING order="19" place="19" resultid="100395" />
                    <RANKING order="20" place="20" resultid="102468" />
                    <RANKING order="21" place="20" resultid="103228" />
                    <RANKING order="22" place="22" resultid="103554" />
                    <RANKING order="23" place="23" resultid="101638" />
                    <RANKING order="24" place="24" resultid="100857" />
                    <RANKING order="25" place="-1" resultid="101423" />
                    <RANKING order="26" place="-1" resultid="101260" />
                    <RANKING order="27" place="-1" resultid="101339" />
                    <RANKING order="28" place="-1" resultid="101778" />
                    <RANKING order="29" place="-1" resultid="101999" />
                    <RANKING order="30" place="-1" resultid="103071" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99683" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101608" />
                    <RANKING order="2" place="2" resultid="102855" />
                    <RANKING order="3" place="3" resultid="102383" />
                    <RANKING order="4" place="4" resultid="100127" />
                    <RANKING order="5" place="5" resultid="101499" />
                    <RANKING order="6" place="6" resultid="105043" />
                    <RANKING order="7" place="7" resultid="101478" />
                    <RANKING order="8" place="8" resultid="101631" />
                    <RANKING order="9" place="9" resultid="103210" />
                    <RANKING order="10" place="10" resultid="103217" />
                    <RANKING order="11" place="11" resultid="103204" />
                    <RANKING order="12" place="12" resultid="101735" />
                    <RANKING order="13" place="-1" resultid="101657" />
                    <RANKING order="14" place="-1" resultid="103223" />
                    <RANKING order="15" place="-1" resultid="103321" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99684" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103502" />
                    <RANKING order="2" place="2" resultid="102259" />
                    <RANKING order="3" place="3" resultid="102827" />
                    <RANKING order="4" place="4" resultid="100989" />
                    <RANKING order="5" place="5" resultid="103604" />
                    <RANKING order="6" place="6" resultid="102264" />
                    <RANKING order="7" place="7" resultid="100942" />
                    <RANKING order="8" place="8" resultid="103069" />
                    <RANKING order="9" place="9" resultid="101666" />
                    <RANKING order="10" place="10" resultid="103193" />
                    <RANKING order="11" place="11" resultid="103360" />
                    <RANKING order="12" place="-1" resultid="103187" />
                    <RANKING order="13" place="-1" resultid="100620" />
                    <RANKING order="14" place="-1" resultid="100666" />
                    <RANKING order="15" place="-1" resultid="100928" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99685" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100269" />
                    <RANKING order="2" place="2" resultid="102193" />
                    <RANKING order="3" place="3" resultid="101770" />
                    <RANKING order="4" place="4" resultid="101057" />
                    <RANKING order="5" place="4" resultid="101446" />
                    <RANKING order="6" place="6" resultid="103181" />
                    <RANKING order="7" place="7" resultid="101027" />
                    <RANKING order="8" place="8" resultid="103034" />
                    <RANKING order="9" place="9" resultid="103176" />
                    <RANKING order="10" place="10" resultid="102562" />
                    <RANKING order="11" place="11" resultid="102634" />
                    <RANKING order="12" place="-1" resultid="101322" />
                    <RANKING order="13" place="-1" resultid="103170" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99686" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102525" />
                    <RANKING order="2" place="2" resultid="100695" />
                    <RANKING order="3" place="3" resultid="100349" />
                    <RANKING order="4" place="4" resultid="100769" />
                    <RANKING order="5" place="5" resultid="100573" />
                    <RANKING order="6" place="6" resultid="101484" />
                    <RANKING order="7" place="7" resultid="103372" />
                    <RANKING order="8" place="8" resultid="103148" />
                    <RANKING order="9" place="9" resultid="100569" />
                    <RANKING order="10" place="10" resultid="103162" />
                    <RANKING order="11" place="11" resultid="100084" />
                    <RANKING order="12" place="12" resultid="100564" />
                    <RANKING order="13" place="13" resultid="101739" />
                    <RANKING order="14" place="14" resultid="101278" />
                    <RANKING order="15" place="15" resultid="100717" />
                    <RANKING order="16" place="16" resultid="102946" />
                    <RANKING order="17" place="17" resultid="103548" />
                    <RANKING order="18" place="-1" resultid="102126" />
                    <RANKING order="19" place="-1" resultid="103154" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99687" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101676" />
                    <RANKING order="2" place="2" resultid="102555" />
                    <RANKING order="3" place="3" resultid="102974" />
                    <RANKING order="4" place="4" resultid="102139" />
                    <RANKING order="5" place="5" resultid="102518" />
                    <RANKING order="6" place="-1" resultid="103407" />
                    <RANKING order="7" place="-1" resultid="100367" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99688" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100402" />
                    <RANKING order="2" place="2" resultid="100978" />
                    <RANKING order="3" place="3" resultid="102134" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99689" agemax="84" agemin="80" name="KAT.L, 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100994" />
                    <RANKING order="2" place="2" resultid="104988" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99690" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99691" agemax="94" agemin="90" name="KAT.N, 90-94 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100615" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105123" daytime="16:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105124" daytime="16:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105125" daytime="16:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105126" daytime="16:27" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="105127" daytime="16:29" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="105128" daytime="16:31" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="105129" daytime="16:33" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="105130" daytime="16:35" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="105131" daytime="16:37" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="105132" daytime="16:39" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="105133" daytime="16:42" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="105134" daytime="16:44" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="105135" daytime="16:46" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="105136" daytime="16:48" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="105137" daytime="16:49" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="105138" daytime="16:51" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="105139" daytime="16:53" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="105140" daytime="16:55" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="105141" daytime="16:57" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="105142" daytime="16:59" number="20" order="20" status="OFFICIAL" />
                <HEAT heatid="105143" daytime="17:01" number="21" order="21" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="98814" daytime="17:04" gender="F" number="3" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99692" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102997" />
                    <RANKING order="2" place="2" resultid="100906" />
                    <RANKING order="3" place="3" resultid="100887" />
                    <RANKING order="4" place="-1" resultid="102105" />
                    <RANKING order="5" place="-1" resultid="103058" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99693" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103138" />
                    <RANKING order="2" place="2" resultid="103390" />
                    <RANKING order="3" place="3" resultid="102172" />
                    <RANKING order="4" place="4" resultid="103559" />
                    <RANKING order="5" place="5" resultid="101591" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99694" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103354" />
                    <RANKING order="2" place="2" resultid="100580" />
                    <RANKING order="3" place="-1" resultid="102955" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99695" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102091" />
                    <RANKING order="2" place="-1" resultid="101304" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99696" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100608" />
                    <RANKING order="2" place="2" resultid="100965" />
                    <RANKING order="3" place="3" resultid="101799" />
                    <RANKING order="4" place="4" resultid="103131" />
                    <RANKING order="5" place="5" resultid="102896" />
                    <RANKING order="6" place="6" resultid="103343" />
                    <RANKING order="7" place="-1" resultid="100699" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99697" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100549" />
                    <RANKING order="2" place="2" resultid="100815" />
                    <RANKING order="3" place="3" resultid="103493" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99698" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101457" />
                    <RANKING order="2" place="2" resultid="103112" />
                    <RANKING order="3" place="3" resultid="103462" />
                    <RANKING order="4" place="-1" resultid="102548" />
                    <RANKING order="5" place="-1" resultid="102755" />
                    <RANKING order="6" place="-1" resultid="103105" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99699" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101990" />
                    <RANKING order="2" place="2" resultid="103088" />
                    <RANKING order="3" place="3" resultid="102541" />
                    <RANKING order="4" place="4" resultid="102788" />
                    <RANKING order="5" place="5" resultid="102779" />
                    <RANKING order="6" place="-1" resultid="102697" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99700" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102711" />
                    <RANKING order="2" place="2" resultid="101434" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99701" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103382" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99702" agemax="74" agemin="70" name="KAT.J, 70-74 lat" />
                <AGEGROUP agegroupid="99703" agemax="79" agemin="75" name="KAT.K, 75-79 lat" />
                <AGEGROUP agegroupid="99704" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99705" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99706" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105144" daytime="17:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105145" daytime="17:11" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105146" daytime="17:16" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105147" daytime="17:20" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="98830" daytime="17:25" gender="M" number="4" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99707" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100899" />
                    <RANKING order="2" place="2" resultid="102901" />
                    <RANKING order="3" place="3" resultid="100970" />
                    <RANKING order="4" place="4" resultid="104954" />
                    <RANKING order="5" place="5" resultid="100796" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99708" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101144" />
                    <RANKING order="2" place="2" resultid="100158" />
                    <RANKING order="3" place="3" resultid="103022" />
                    <RANKING order="4" place="4" resultid="100284" />
                    <RANKING order="5" place="-1" resultid="102863" />
                    <RANKING order="6" place="-1" resultid="103008" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99709" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102062" />
                    <RANKING order="2" place="2" resultid="101008" />
                    <RANKING order="3" place="3" resultid="100278" />
                    <RANKING order="4" place="4" resultid="103537" />
                    <RANKING order="5" place="5" resultid="102374" />
                    <RANKING order="6" place="6" resultid="102181" />
                    <RANKING order="7" place="7" resultid="102988" />
                    <RANKING order="8" place="8" resultid="102145" />
                    <RANKING order="9" place="-1" resultid="101650" />
                    <RANKING order="10" place="-1" resultid="103452" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99710" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102154" />
                    <RANKING order="2" place="2" resultid="102162" />
                    <RANKING order="3" place="3" resultid="101920" />
                    <RANKING order="4" place="4" resultid="100832" />
                    <RANKING order="5" place="5" resultid="100752" />
                    <RANKING order="6" place="6" resultid="101195" />
                    <RANKING order="7" place="7" resultid="101713" />
                    <RANKING order="8" place="8" resultid="100595" />
                    <RANKING order="9" place="9" resultid="103048" />
                    <RANKING order="10" place="10" resultid="104399" />
                    <RANKING order="11" place="11" resultid="100105" />
                    <RANKING order="12" place="12" resultid="102247" />
                    <RANKING order="13" place="-1" resultid="102963" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99711" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100761" />
                    <RANKING order="2" place="2" resultid="101402" />
                    <RANKING order="3" place="3" resultid="101212" />
                    <RANKING order="4" place="4" resultid="101187" />
                    <RANKING order="5" place="5" resultid="103511" />
                    <RANKING order="6" place="6" resultid="101178" />
                    <RANKING order="7" place="7" resultid="101413" />
                    <RANKING order="8" place="8" resultid="101473" />
                    <RANKING order="9" place="9" resultid="100188" />
                    <RANKING order="10" place="10" resultid="105073" />
                    <RANKING order="11" place="11" resultid="100779" />
                    <RANKING order="12" place="-1" resultid="101234" />
                    <RANKING order="13" place="-1" resultid="101929" />
                    <RANKING order="14" place="-1" resultid="101935" />
                    <RANKING order="15" place="-1" resultid="102980" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99712" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101830" />
                    <RANKING order="2" place="2" resultid="105000" />
                    <RANKING order="3" place="3" resultid="100720" />
                    <RANKING order="4" place="4" resultid="104973" />
                    <RANKING order="5" place="5" resultid="101697" />
                    <RANKING order="6" place="6" resultid="101559" />
                    <RANKING order="7" place="7" resultid="103574" />
                    <RANKING order="8" place="8" resultid="102840" />
                    <RANKING order="9" place="9" resultid="101312" />
                    <RANKING order="10" place="10" resultid="101261" />
                    <RANKING order="11" place="11" resultid="100915" />
                    <RANKING order="12" place="12" resultid="103596" />
                    <RANKING order="13" place="13" resultid="101779" />
                    <RANKING order="14" place="-1" resultid="100858" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99713" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100128" />
                    <RANKING order="2" place="2" resultid="104978" />
                    <RANKING order="3" place="3" resultid="101442" />
                    <RANKING order="4" place="4" resultid="100787" />
                    <RANKING order="5" place="5" resultid="101632" />
                    <RANKING order="6" place="6" resultid="102361" />
                    <RANKING order="7" place="7" resultid="103015" />
                    <RANKING order="8" place="8" resultid="103543" />
                    <RANKING order="9" place="-1" resultid="100120" />
                    <RANKING order="10" place="-1" resultid="101658" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99714" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103503" />
                    <RANKING order="2" place="2" resultid="100621" />
                    <RANKING order="3" place="3" resultid="100555" />
                    <RANKING order="4" place="4" resultid="102568" />
                    <RANKING order="5" place="5" resultid="101157" />
                    <RANKING order="6" place="6" resultid="100600" />
                    <RANKING order="7" place="7" resultid="101667" />
                    <RANKING order="8" place="8" resultid="102027" />
                    <RANKING order="9" place="9" resultid="102045" />
                    <RANKING order="10" place="10" resultid="102033" />
                    <RANKING order="11" place="11" resultid="101087" />
                    <RANKING order="12" place="-1" resultid="102011" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99715" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101577" />
                    <RANKING order="2" place="2" resultid="102201" />
                    <RANKING order="3" place="3" resultid="102504" />
                    <RANKING order="4" place="4" resultid="102194" />
                    <RANKING order="5" place="5" resultid="100376" />
                    <RANKING order="6" place="6" resultid="105008" />
                    <RANKING order="7" place="7" resultid="102734" />
                    <RANKING order="8" place="8" resultid="102114" />
                    <RANKING order="9" place="9" resultid="102121" />
                    <RANKING order="10" place="10" resultid="102635" />
                    <RANKING order="11" place="11" resultid="100385" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99716" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100770" />
                    <RANKING order="2" place="2" resultid="100350" />
                    <RANKING order="3" place="3" resultid="103163" />
                    <RANKING order="4" place="4" resultid="101288" />
                    <RANKING order="5" place="5" resultid="105054" />
                    <RANKING order="6" place="6" resultid="102947" />
                    <RANKING order="7" place="7" resultid="101015" />
                    <RANKING order="8" place="-1" resultid="102127" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99717" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102556" />
                    <RANKING order="2" place="2" resultid="100368" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99718" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102745" />
                    <RANKING order="2" place="2" resultid="100403" />
                    <RANKING order="3" place="3" resultid="101582" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99719" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99720" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99721" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105148" daytime="17:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105149" daytime="17:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105150" daytime="17:38" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105151" daytime="17:43" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="105152" daytime="17:48" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="105153" daytime="17:53" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="105154" daytime="17:57" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="105155" daytime="18:02" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="105156" daytime="18:06" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="105157" daytime="18:10" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="105158" daytime="18:14" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="98846" daytime="18:19" gender="X" number="5" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="98847" agemax="96" agemin="80" name="KAT.0, 80-96 lat" calculate="TOTAL" />
                <AGEGROUP agegroupid="98848" agemax="119" agemin="100" name="KAT.A, 100-119 lat" calculate="TOTAL" />
                <AGEGROUP agegroupid="98849" agemax="159" agemin="120" name="KAT.B, 120-159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102294" />
                    <RANKING order="2" place="2" resultid="101869" />
                    <RANKING order="3" place="3" resultid="102216" />
                    <RANKING order="4" place="4" resultid="100248" />
                    <RANKING order="5" place="5" resultid="104098" />
                    <RANKING order="6" place="6" resultid="101868" />
                    <RANKING order="7" place="7" resultid="103420" />
                    <RANKING order="8" place="8" resultid="101881" />
                    <RANKING order="9" place="-1" resultid="101360" />
                    <RANKING order="10" place="-1" resultid="103281" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98850" agemax="199" agemin="160" name="KAT.C,160-199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101361" />
                    <RANKING order="2" place="2" resultid="103418" />
                    <RANKING order="3" place="3" resultid="103266" />
                    <RANKING order="4" place="4" resultid="100634" />
                    <RANKING order="5" place="5" resultid="100249" />
                    <RANKING order="6" place="6" resultid="102488" />
                    <RANKING order="7" place="-1" resultid="102585" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98851" agemax="239" agemin="200" name="KAT.D, 200-239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103279" />
                    <RANKING order="2" place="2" resultid="104097" />
                    <RANKING order="3" place="3" resultid="100636" />
                    <RANKING order="4" place="4" resultid="105065" />
                    <RANKING order="5" place="-1" resultid="105039" />
                    <RANKING order="6" place="-1" resultid="101363" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98852" agemax="279" agemin="240" name="KAT.E, 240-279 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103268" />
                    <RANKING order="2" place="2" resultid="100731" />
                    <RANKING order="3" place="3" resultid="103416" />
                    <RANKING order="4" place="4" resultid="101365" />
                    <RANKING order="5" place="-1" resultid="102766" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="98853" agemax="-1" agemin="280" name="KAT.F, 280+ lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100730" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105159" daytime="18:19" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105160" daytime="18:24" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105161" daytime="18:28" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="98863" daytime="18:32" gender="F" number="6" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99722" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103613" />
                    <RANKING order="2" place="2" resultid="100311" />
                    <RANKING order="3" place="3" resultid="102106" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99723" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102285" />
                    <RANKING order="2" place="2" resultid="101138" />
                    <RANKING order="3" place="3" resultid="102497" />
                    <RANKING order="4" place="4" resultid="100432" />
                    <RANKING order="5" place="-1" resultid="101846" />
                    <RANKING order="6" place="-1" resultid="101346" />
                    <RANKING order="7" place="-1" resultid="101617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99724" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103531" />
                    <RANKING order="2" place="2" resultid="103523" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99725" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100923" />
                    <RANKING order="2" place="2" resultid="100164" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99726" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100700" />
                    <RANKING order="2" place="2" resultid="100966" />
                    <RANKING order="3" place="3" resultid="100233" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99727" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="105014" />
                    <RANKING order="2" place="2" resultid="100550" />
                    <RANKING order="3" place="3" resultid="103494" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99728" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102835" />
                    <RANKING order="2" place="2" resultid="100437" />
                    <RANKING order="3" place="-1" resultid="100540" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99729" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101991" />
                    <RANKING order="2" place="2" resultid="102698" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99730" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100444" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99731" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101839" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99732" agemax="74" agemin="70" name="KAT.J, 70-74 lat" />
                <AGEGROUP agegroupid="99733" agemax="79" agemin="75" name="KAT.K, 75-79 lat" />
                <AGEGROUP agegroupid="99734" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99735" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99736" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105404" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105405" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105406" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="98891" daytime="19:19" gender="M" number="7" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99737" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100797" />
                    <RANKING order="2" place="2" resultid="104955" />
                    <RANKING order="3" place="3" resultid="100681" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99738" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102276" />
                    <RANKING order="2" place="2" resultid="105089" />
                    <RANKING order="3" place="3" resultid="100285" />
                    <RANKING order="4" place="4" resultid="101316" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99739" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101009" />
                    <RANKING order="2" place="2" resultid="102375" />
                    <RANKING order="3" place="3" resultid="100866" />
                    <RANKING order="4" place="-1" resultid="101050" />
                    <RANKING order="5" place="-1" resultid="101767" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99740" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102881" />
                    <RANKING order="2" place="2" resultid="102163" />
                    <RANKING order="3" place="3" resultid="100806" />
                    <RANKING order="4" place="4" resultid="102801" />
                    <RANKING order="5" place="-1" resultid="102006" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99741" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103396" />
                    <RANKING order="2" place="2" resultid="105034" />
                    <RANKING order="3" place="3" resultid="101408" />
                    <RANKING order="4" place="4" resultid="102069" />
                    <RANKING order="5" place="5" resultid="101604" />
                    <RANKING order="6" place="-1" resultid="104996" />
                    <RANKING order="7" place="-1" resultid="100211" />
                    <RANKING order="8" place="-1" resultid="101942" />
                    <RANKING order="9" place="-1" resultid="102982" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99742" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101692" />
                    <RANKING order="2" place="2" resultid="103246" />
                    <RANKING order="3" place="3" resultid="104965" />
                    <RANKING order="4" place="4" resultid="102355" />
                    <RANKING order="5" place="5" resultid="105079" />
                    <RANKING order="6" place="6" resultid="102845" />
                    <RANKING order="7" place="-1" resultid="103234" />
                    <RANKING order="8" place="-1" resultid="103567" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99743" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="105044" />
                    <RANKING order="2" place="2" resultid="104388" />
                    <RANKING order="3" place="3" resultid="100788" />
                    <RANKING order="4" place="4" resultid="102393" />
                    <RANKING order="5" place="5" resultid="103211" />
                    <RANKING order="6" place="6" resultid="102349" />
                    <RANKING order="7" place="7" resultid="103205" />
                    <RANKING order="8" place="8" resultid="103322" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99744" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102012" />
                    <RANKING order="2" place="2" resultid="100943" />
                    <RANKING order="3" place="3" resultid="101158" />
                    <RANKING order="4" place="4" resultid="103194" />
                    <RANKING order="5" place="-1" resultid="102995" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99745" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101771" />
                    <RANKING order="2" place="2" resultid="100377" />
                    <RANKING order="3" place="3" resultid="101058" />
                    <RANKING order="4" place="4" resultid="100386" />
                    <RANKING order="5" place="-1" resultid="100270" />
                    <RANKING order="6" place="-1" resultid="101028" />
                    <RANKING order="7" place="-1" resultid="102021" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99746" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101485" />
                    <RANKING order="2" place="2" resultid="105055" />
                    <RANKING order="3" place="3" resultid="100085" />
                    <RANKING order="4" place="4" resultid="103373" />
                    <RANKING order="5" place="-1" resultid="103155" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99747" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102975" />
                    <RANKING order="2" place="2" resultid="103408" />
                    <RANKING order="3" place="3" resultid="101677" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99748" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100691" />
                    <RANKING order="2" place="2" resultid="100979" />
                    <RANKING order="3" place="3" resultid="101583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99749" agemax="84" agemin="80" name="KAT.L, 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="104992" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99750" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99751" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105420" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105421" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105422" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105423" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="105424" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="105425" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2014-06-28" daytime="09:00" number="2" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="98907" daytime="09:00" gender="F" number="8" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99752" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100312" />
                    <RANKING order="2" place="2" resultid="103470" />
                    <RANKING order="3" place="3" resultid="102414" />
                    <RANKING order="4" place="4" resultid="100888" />
                    <RANKING order="5" place="5" resultid="103059" />
                    <RANKING order="6" place="6" resultid="100907" />
                    <RANKING order="7" place="7" resultid="104377" />
                    <RANKING order="8" place="8" resultid="103476" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99753" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101139" />
                    <RANKING order="2" place="2" resultid="103391" />
                    <RANKING order="3" place="3" resultid="102944" />
                    <RANKING order="4" place="4" resultid="102173" />
                    <RANKING order="5" place="5" resultid="101166" />
                    <RANKING order="6" place="6" resultid="103027" />
                    <RANKING order="7" place="7" resultid="101787" />
                    <RANKING order="8" place="-1" resultid="101847" />
                    <RANKING order="9" place="-1" resultid="102389" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99754" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101085" />
                    <RANKING order="2" place="2" resultid="103519" />
                    <RANKING order="3" place="3" resultid="100581" />
                    <RANKING order="4" place="-1" resultid="102956" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99755" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100165" />
                    <RANKING order="2" place="2" resultid="101703" />
                    <RANKING order="3" place="3" resultid="102092" />
                    <RANKING order="4" place="4" resultid="100173" />
                    <RANKING order="5" place="5" resultid="101686" />
                    <RANKING order="6" place="-1" resultid="101305" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99756" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100609" />
                    <RANKING order="2" place="2" resultid="103331" />
                    <RANKING order="3" place="3" resultid="103125" />
                    <RANKING order="4" place="4" resultid="100234" />
                    <RANKING order="5" place="5" resultid="102897" />
                    <RANKING order="6" place="-1" resultid="103344" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99757" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100727" />
                    <RANKING order="2" place="2" resultid="103348" />
                    <RANKING order="3" place="3" resultid="103427" />
                    <RANKING order="4" place="4" resultid="101072" />
                    <RANKING order="5" place="5" resultid="105031" />
                    <RANKING order="6" place="6" resultid="100872" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99758" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103100" />
                    <RANKING order="2" place="2" resultid="101270" />
                    <RANKING order="3" place="3" resultid="100588" />
                    <RANKING order="4" place="4" resultid="102457" />
                    <RANKING order="5" place="5" resultid="101458" />
                    <RANKING order="6" place="6" resultid="102728" />
                    <RANKING order="7" place="7" resultid="103113" />
                    <RANKING order="8" place="-1" resultid="103106" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99759" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101992" />
                    <RANKING order="2" place="2" resultid="101294" />
                    <RANKING order="3" place="3" resultid="102542" />
                    <RANKING order="4" place="4" resultid="105021" />
                    <RANKING order="5" place="5" resultid="102789" />
                    <RANKING order="6" place="-1" resultid="100935" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99760" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102462" />
                    <RANKING order="2" place="2" resultid="102534" />
                    <RANKING order="3" place="3" resultid="100952" />
                    <RANKING order="4" place="4" resultid="100445" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99761" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101568" />
                    <RANKING order="2" place="2" resultid="101494" />
                    <RANKING order="3" place="3" resultid="101284" />
                    <RANKING order="4" place="-1" resultid="101840" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99762" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100686" />
                    <RANKING order="2" place="2" resultid="102741" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99763" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100464" />
                    <RANKING order="2" place="2" resultid="101573" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99764" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99765" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99766" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105172" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105173" daytime="09:03" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105174" daytime="09:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105175" daytime="09:08" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="105176" daytime="09:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="105177" daytime="09:13" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="105178" daytime="09:15" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="98924" daytime="09:17" gender="M" number="9" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99767" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100971" />
                    <RANKING order="2" place="2" resultid="102410" />
                    <RANKING order="3" place="3" resultid="102806" />
                    <RANKING order="4" place="4" resultid="100798" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99768" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="105090" />
                    <RANKING order="2" place="2" resultid="101002" />
                    <RANKING order="3" place="3" resultid="101145" />
                    <RANKING order="4" place="4" resultid="102277" />
                    <RANKING order="5" place="5" resultid="103442" />
                    <RANKING order="6" place="6" resultid="101645" />
                    <RANKING order="7" place="7" resultid="100296" />
                    <RANKING order="8" place="8" resultid="101856" />
                    <RANKING order="9" place="-1" resultid="102864" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99769" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102063" />
                    <RANKING order="2" place="2" resultid="102368" />
                    <RANKING order="3" place="3" resultid="102475" />
                    <RANKING order="4" place="4" resultid="102182" />
                    <RANKING order="5" place="5" resultid="102887" />
                    <RANKING order="6" place="6" resultid="102207" />
                    <RANKING order="7" place="7" resultid="101651" />
                    <RANKING order="8" place="8" resultid="101805" />
                    <RANKING order="9" place="-1" resultid="100305" />
                    <RANKING order="10" place="-1" resultid="102146" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99770" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102821" />
                    <RANKING order="2" place="2" resultid="100753" />
                    <RANKING order="3" place="3" resultid="102164" />
                    <RANKING order="4" place="4" resultid="103049" />
                    <RANKING order="5" place="5" resultid="101196" />
                    <RANKING order="6" place="6" resultid="102099" />
                    <RANKING order="7" place="7" resultid="104400" />
                    <RANKING order="8" place="8" resultid="100206" />
                    <RANKING order="9" place="9" resultid="102580" />
                    <RANKING order="10" place="10" resultid="100106" />
                    <RANKING order="11" place="11" resultid="102253" />
                    <RANKING order="12" place="-1" resultid="101815" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99771" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101188" />
                    <RANKING order="2" place="2" resultid="101474" />
                    <RANKING order="3" place="3" resultid="100762" />
                    <RANKING order="4" place="4" resultid="101179" />
                    <RANKING order="5" place="5" resultid="101414" />
                    <RANKING order="6" place="6" resultid="100212" />
                    <RANKING order="7" place="7" resultid="102271" />
                    <RANKING order="8" place="8" resultid="102511" />
                    <RANKING order="9" place="-1" resultid="100959" />
                    <RANKING order="10" place="-1" resultid="101930" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99772" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100721" />
                    <RANKING order="2" place="2" resultid="101831" />
                    <RANKING order="3" place="3" resultid="101698" />
                    <RANKING order="4" place="4" resultid="104966" />
                    <RANKING order="5" place="5" resultid="100459" />
                    <RANKING order="6" place="6" resultid="103241" />
                    <RANKING order="7" place="7" resultid="101037" />
                    <RANKING order="8" place="8" resultid="102356" />
                    <RANKING order="9" place="9" resultid="103490" />
                    <RANKING order="10" place="10" resultid="103575" />
                    <RANKING order="11" place="11" resultid="100824" />
                    <RANKING order="12" place="12" resultid="100916" />
                    <RANKING order="13" place="13" resultid="101313" />
                    <RANKING order="14" place="14" resultid="103555" />
                    <RANKING order="15" place="15" resultid="103597" />
                    <RANKING order="16" place="-1" resultid="102000" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99773" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101479" />
                    <RANKING order="2" place="2" resultid="102856" />
                    <RANKING order="3" place="3" resultid="100659" />
                    <RANKING order="4" place="4" resultid="103016" />
                    <RANKING order="5" place="5" resultid="103218" />
                    <RANKING order="6" place="-1" resultid="103212" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99774" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103504" />
                    <RANKING order="2" place="2" resultid="102828" />
                    <RANKING order="3" place="3" resultid="100622" />
                    <RANKING order="4" place="4" resultid="103605" />
                    <RANKING order="5" place="5" resultid="103188" />
                    <RANKING order="6" place="6" resultid="101159" />
                    <RANKING order="7" place="7" resultid="102569" />
                    <RANKING order="8" place="8" resultid="102028" />
                    <RANKING order="9" place="9" resultid="101668" />
                    <RANKING order="10" place="10" resultid="102034" />
                    <RANKING order="11" place="11" resultid="101088" />
                    <RANKING order="12" place="12" resultid="103361" />
                    <RANKING order="13" place="-1" resultid="100673" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99775" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101274" />
                    <RANKING order="2" place="2" resultid="101059" />
                    <RANKING order="3" place="3" resultid="101772" />
                    <RANKING order="4" place="4" resultid="100271" />
                    <RANKING order="5" place="5" resultid="100378" />
                    <RANKING order="6" place="6" resultid="101029" />
                    <RANKING order="7" place="7" resultid="103182" />
                    <RANKING order="8" place="8" resultid="102563" />
                    <RANKING order="9" place="-1" resultid="103171" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99776" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102526" />
                    <RANKING order="2" place="2" resultid="101486" />
                    <RANKING order="3" place="3" resultid="100771" />
                    <RANKING order="4" place="4" resultid="100677" />
                    <RANKING order="5" place="5" resultid="103149" />
                    <RANKING order="6" place="6" resultid="101279" />
                    <RANKING order="7" place="7" resultid="102948" />
                    <RANKING order="8" place="8" resultid="102128" />
                    <RANKING order="9" place="9" resultid="101335" />
                    <RANKING order="10" place="10" resultid="103402" />
                    <RANKING order="11" place="11" resultid="101016" />
                    <RANKING order="12" place="12" resultid="101740" />
                    <RANKING order="13" place="-1" resultid="103156" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99777" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102557" />
                    <RANKING order="2" place="2" resultid="101678" />
                    <RANKING order="3" place="3" resultid="102973" />
                    <RANKING order="4" place="4" resultid="100369" />
                    <RANKING order="5" place="5" resultid="102140" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99778" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102746" />
                    <RANKING order="2" place="2" resultid="100404" />
                    <RANKING order="3" place="3" resultid="101584" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99779" agemax="84" agemin="80" name="KAT.L, 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102706" />
                    <RANKING order="2" place="2" resultid="100995" />
                    <RANKING order="3" place="3" resultid="104989" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99780" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99781" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105179" daytime="09:17" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105180" daytime="09:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105181" daytime="09:23" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105182" daytime="09:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="105183" daytime="09:28" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="105184" daytime="09:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="105185" daytime="09:32" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="105186" daytime="09:34" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="105187" daytime="09:36" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="105188" daytime="09:39" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="105189" daytime="09:41" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="105190" daytime="09:43" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="98940" daytime="09:45" gender="F" number="10" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99782" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102998" />
                    <RANKING order="2" place="2" resultid="103060" />
                    <RANKING order="3" place="3" resultid="100908" />
                    <RANKING order="4" place="4" resultid="102107" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99783" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103560" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99784" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103532" />
                    <RANKING order="2" place="2" resultid="103355" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99785" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100166" />
                    <RANKING order="2" place="2" resultid="101242" />
                    <RANKING order="3" place="3" resultid="100184" />
                    <RANKING order="4" place="4" resultid="102093" />
                    <RANKING order="5" place="5" resultid="100880" />
                    <RANKING order="6" place="6" resultid="102797" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99786" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100701" />
                    <RANKING order="2" place="2" resultid="101800" />
                    <RANKING order="3" place="-1" resultid="100114" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99787" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100816" />
                    <RANKING order="2" place="2" resultid="103495" />
                    <RANKING order="3" place="3" resultid="100873" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99788" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101745" />
                    <RANKING order="2" place="2" resultid="101459" />
                    <RANKING order="3" place="3" resultid="103114" />
                    <RANKING order="4" place="4" resultid="103463" />
                    <RANKING order="5" place="5" resultid="100426" />
                    <RANKING order="6" place="-1" resultid="101327" />
                    <RANKING order="7" place="-1" resultid="102549" />
                    <RANKING order="8" place="-1" resultid="102756" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99789" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103413" />
                    <RANKING order="2" place="2" resultid="102543" />
                    <RANKING order="3" place="3" resultid="103083" />
                    <RANKING order="4" place="4" resultid="105062" />
                    <RANKING order="5" place="5" resultid="102790" />
                    <RANKING order="6" place="6" resultid="102780" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99790" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102712" />
                    <RANKING order="2" place="2" resultid="101435" />
                    <RANKING order="3" place="-1" resultid="100446" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99791" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101453" />
                    <RANKING order="2" place="2" resultid="103383" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99792" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100711" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99793" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="105026" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99794" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99795" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99796" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105191" daytime="09:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105192" daytime="09:53" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105193" daytime="09:59" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105194" daytime="10:05" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="98956" daytime="10:15" gender="M" number="11" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99797" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102902" />
                    <RANKING order="2" place="2" resultid="104383" />
                    <RANKING order="3" place="3" resultid="104956" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99798" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100159" />
                    <RANKING order="2" place="2" resultid="103438" />
                    <RANKING order="3" place="3" resultid="101761" />
                    <RANKING order="4" place="4" resultid="101172" />
                    <RANKING order="5" place="5" resultid="101822" />
                    <RANKING order="6" place="-1" resultid="100286" />
                    <RANKING order="7" place="-1" resultid="100300" />
                    <RANKING order="8" place="-1" resultid="103009" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99799" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103538" />
                    <RANKING order="2" place="2" resultid="101730" />
                    <RANKING order="3" place="3" resultid="102376" />
                    <RANKING order="4" place="4" resultid="100325" />
                    <RANKING order="5" place="5" resultid="100153" />
                    <RANKING order="6" place="-1" resultid="101041" />
                    <RANKING order="7" place="-1" resultid="102183" />
                    <RANKING order="8" place="-1" resultid="103600" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99800" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102072" />
                    <RANKING order="2" place="2" resultid="102155" />
                    <RANKING order="3" place="3" resultid="100596" />
                    <RANKING order="4" place="4" resultid="100833" />
                    <RANKING order="5" place="5" resultid="101921" />
                    <RANKING order="6" place="6" resultid="101265" />
                    <RANKING order="7" place="7" resultid="101987" />
                    <RANKING order="8" place="-1" resultid="103050" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99801" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101235" />
                    <RANKING order="2" place="2" resultid="101213" />
                    <RANKING order="3" place="3" resultid="100189" />
                    <RANKING order="4" place="4" resultid="102040" />
                    <RANKING order="5" place="5" resultid="100242" />
                    <RANKING order="6" place="6" resultid="100984" />
                    <RANKING order="7" place="7" resultid="100780" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99802" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="105001" />
                    <RANKING order="2" place="2" resultid="101751" />
                    <RANKING order="3" place="3" resultid="101419" />
                    <RANKING order="4" place="4" resultid="100396" />
                    <RANKING order="5" place="5" resultid="105080" />
                    <RANKING order="6" place="6" resultid="103072" />
                    <RANKING order="7" place="7" resultid="101639" />
                    <RANKING order="8" place="8" resultid="100859" />
                    <RANKING order="9" place="9" resultid="101780" />
                    <RANKING order="10" place="10" resultid="102846" />
                    <RANKING order="11" place="-1" resultid="102574" />
                    <RANKING order="12" place="-1" resultid="103229" />
                    <RANKING order="13" place="-1" resultid="103617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99803" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101609" />
                    <RANKING order="2" place="2" resultid="102362" />
                    <RANKING order="3" place="3" resultid="101633" />
                    <RANKING order="4" place="4" resultid="103017" />
                    <RANKING order="5" place="5" resultid="103206" />
                    <RANKING order="6" place="6" resultid="102394" />
                    <RANKING order="7" place="-1" resultid="101659" />
                    <RANKING order="8" place="-1" resultid="103224" />
                    <RANKING order="9" place="-1" resultid="103323" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99804" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102265" />
                    <RANKING order="2" place="2" resultid="100556" />
                    <RANKING order="3" place="3" resultid="103189" />
                    <RANKING order="4" place="4" resultid="102035" />
                    <RANKING order="5" place="5" resultid="102013" />
                    <RANKING order="6" place="6" resultid="100601" />
                    <RANKING order="7" place="7" resultid="101160" />
                    <RANKING order="8" place="8" resultid="102046" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99805" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102505" />
                    <RANKING order="2" place="2" resultid="102202" />
                    <RANKING order="3" place="3" resultid="105009" />
                    <RANKING order="4" place="4" resultid="103035" />
                    <RANKING order="5" place="5" resultid="102122" />
                    <RANKING order="6" place="6" resultid="102022" />
                    <RANKING order="7" place="7" resultid="100387" />
                    <RANKING order="8" place="8" resultid="102636" />
                    <RANKING order="9" place="9" resultid="103586" />
                    <RANKING order="10" place="10" resultid="102115" />
                    <RANKING order="11" place="11" resultid="100892" />
                    <RANKING order="12" place="-1" resultid="102735" />
                    <RANKING order="13" place="-1" resultid="103172" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99806" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100565" />
                    <RANKING order="2" place="2" resultid="100351" />
                    <RANKING order="3" place="3" resultid="100772" />
                    <RANKING order="4" place="4" resultid="102129" />
                    <RANKING order="5" place="-1" resultid="103157" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99807" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100706" />
                    <RANKING order="2" place="2" resultid="100136" />
                    <RANKING order="3" place="-1" resultid="102519" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99808" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101585" />
                    <RANKING order="2" place="-1" resultid="102747" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99809" agemax="84" agemin="80" name="KAT.L, 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="102707" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99810" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99811" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105196" daytime="10:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105197" daytime="10:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105198" daytime="10:27" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105199" daytime="10:32" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="105200" daytime="10:38" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="105201" daytime="10:43" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="105202" daytime="10:47" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="105203" daytime="10:52" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="105204" daytime="10:56" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="98972" daytime="11:01" gender="F" number="12" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99812" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103471" />
                    <RANKING order="2" place="2" resultid="102999" />
                    <RANKING order="3" place="3" resultid="103610" />
                    <RANKING order="4" place="4" resultid="104378" />
                    <RANKING order="5" place="5" resultid="105069" />
                    <RANKING order="6" place="-1" resultid="100193" />
                    <RANKING order="7" place="-1" resultid="101720" />
                    <RANKING order="8" place="-1" resultid="102108" />
                    <RANKING order="9" place="-1" resultid="102415" />
                    <RANKING order="10" place="-1" resultid="103477" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99813" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103143" />
                    <RANKING order="2" place="2" resultid="101140" />
                    <RANKING order="3" place="3" resultid="102286" />
                    <RANKING order="4" place="4" resultid="103005" />
                    <RANKING order="5" place="5" resultid="101592" />
                    <RANKING order="6" place="6" resultid="102498" />
                    <RANKING order="7" place="7" resultid="101167" />
                    <RANKING order="8" place="8" resultid="101624" />
                    <RANKING order="9" place="9" resultid="101788" />
                    <RANKING order="10" place="10" resultid="100433" />
                    <RANKING order="11" place="-1" resultid="103055" />
                    <RANKING order="12" place="-1" resultid="101225" />
                    <RANKING order="13" place="-1" resultid="101347" />
                    <RANKING order="14" place="-1" resultid="102390" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99814" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101708" />
                    <RANKING order="2" place="2" resultid="102291" />
                    <RANKING order="3" place="3" resultid="101850" />
                    <RANKING order="4" place="-1" resultid="100582" />
                    <RANKING order="5" place="-1" resultid="102957" />
                    <RANKING order="6" place="-1" resultid="103524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99815" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100924" />
                    <RANKING order="2" place="2" resultid="100179" />
                    <RANKING order="3" place="3" resultid="105050" />
                    <RANKING order="4" place="4" resultid="101704" />
                    <RANKING order="5" place="5" resultid="100174" />
                    <RANKING order="6" place="6" resultid="101687" />
                    <RANKING order="7" place="-1" resultid="100881" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99816" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103332" />
                    <RANKING order="2" place="2" resultid="101357" />
                    <RANKING order="3" place="3" resultid="103132" />
                    <RANKING order="4" place="4" resultid="103126" />
                    <RANKING order="5" place="5" resultid="102898" />
                    <RANKING order="6" place="6" resultid="100115" />
                    <RANKING order="7" place="-1" resultid="100235" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99817" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103120" />
                    <RANKING order="2" place="2" resultid="105015" />
                    <RANKING order="3" place="3" resultid="103349" />
                    <RANKING order="4" place="4" resultid="103496" />
                    <RANKING order="5" place="5" resultid="101073" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99818" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101271" />
                    <RANKING order="2" place="2" resultid="100630" />
                    <RANKING order="3" place="3" resultid="103095" />
                    <RANKING order="4" place="4" resultid="102729" />
                    <RANKING order="5" place="5" resultid="103464" />
                    <RANKING order="6" place="-1" resultid="100542" />
                    <RANKING order="7" place="-1" resultid="100589" />
                    <RANKING order="8" place="-1" resultid="102836" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99819" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103089" />
                    <RANKING order="2" place="2" resultid="103338" />
                    <RANKING order="3" place="3" resultid="105022" />
                    <RANKING order="4" place="4" resultid="102720" />
                    <RANKING order="5" place="5" resultid="100936" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99820" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102535" />
                    <RANKING order="2" place="2" resultid="102713" />
                    <RANKING order="3" place="3" resultid="100953" />
                    <RANKING order="4" place="4" resultid="100670" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99821" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101495" />
                    <RANKING order="2" place="2" resultid="101569" />
                    <RANKING order="3" place="3" resultid="101841" />
                    <RANKING order="4" place="4" resultid="103384" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99822" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100687" />
                    <RANKING order="2" place="-1" resultid="102742" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99823" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103078" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99824" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99825" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99826" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105205" daytime="11:01" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105206" daytime="11:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105207" daytime="11:08" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105208" daytime="11:11" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="105209" daytime="11:14" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="105210" daytime="11:17" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="105211" daytime="11:20" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="105212" daytime="11:23" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="98988" daytime="11:26" gender="M" number="13" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99827" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100900" />
                    <RANKING order="2" place="2" resultid="103043" />
                    <RANKING order="3" place="3" resultid="102903" />
                    <RANKING order="4" place="4" resultid="102419" />
                    <RANKING order="5" place="5" resultid="103029" />
                    <RANKING order="6" place="-1" resultid="101046" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99828" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102278" />
                    <RANKING order="2" place="2" resultid="101151" />
                    <RANKING order="3" place="3" resultid="104370" />
                    <RANKING order="4" place="4" resultid="101726" />
                    <RANKING order="5" place="5" resultid="101857" />
                    <RANKING order="6" place="6" resultid="103367" />
                    <RANKING order="7" place="7" resultid="100297" />
                    <RANKING order="8" place="8" resultid="100318" />
                    <RANKING order="9" place="9" resultid="101823" />
                    <RANKING order="10" place="10" resultid="100664" />
                    <RANKING order="11" place="11" resultid="101103" />
                    <RANKING order="12" place="12" resultid="101319" />
                    <RANKING order="13" place="-1" resultid="101208" />
                    <RANKING order="14" place="-1" resultid="101229" />
                    <RANKING order="15" place="-1" resultid="102865" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99829" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102064" />
                    <RANKING order="2" place="2" resultid="100279" />
                    <RANKING order="3" place="3" resultid="100867" />
                    <RANKING order="4" place="4" resultid="102989" />
                    <RANKING order="5" place="5" resultid="103318" />
                    <RANKING order="6" place="6" resultid="102892" />
                    <RANKING order="7" place="7" resultid="101051" />
                    <RANKING order="8" place="8" resultid="102377" />
                    <RANKING order="9" place="9" resultid="101652" />
                    <RANKING order="10" place="10" resultid="101251" />
                    <RANKING order="11" place="11" resultid="101793" />
                    <RANKING order="12" place="12" resultid="102213" />
                    <RANKING order="13" place="13" resultid="100306" />
                    <RANKING order="14" place="14" resultid="101806" />
                    <RANKING order="15" place="-1" resultid="101221" />
                    <RANKING order="16" place="-1" resultid="102369" />
                    <RANKING order="17" place="-1" resultid="104373" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99830" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102156" />
                    <RANKING order="2" place="2" resultid="100754" />
                    <RANKING order="3" place="3" resultid="101810" />
                    <RANKING order="4" place="4" resultid="101133" />
                    <RANKING order="5" place="5" resultid="102581" />
                    <RANKING order="6" place="6" resultid="102100" />
                    <RANKING order="7" place="7" resultid="100292" />
                    <RANKING order="8" place="8" resultid="101599" />
                    <RANKING order="9" place="9" resultid="102478" />
                    <RANKING order="10" place="10" resultid="103447" />
                    <RANKING order="11" place="11" resultid="102492" />
                    <RANKING order="12" place="12" resultid="100107" />
                    <RANKING order="13" place="13" resultid="105390" />
                    <RANKING order="14" place="14" resultid="102248" />
                    <RANKING order="15" place="15" resultid="102254" />
                    <RANKING order="16" place="-1" resultid="100220" />
                    <RANKING order="17" place="-1" resultid="102007" />
                    <RANKING order="18" place="-1" resultid="102914" />
                    <RANKING order="19" place="-1" resultid="102964" />
                    <RANKING order="20" place="-1" resultid="103257" />
                    <RANKING order="21" place="-1" resultid="103263" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99831" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101403" />
                    <RANKING order="2" place="2" resultid="101352" />
                    <RANKING order="3" place="3" resultid="103252" />
                    <RANKING order="4" place="4" resultid="103512" />
                    <RANKING order="5" place="5" resultid="101214" />
                    <RANKING order="6" place="6" resultid="101409" />
                    <RANKING order="7" place="7" resultid="101189" />
                    <RANKING order="8" place="8" resultid="101180" />
                    <RANKING order="9" place="9" resultid="100213" />
                    <RANKING order="10" place="10" resultid="101106" />
                    <RANKING order="11" place="11" resultid="105035" />
                    <RANKING order="12" place="12" resultid="101099" />
                    <RANKING order="13" place="13" resultid="103591" />
                    <RANKING order="14" place="14" resultid="100243" />
                    <RANKING order="15" place="15" resultid="102512" />
                    <RANKING order="16" place="16" resultid="100200" />
                    <RANKING order="17" place="17" resultid="100781" />
                    <RANKING order="18" place="18" resultid="101096" />
                    <RANKING order="19" place="19" resultid="101756" />
                    <RANKING order="20" place="20" resultid="103583" />
                    <RANKING order="21" place="21" resultid="100976" />
                    <RANKING order="22" place="22" resultid="102272" />
                    <RANKING order="23" place="-1" resultid="101341" />
                    <RANKING order="24" place="-1" resultid="102983" />
                    <RANKING order="25" place="-1" resultid="101943" />
                    <RANKING order="26" place="-1" resultid="105076" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99832" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="104974" />
                    <RANKING order="2" place="2" resultid="105002" />
                    <RANKING order="3" place="3" resultid="101752" />
                    <RANKING order="4" place="4" resultid="100478" />
                    <RANKING order="5" place="5" resultid="104967" />
                    <RANKING order="6" place="6" resultid="101560" />
                    <RANKING order="7" place="7" resultid="103247" />
                    <RANKING order="8" place="8" resultid="103235" />
                    <RANKING order="9" place="9" resultid="100825" />
                    <RANKING order="10" place="10" resultid="103576" />
                    <RANKING order="11" place="11" resultid="102357" />
                    <RANKING order="12" place="12" resultid="105081" />
                    <RANKING order="13" place="13" resultid="101259" />
                    <RANKING order="14" place="14" resultid="101424" />
                    <RANKING order="15" place="15" resultid="101640" />
                    <RANKING order="16" place="16" resultid="101081" />
                    <RANKING order="17" place="-1" resultid="101699" />
                    <RANKING order="18" place="-1" resultid="102001" />
                    <RANKING order="19" place="-1" resultid="103242" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99833" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101610" />
                    <RANKING order="2" place="2" resultid="102384" />
                    <RANKING order="3" place="3" resultid="102857" />
                    <RANKING order="4" place="4" resultid="100129" />
                    <RANKING order="5" place="5" resultid="105045" />
                    <RANKING order="6" place="6" resultid="103213" />
                    <RANKING order="7" place="7" resultid="101634" />
                    <RANKING order="8" place="8" resultid="100789" />
                    <RANKING order="9" place="9" resultid="103544" />
                    <RANKING order="10" place="10" resultid="103219" />
                    <RANKING order="11" place="11" resultid="101736" />
                    <RANKING order="12" place="-1" resultid="103324" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99834" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103505" />
                    <RANKING order="2" place="2" resultid="102829" />
                    <RANKING order="3" place="3" resultid="100623" />
                    <RANKING order="4" place="4" resultid="100990" />
                    <RANKING order="5" place="5" resultid="103606" />
                    <RANKING order="6" place="6" resultid="102260" />
                    <RANKING order="7" place="7" resultid="101669" />
                    <RANKING order="8" place="8" resultid="103195" />
                    <RANKING order="9" place="-1" resultid="100929" />
                    <RANKING order="10" place="-1" resultid="100944" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99835" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101578" />
                    <RANKING order="2" place="2" resultid="101323" />
                    <RANKING order="3" place="3" resultid="100272" />
                    <RANKING order="4" place="4" resultid="102195" />
                    <RANKING order="5" place="5" resultid="101773" />
                    <RANKING order="6" place="6" resultid="101447" />
                    <RANKING order="7" place="7" resultid="101030" />
                    <RANKING order="8" place="8" resultid="103183" />
                    <RANKING order="9" place="9" resultid="103177" />
                    <RANKING order="10" place="10" resultid="102637" />
                    <RANKING order="11" place="-1" resultid="100379" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99836" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102527" />
                    <RANKING order="2" place="2" resultid="100696" />
                    <RANKING order="3" place="3" resultid="100574" />
                    <RANKING order="4" place="4" resultid="103164" />
                    <RANKING order="5" place="5" resultid="101487" />
                    <RANKING order="6" place="6" resultid="103374" />
                    <RANKING order="7" place="7" resultid="100086" />
                    <RANKING order="8" place="8" resultid="101280" />
                    <RANKING order="9" place="9" resultid="101741" />
                    <RANKING order="10" place="10" resultid="103550" />
                    <RANKING order="11" place="-1" resultid="103150" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99837" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101679" />
                    <RANKING order="2" place="2" resultid="102558" />
                    <RANKING order="3" place="3" resultid="102976" />
                    <RANKING order="4" place="4" resultid="102141" />
                    <RANKING order="5" place="5" resultid="103409" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99838" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100405" />
                    <RANKING order="2" place="2" resultid="100980" />
                    <RANKING order="3" place="-1" resultid="102135" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99839" agemax="84" agemin="80" name="KAT.L, 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100996" />
                    <RANKING order="2" place="2" resultid="104993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99840" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99841" agemax="94" agemin="90" name="KAT.N, 90-94 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100616" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105213" daytime="11:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105214" daytime="11:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105215" daytime="11:33" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105216" daytime="11:36" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="105217" daytime="11:39" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="105218" daytime="11:42" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="105219" daytime="11:44" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="105220" daytime="11:47" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="105221" daytime="11:50" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="105222" daytime="11:52" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="105223" daytime="11:55" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="105224" daytime="11:57" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="105225" daytime="12:00" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="105226" daytime="12:02" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="105227" daytime="12:05" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="105228" daytime="12:07" number="16" order="16" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99004" daytime="12:10" gender="F" number="14" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99005" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100194" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99006" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103561" />
                    <RANKING order="2" place="2" resultid="102174" />
                    <RANKING order="3" place="3" resultid="101625" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99007" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103525" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99008" agemax="39" agemin="35" name="KAT.C, 35-39 lat" />
                <AGEGROUP agegroupid="99009" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100610" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99010" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100817" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99011" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100438" />
                    <RANKING order="2" place="-1" resultid="102757" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99012" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101993" />
                    <RANKING order="2" place="-1" resultid="102700" />
                    <RANKING order="3" place="-1" resultid="102721" />
                    <RANKING order="4" place="-1" resultid="102781" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99013" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101436" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99014" agemax="69" agemin="65" name="KAT.I, 65-69 lat" />
                <AGEGROUP agegroupid="99015" agemax="74" agemin="70" name="KAT.J, 70-74 lat" />
                <AGEGROUP agegroupid="99016" agemax="79" agemin="75" name="KAT.K, 75-79 lat" />
                <AGEGROUP agegroupid="99017" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99018" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99019" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105229" daytime="12:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105230" daytime="12:17" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99020" daytime="12:23" gender="M" number="15" order="8" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99021" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="104957" />
                    <RANKING order="2" place="2" resultid="100799" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99022" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100287" />
                    <RANKING order="2" place="-1" resultid="100319" />
                    <RANKING order="3" place="-1" resultid="103010" />
                    <RANKING order="4" place="-1" resultid="103023" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99023" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102990" />
                    <RANKING order="2" place="2" resultid="102147" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99024" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101922" />
                    <RANKING order="2" place="2" resultid="102165" />
                    <RANKING order="3" place="3" resultid="101714" />
                    <RANKING order="4" place="4" resultid="104401" />
                    <RANKING order="5" place="5" resultid="100808" />
                    <RANKING order="6" place="-1" resultid="102965" />
                    <RANKING order="7" place="-1" resultid="100221" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99025" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100763" />
                    <RANKING order="2" place="2" resultid="103397" />
                    <RANKING order="3" place="3" resultid="100471" />
                    <RANKING order="4" place="-1" resultid="101936" />
                    <RANKING order="5" place="-1" resultid="101093" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99026" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101832" />
                    <RANKING order="2" place="2" resultid="100453" />
                    <RANKING order="3" place="3" resultid="101466" />
                    <RANKING order="4" place="4" resultid="103568" />
                    <RANKING order="5" place="5" resultid="100917" />
                    <RANKING order="6" place="-1" resultid="101781" />
                    <RANKING order="7" place="-1" resultid="102841" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99027" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103199" />
                    <RANKING order="2" place="2" resultid="101443" />
                    <RANKING order="3" place="3" resultid="104979" />
                    <RANKING order="4" place="4" resultid="100790" />
                    <RANKING order="5" place="5" resultid="102350" />
                    <RANKING order="6" place="6" resultid="102395" />
                    <RANKING order="7" place="-1" resultid="100121" />
                    <RANKING order="8" place="-1" resultid="101660" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99028" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100557" />
                    <RANKING order="2" place="2" resultid="102014" />
                    <RANKING order="3" place="3" resultid="102029" />
                    <RANKING order="4" place="4" resultid="101089" />
                    <RANKING order="5" place="-1" resultid="100602" />
                    <RANKING order="6" place="-1" resultid="100945" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99029" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102023" />
                    <RANKING order="2" place="2" resultid="105096" />
                    <RANKING order="3" place="3" resultid="101060" />
                    <RANKING order="4" place="4" resultid="100388" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99030" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100352" />
                    <RANKING order="2" place="2" resultid="101289" />
                    <RANKING order="3" place="3" resultid="105056" />
                    <RANKING order="4" place="4" resultid="102949" />
                    <RANKING order="5" place="5" resultid="101017" />
                    <RANKING order="6" place="-1" resultid="100575" />
                    <RANKING order="7" place="-1" resultid="103375" />
                    <RANKING order="8" place="-1" resultid="102969" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99031" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100137" />
                    <RANKING order="2" place="2" resultid="100370" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99032" agemax="79" agemin="75" name="KAT.K, 75-79 lat" />
                <AGEGROUP agegroupid="99033" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99034" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99035" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105231" daytime="12:23" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105232" daytime="12:29" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105233" daytime="12:36" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105234" daytime="12:42" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="105235" daytime="12:47" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="105236" daytime="12:51" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99036" daytime="12:56" gender="F" number="16" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99512" agemax="96" agemin="80" name="KAT.0, 80-96 lat" calculate="TOTAL" />
                <AGEGROUP agegroupid="99513" agemax="119" agemin="100" name="KAT.A, 100-119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101871" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99514" agemax="159" agemin="120" name="KAT.B, 120-159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101870" />
                    <RANKING order="2" place="2" resultid="104099" />
                    <RANKING order="3" place="3" resultid="100252" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99515" agemax="199" agemin="160" name="KAT.C,160-199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103270" />
                    <RANKING order="2" place="2" resultid="100638" />
                    <RANKING order="3" place="-1" resultid="101371" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99516" agemax="239" agemin="200" name="KAT.D, 200-239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103422" />
                    <RANKING order="2" place="2" resultid="103272" />
                    <RANKING order="3" place="3" resultid="101373" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99517" agemax="279" agemin="240" name="KAT.E, 240-279 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100732" />
                    <RANKING order="2" place="2" resultid="102762" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99518" agemax="-1" agemin="280" name="KAT.F, 280+ lat" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105237" daytime="12:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105238" daytime="13:31" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99059" daytime="13:36" gender="M" number="17" order="10" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99519" agemax="96" agemin="80" name="KAT.0, 80-96 lat" calculate="TOTAL" />
                <AGEGROUP agegroupid="99520" agemax="119" agemin="100" name="KAT.A, 100-119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101872" />
                    <RANKING order="2" place="2" resultid="103480" />
                    <RANKING order="3" place="3" resultid="100329" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99521" agemax="159" agemin="120" name="KAT.B, 120-159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101874" />
                    <RANKING order="2" place="2" resultid="100254" />
                    <RANKING order="3" place="3" resultid="103431" />
                    <RANKING order="4" place="4" resultid="100331" />
                    <RANKING order="5" place="5" resultid="104101" />
                    <RANKING order="6" place="6" resultid="101367" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99522" agemax="199" agemin="160" name="KAT.C,160-199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100837" />
                    <RANKING order="2" place="2" resultid="101873" />
                    <RANKING order="3" place="3" resultid="105085" />
                    <RANKING order="4" place="4" resultid="102220" />
                    <RANKING order="5" place="5" resultid="104100" />
                    <RANKING order="6" place="6" resultid="102295" />
                    <RANKING order="7" place="7" resultid="103278" />
                    <RANKING order="8" place="8" resultid="100255" />
                    <RANKING order="9" place="9" resultid="101111" />
                    <RANKING order="10" place="10" resultid="102869" />
                    <RANKING order="11" place="11" resultid="102222" />
                    <RANKING order="12" place="12" resultid="103425" />
                    <RANKING order="13" place="13" resultid="104102" />
                    <RANKING order="14" place="14" resultid="101113" />
                    <RANKING order="15" place="-1" resultid="101947" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99523" agemax="239" agemin="200" name="KAT.D, 200-239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103275" />
                    <RANKING order="2" place="2" resultid="102398" />
                    <RANKING order="3" place="-1" resultid="101369" />
                    <RANKING order="4" place="-1" resultid="101882" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99524" agemax="279" agemin="240" name="KAT.E, 240-279 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100640" />
                    <RANKING order="2" place="2" resultid="103273" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99525" agemax="-1" agemin="280" name="KAT.F, 280+ lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100733" />
                    <RANKING order="2" place="2" resultid="102765" />
                    <RANKING order="3" place="3" resultid="102218" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105239" daytime="13:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105240" daytime="13:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105241" daytime="13:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105242" daytime="13:49" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2014-06-28" daytime="16:00" number="3" warmupfrom="15:00">
          <EVENTS>
            <EVENT eventid="99089" daytime="16:00" gender="F" number="18" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99109" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103000" />
                    <RANKING order="2" place="2" resultid="100909" />
                    <RANKING order="3" place="3" resultid="103061" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99110" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102499" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99111" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103533" />
                    <RANKING order="2" place="2" resultid="103356" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99112" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100167" />
                    <RANKING order="2" place="2" resultid="101243" />
                    <RANKING order="3" place="3" resultid="100185" />
                    <RANKING order="4" place="4" resultid="102094" />
                    <RANKING order="5" place="5" resultid="100882" />
                    <RANKING order="6" place="-1" resultid="102798" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99113" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100702" />
                    <RANKING order="2" place="2" resultid="101801" />
                    <RANKING order="3" place="3" resultid="100116" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99114" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103350" />
                    <RANKING order="2" place="2" resultid="101074" />
                    <RANKING order="3" place="3" resultid="100818" />
                    <RANKING order="4" place="4" resultid="100874" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99115" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100631" />
                    <RANKING order="2" place="2" resultid="101746" />
                    <RANKING order="3" place="3" resultid="101460" />
                    <RANKING order="4" place="4" resultid="103465" />
                    <RANKING order="5" place="5" resultid="100427" />
                    <RANKING order="6" place="-1" resultid="101328" />
                    <RANKING order="7" place="-1" resultid="102550" />
                    <RANKING order="8" place="-1" resultid="103115" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99116" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103414" />
                    <RANKING order="2" place="2" resultid="102544" />
                    <RANKING order="3" place="3" resultid="103084" />
                    <RANKING order="4" place="4" resultid="102722" />
                    <RANKING order="5" place="5" resultid="105063" />
                    <RANKING order="6" place="6" resultid="102791" />
                    <RANKING order="7" place="7" resultid="102782" />
                    <RANKING order="8" place="-1" resultid="101297" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99117" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102714" />
                    <RANKING order="2" place="2" resultid="100447" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99118" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101454" />
                    <RANKING order="2" place="2" resultid="101285" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99119" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100712" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99120" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="105027" />
                    <RANKING order="2" place="2" resultid="103079" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99121" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99122" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99123" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105243" daytime="16:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105244" daytime="16:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105245" daytime="16:07" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105246" daytime="16:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="105247" daytime="16:12" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99091" daytime="16:15" gender="M" number="19" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99124" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102904" />
                    <RANKING order="2" place="2" resultid="104958" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99125" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="105109" />
                    <RANKING order="2" place="2" resultid="100160" />
                    <RANKING order="3" place="3" resultid="101762" />
                    <RANKING order="4" place="4" resultid="103439" />
                    <RANKING order="5" place="5" resultid="101173" />
                    <RANKING order="6" place="6" resultid="101824" />
                    <RANKING order="7" place="7" resultid="100301" />
                    <RANKING order="8" place="-1" resultid="101301" />
                    <RANKING order="9" place="-1" resultid="103011" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99126" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103453" />
                    <RANKING order="2" place="2" resultid="101731" />
                    <RANKING order="3" place="3" resultid="100326" />
                    <RANKING order="4" place="4" resultid="100154" />
                    <RANKING order="5" place="5" resultid="101250" />
                    <RANKING order="6" place="6" resultid="102214" />
                    <RANKING order="7" place="-1" resultid="103539" />
                    <RANKING order="8" place="-1" resultid="100307" />
                    <RANKING order="9" place="-1" resultid="101042" />
                    <RANKING order="10" place="-1" resultid="102991" />
                    <RANKING order="11" place="-1" resultid="103601" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99127" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102073" />
                    <RANKING order="2" place="2" resultid="102157" />
                    <RANKING order="3" place="3" resultid="100834" />
                    <RANKING order="4" place="4" resultid="100597" />
                    <RANKING order="5" place="5" resultid="101266" />
                    <RANKING order="6" place="6" resultid="102582" />
                    <RANKING order="7" place="7" resultid="101600" />
                    <RANKING order="8" place="8" resultid="100809" />
                    <RANKING order="9" place="9" resultid="100413" />
                    <RANKING order="10" place="10" resultid="101816" />
                    <RANKING order="11" place="11" resultid="102493" />
                    <RANKING order="12" place="-1" resultid="102915" />
                    <RANKING order="13" place="-1" resultid="103258" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99128" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101404" />
                    <RANKING order="2" place="2" resultid="100764" />
                    <RANKING order="3" place="3" resultid="101236" />
                    <RANKING order="4" place="4" resultid="100190" />
                    <RANKING order="5" place="5" resultid="101110" />
                    <RANKING order="6" place="6" resultid="100244" />
                    <RANKING order="7" place="7" resultid="102041" />
                    <RANKING order="8" place="8" resultid="100985" />
                    <RANKING order="9" place="-1" resultid="100655" />
                    <RANKING order="10" place="-1" resultid="100960" />
                    <RANKING order="11" place="-1" resultid="101204" />
                    <RANKING order="12" place="-1" resultid="101215" />
                    <RANKING order="13" place="-1" resultid="101931" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99129" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101753" />
                    <RANKING order="2" place="2" resultid="101038" />
                    <RANKING order="3" place="3" resultid="101420" />
                    <RANKING order="4" place="4" resultid="103616" />
                    <RANKING order="5" place="5" resultid="102575" />
                    <RANKING order="6" place="6" resultid="101561" />
                    <RANKING order="7" place="7" resultid="100397" />
                    <RANKING order="8" place="8" resultid="101641" />
                    <RANKING order="9" place="9" resultid="100860" />
                    <RANKING order="10" place="10" resultid="101782" />
                    <RANKING order="11" place="11" resultid="100467" />
                    <RANKING order="12" place="-1" resultid="101332" />
                    <RANKING order="13" place="-1" resultid="102002" />
                    <RANKING order="14" place="-1" resultid="102847" />
                    <RANKING order="15" place="-1" resultid="103073" />
                    <RANKING order="16" place="-1" resultid="103230" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99130" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101611" />
                    <RANKING order="2" place="2" resultid="101635" />
                    <RANKING order="3" place="3" resultid="101480" />
                    <RANKING order="4" place="4" resultid="102363" />
                    <RANKING order="5" place="5" resultid="103207" />
                    <RANKING order="6" place="6" resultid="103325" />
                    <RANKING order="7" place="-1" resultid="103225" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99131" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102266" />
                    <RANKING order="2" place="2" resultid="100558" />
                    <RANKING order="3" place="3" resultid="103190" />
                    <RANKING order="4" place="4" resultid="100603" />
                    <RANKING order="5" place="5" resultid="102036" />
                    <RANKING order="6" place="6" resultid="102047" />
                    <RANKING order="7" place="7" resultid="103362" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99132" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102506" />
                    <RANKING order="2" place="2" resultid="102203" />
                    <RANKING order="3" place="3" resultid="105010" />
                    <RANKING order="4" place="4" resultid="103036" />
                    <RANKING order="5" place="5" resultid="102123" />
                    <RANKING order="6" place="6" resultid="102638" />
                    <RANKING order="7" place="7" resultid="102736" />
                    <RANKING order="8" place="8" resultid="103587" />
                    <RANKING order="9" place="9" resultid="100389" />
                    <RANKING order="10" place="10" resultid="102116" />
                    <RANKING order="11" place="11" resultid="100893" />
                    <RANKING order="12" place="-1" resultid="101275" />
                    <RANKING order="13" place="-1" resultid="101324" />
                    <RANKING order="14" place="-1" resultid="103173" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99133" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100566" />
                    <RANKING order="2" place="2" resultid="100570" />
                    <RANKING order="3" place="3" resultid="102130" />
                    <RANKING order="4" place="-1" resultid="103158" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99134" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100707" />
                    <RANKING order="2" place="2" resultid="100138" />
                    <RANKING order="3" place="3" resultid="102520" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99135" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102748" />
                    <RANKING order="2" place="2" resultid="102136" />
                    <RANKING order="3" place="-1" resultid="101586" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99136" agemax="84" agemin="80" name="KAT.L, 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102708" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99137" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99138" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105248" daytime="16:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105249" daytime="16:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105250" daytime="16:24" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105251" daytime="16:27" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="105252" daytime="16:30" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="105253" daytime="16:32" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="105254" daytime="16:35" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="105255" daytime="16:37" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="105256" daytime="16:40" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="105257" daytime="16:42" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="105258" daytime="16:44" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99154" daytime="16:47" gender="F" number="20" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99842" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103472" />
                    <RANKING order="2" place="2" resultid="103614" />
                    <RANKING order="3" place="3" resultid="102416" />
                    <RANKING order="4" place="4" resultid="100313" />
                    <RANKING order="5" place="5" resultid="100195" />
                    <RANKING order="6" place="6" resultid="104379" />
                    <RANKING order="7" place="-1" resultid="101721" />
                    <RANKING order="8" place="-1" resultid="103062" />
                    <RANKING order="9" place="-1" resultid="103478" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99843" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103144" />
                    <RANKING order="2" place="2" resultid="103139" />
                    <RANKING order="3" place="3" resultid="102175" />
                    <RANKING order="4" place="4" resultid="103562" />
                    <RANKING order="5" place="5" resultid="101593" />
                    <RANKING order="6" place="6" resultid="101626" />
                    <RANKING order="7" place="7" resultid="103056" />
                    <RANKING order="8" place="8" resultid="101618" />
                    <RANKING order="9" place="-1" resultid="101226" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99844" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101709" />
                    <RANKING order="2" place="2" resultid="102292" />
                    <RANKING order="3" place="3" resultid="105084" />
                    <RANKING order="4" place="4" resultid="101851" />
                    <RANKING order="5" place="5" resultid="103526" />
                    <RANKING order="6" place="-1" resultid="100583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99845" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100180" />
                    <RANKING order="2" place="2" resultid="105051" />
                    <RANKING order="3" place="3" resultid="102095" />
                    <RANKING order="4" place="-1" resultid="101306" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99846" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100611" />
                    <RANKING order="2" place="2" resultid="103333" />
                    <RANKING order="3" place="3" resultid="100967" />
                    <RANKING order="4" place="4" resultid="101802" />
                    <RANKING order="5" place="5" resultid="103133" />
                    <RANKING order="6" place="-1" resultid="102054" />
                    <RANKING order="7" place="-1" resultid="103345" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99847" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103121" />
                    <RANKING order="2" place="2" resultid="103351" />
                    <RANKING order="3" place="3" resultid="100819" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99848" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101272" />
                    <RANKING order="2" place="2" resultid="100590" />
                    <RANKING order="3" place="3" resultid="102458" />
                    <RANKING order="4" place="4" resultid="103466" />
                    <RANKING order="5" place="-1" resultid="100428" />
                    <RANKING order="6" place="-1" resultid="101310" />
                    <RANKING order="7" place="-1" resultid="102551" />
                    <RANKING order="8" place="-1" resultid="102730" />
                    <RANKING order="9" place="-1" resultid="102758" />
                    <RANKING order="10" place="-1" resultid="103101" />
                    <RANKING order="11" place="-1" resultid="103107" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99849" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103090" />
                    <RANKING order="2" place="2" resultid="102545" />
                    <RANKING order="3" place="3" resultid="102723" />
                    <RANKING order="4" place="4" resultid="103339" />
                    <RANKING order="5" place="5" resultid="102783" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99850" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102536" />
                    <RANKING order="2" place="2" resultid="102463" />
                    <RANKING order="3" place="3" resultid="100954" />
                    <RANKING order="4" place="4" resultid="101437" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99851" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103385" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99852" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100713" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99853" agemax="79" agemin="75" name="KAT.K, 75-79 lat" />
                <AGEGROUP agegroupid="99854" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99855" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99856" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105259" daytime="16:47" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105260" daytime="16:49" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105261" daytime="16:51" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105262" daytime="16:52" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="105263" daytime="16:54" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="105264" daytime="16:55" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99170" daytime="16:57" gender="M" number="21" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99857" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102411" />
                    <RANKING order="2" place="2" resultid="100901" />
                    <RANKING order="3" place="3" resultid="102420" />
                    <RANKING order="4" place="4" resultid="101047" />
                    <RANKING order="5" place="5" resultid="103030" />
                    <RANKING order="6" place="-1" resultid="102808" />
                    <RANKING order="7" place="-1" resultid="103044" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99858" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102279" />
                    <RANKING order="2" place="2" resultid="101003" />
                    <RANKING order="3" place="3" resultid="101152" />
                    <RANKING order="4" place="4" resultid="101727" />
                    <RANKING order="5" place="5" resultid="103457" />
                    <RANKING order="6" place="6" resultid="101858" />
                    <RANKING order="7" place="7" resultid="100161" />
                    <RANKING order="8" place="8" resultid="103368" />
                    <RANKING order="9" place="9" resultid="100320" />
                    <RANKING order="10" place="10" resultid="101825" />
                    <RANKING order="11" place="-1" resultid="101209" />
                    <RANKING order="12" place="-1" resultid="101320" />
                    <RANKING order="13" place="-1" resultid="101763" />
                    <RANKING order="14" place="-1" resultid="102866" />
                    <RANKING order="15" place="-1" resultid="103012" />
                    <RANKING order="16" place="-1" resultid="105106" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99859" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102065" />
                    <RANKING order="2" place="2" resultid="105112" />
                    <RANKING order="3" place="3" resultid="101768" />
                    <RANKING order="4" place="4" resultid="102893" />
                    <RANKING order="5" place="5" resultid="103319" />
                    <RANKING order="6" place="6" resultid="101052" />
                    <RANKING order="7" place="7" resultid="101653" />
                    <RANKING order="8" place="8" resultid="101807" />
                    <RANKING order="9" place="-1" resultid="101794" />
                    <RANKING order="10" place="-1" resultid="102208" />
                    <RANKING order="11" place="-1" resultid="102370" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99860" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102822" />
                    <RANKING order="2" place="2" resultid="103051" />
                    <RANKING order="3" place="3" resultid="102882" />
                    <RANKING order="4" place="4" resultid="101811" />
                    <RANKING order="5" place="5" resultid="100414" />
                    <RANKING order="6" place="6" resultid="102583" />
                    <RANKING order="7" place="7" resultid="100222" />
                    <RANKING order="8" place="8" resultid="104402" />
                    <RANKING order="9" place="9" resultid="100207" />
                    <RANKING order="10" place="10" resultid="102101" />
                    <RANKING order="11" place="11" resultid="101817" />
                    <RANKING order="12" place="12" resultid="101068" />
                    <RANKING order="13" place="13" resultid="102249" />
                    <RANKING order="14" place="14" resultid="100108" />
                    <RANKING order="15" place="15" resultid="102255" />
                    <RANKING order="16" place="-1" resultid="102189" />
                    <RANKING order="17" place="-1" resultid="102472" />
                    <RANKING order="18" place="-1" resultid="103259" />
                    <RANKING order="19" place="-1" resultid="103264" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99861" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101353" />
                    <RANKING order="2" place="2" resultid="100472" />
                    <RANKING order="3" place="3" resultid="103513" />
                    <RANKING order="4" place="4" resultid="101094" />
                    <RANKING order="5" place="5" resultid="101100" />
                    <RANKING order="6" place="6" resultid="100214" />
                    <RANKING order="7" place="7" resultid="101107" />
                    <RANKING order="8" place="8" resultid="103398" />
                    <RANKING order="9" place="9" resultid="102513" />
                    <RANKING order="10" place="10" resultid="100986" />
                    <RANKING order="11" place="11" resultid="103592" />
                    <RANKING order="12" place="12" resultid="100245" />
                    <RANKING order="13" place="13" resultid="105074" />
                    <RANKING order="14" place="14" resultid="100782" />
                    <RANKING order="15" place="15" resultid="100201" />
                    <RANKING order="16" place="16" resultid="101757" />
                    <RANKING order="17" place="-1" resultid="100656" />
                    <RANKING order="18" place="-1" resultid="101937" />
                    <RANKING order="19" place="-1" resultid="101944" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99862" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="105003" />
                    <RANKING order="2" place="2" resultid="101833" />
                    <RANKING order="3" place="3" resultid="100479" />
                    <RANKING order="4" place="4" resultid="100460" />
                    <RANKING order="5" place="5" resultid="101467" />
                    <RANKING order="6" place="6" resultid="100826" />
                    <RANKING order="7" place="7" resultid="103491" />
                    <RANKING order="8" place="8" resultid="103236" />
                    <RANKING order="9" place="9" resultid="104382" />
                    <RANKING order="10" place="10" resultid="105095" />
                    <RANKING order="11" place="11" resultid="103598" />
                    <RANKING order="12" place="12" resultid="101642" />
                    <RANKING order="13" place="13" resultid="101082" />
                    <RANKING order="14" place="-1" resultid="100861" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99863" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100130" />
                    <RANKING order="2" place="2" resultid="101500" />
                    <RANKING order="3" place="3" resultid="102858" />
                    <RANKING order="4" place="4" resultid="103220" />
                    <RANKING order="5" place="5" resultid="103214" />
                    <RANKING order="6" place="-1" resultid="100122" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99864" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102830" />
                    <RANKING order="2" place="2" resultid="102261" />
                    <RANKING order="3" place="3" resultid="100946" />
                    <RANKING order="4" place="4" resultid="100991" />
                    <RANKING order="5" place="5" resultid="102048" />
                    <RANKING order="6" place="6" resultid="101670" />
                    <RANKING order="7" place="7" resultid="101090" />
                    <RANKING order="8" place="-1" resultid="100604" />
                    <RANKING order="9" place="-1" resultid="100930" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99865" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102196" />
                    <RANKING order="2" place="2" resultid="100380" />
                    <RANKING order="3" place="3" resultid="103178" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99866" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102528" />
                    <RANKING order="2" place="2" resultid="100353" />
                    <RANKING order="3" place="3" resultid="100697" />
                    <RANKING order="4" place="4" resultid="100576" />
                    <RANKING order="5" place="5" resultid="103165" />
                    <RANKING order="6" place="6" resultid="101742" />
                    <RANKING order="7" place="7" resultid="103151" />
                    <RANKING order="8" place="8" resultid="100718" />
                    <RANKING order="9" place="9" resultid="101018" />
                    <RANKING order="10" place="-1" resultid="100087" />
                    <RANKING order="11" place="-1" resultid="101290" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99867" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100708" />
                    <RANKING order="2" place="2" resultid="100139" />
                    <RANKING order="3" place="-1" resultid="102977" />
                    <RANKING order="4" place="-1" resultid="100371" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99868" agemax="79" agemin="75" name="KAT.K, 75-79 lat" />
                <AGEGROUP agegroupid="99869" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99870" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99871" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105265" daytime="16:57" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105266" daytime="16:59" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105267" daytime="17:01" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105268" daytime="17:02" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="105269" daytime="17:04" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="105270" daytime="17:06" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="105271" daytime="17:07" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="105272" daytime="17:09" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="105273" daytime="17:10" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="105274" daytime="17:12" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="105275" daytime="17:13" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="105276" daytime="17:15" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99186" daytime="17:28" gender="M" number="23" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99887" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100972" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99888" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101004" />
                    <RANKING order="2" place="2" resultid="101146" />
                    <RANKING order="3" place="3" resultid="103443" />
                    <RANKING order="4" place="4" resultid="105091" />
                    <RANKING order="5" place="5" resultid="100298" />
                    <RANKING order="6" place="6" resultid="101646" />
                    <RANKING order="7" place="-1" resultid="102867" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99889" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102371" />
                    <RANKING order="2" place="2" resultid="102184" />
                    <RANKING order="3" place="3" resultid="101732" />
                    <RANKING order="4" place="4" resultid="102888" />
                    <RANKING order="5" place="5" resultid="102209" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99890" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102823" />
                    <RANKING order="2" place="2" resultid="100755" />
                    <RANKING order="3" place="3" resultid="102166" />
                    <RANKING order="4" place="4" resultid="101197" />
                    <RANKING order="5" place="5" resultid="103052" />
                    <RANKING order="6" place="6" resultid="102102" />
                    <RANKING order="7" place="7" resultid="103448" />
                    <RANKING order="8" place="8" resultid="104403" />
                    <RANKING order="9" place="9" resultid="101818" />
                    <RANKING order="10" place="-1" resultid="100208" />
                    <RANKING order="11" place="-1" resultid="102190" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99891" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101190" />
                    <RANKING order="2" place="2" resultid="101405" />
                    <RANKING order="3" place="3" resultid="101475" />
                    <RANKING order="4" place="4" resultid="101181" />
                    <RANKING order="5" place="5" resultid="101415" />
                    <RANKING order="6" place="6" resultid="105075" />
                    <RANKING order="7" place="7" resultid="101097" />
                    <RANKING order="8" place="-1" resultid="100961" />
                    <RANKING order="9" place="-1" resultid="101932" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99892" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100722" />
                    <RANKING order="2" place="2" resultid="104968" />
                    <RANKING order="3" place="3" resultid="101700" />
                    <RANKING order="4" place="4" resultid="102358" />
                    <RANKING order="5" place="5" resultid="100398" />
                    <RANKING order="6" place="6" resultid="100827" />
                    <RANKING order="7" place="7" resultid="100918" />
                    <RANKING order="8" place="8" resultid="103556" />
                    <RANKING order="9" place="-1" resultid="103243" />
                    <RANKING order="10" place="-1" resultid="103577" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99893" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100131" />
                    <RANKING order="2" place="2" resultid="101481" />
                    <RANKING order="3" place="3" resultid="100660" />
                    <RANKING order="4" place="4" resultid="102859" />
                    <RANKING order="5" place="5" resultid="100791" />
                    <RANKING order="6" place="6" resultid="102364" />
                    <RANKING order="7" place="-1" resultid="101661" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99894" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102831" />
                    <RANKING order="2" place="2" resultid="100624" />
                    <RANKING order="3" place="3" resultid="102570" />
                    <RANKING order="4" place="4" resultid="102037" />
                    <RANKING order="5" place="5" resultid="102030" />
                    <RANKING order="6" place="6" resultid="103363" />
                    <RANKING order="7" place="-1" resultid="100674" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99895" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101579" />
                    <RANKING order="2" place="2" resultid="101061" />
                    <RANKING order="3" place="3" resultid="103184" />
                    <RANKING order="4" place="4" resultid="101031" />
                    <RANKING order="5" place="5" resultid="100381" />
                    <RANKING order="6" place="6" resultid="102564" />
                    <RANKING order="7" place="7" resultid="100894" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99896" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100773" />
                    <RANKING order="2" place="2" resultid="101488" />
                    <RANKING order="3" place="3" resultid="100678" />
                    <RANKING order="4" place="4" resultid="101281" />
                    <RANKING order="5" place="5" resultid="102950" />
                    <RANKING order="6" place="6" resultid="103403" />
                    <RANKING order="7" place="7" resultid="101336" />
                    <RANKING order="8" place="8" resultid="102131" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99897" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102559" />
                    <RANKING order="2" place="2" resultid="101680" />
                    <RANKING order="3" place="3" resultid="102142" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99898" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102749" />
                    <RANKING order="2" place="2" resultid="100406" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99899" agemax="84" agemin="80" name="KAT.L, 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100997" />
                    <RANKING order="2" place="2" resultid="104990" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99900" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99901" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105281" daytime="17:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105282" daytime="17:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105283" daytime="17:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105284" daytime="17:37" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="105285" daytime="17:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="105286" daytime="17:42" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="105287" daytime="17:44" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="105288" daytime="17:47" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99202" daytime="17:49" gender="F" number="24" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99902" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103001" />
                    <RANKING order="2" place="2" resultid="103611" />
                    <RANKING order="3" place="3" resultid="105070" />
                    <RANKING order="4" place="-1" resultid="100196" />
                    <RANKING order="5" place="-1" resultid="101722" />
                    <RANKING order="6" place="-1" resultid="102109" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99903" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103145" />
                    <RANKING order="2" place="2" resultid="101141" />
                    <RANKING order="3" place="3" resultid="102287" />
                    <RANKING order="4" place="4" resultid="101594" />
                    <RANKING order="5" place="5" resultid="102500" />
                    <RANKING order="6" place="6" resultid="103006" />
                    <RANKING order="7" place="7" resultid="101169" />
                    <RANKING order="8" place="8" resultid="101627" />
                    <RANKING order="9" place="9" resultid="100434" />
                    <RANKING order="10" place="-1" resultid="101619" />
                    <RANKING order="11" place="-1" resultid="101348" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99904" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103534" />
                    <RANKING order="2" place="2" resultid="103527" />
                    <RANKING order="3" place="3" resultid="101852" />
                    <RANKING order="4" place="4" resultid="100585" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99905" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100925" />
                    <RANKING order="2" place="2" resultid="100181" />
                    <RANKING order="3" place="3" resultid="100175" />
                    <RANKING order="4" place="4" resultid="101689" />
                    <RANKING order="5" place="5" resultid="100883" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99906" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100968" />
                    <RANKING order="2" place="2" resultid="101358" />
                    <RANKING order="3" place="3" resultid="103134" />
                    <RANKING order="4" place="4" resultid="103334" />
                    <RANKING order="5" place="5" resultid="100237" />
                    <RANKING order="6" place="6" resultid="102899" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99907" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103122" />
                    <RANKING order="2" place="2" resultid="100551" />
                    <RANKING order="3" place="3" resultid="105016" />
                    <RANKING order="4" place="4" resultid="103497" />
                    <RANKING order="5" place="5" resultid="101076" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99908" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103096" />
                    <RANKING order="2" place="2" resultid="101449" />
                    <RANKING order="3" place="3" resultid="101747" />
                    <RANKING order="4" place="4" resultid="101462" />
                    <RANKING order="5" place="5" resultid="102731" />
                    <RANKING order="6" place="-1" resultid="100541" />
                    <RANKING order="7" place="-1" resultid="100632" />
                    <RANKING order="8" place="-1" resultid="102837" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99909" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100938" />
                    <RANKING order="2" place="2" resultid="102792" />
                    <RANKING order="3" place="-1" resultid="103340" />
                    <RANKING order="4" place="-1" resultid="105102" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99910" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102537" />
                    <RANKING order="2" place="2" resultid="102715" />
                    <RANKING order="3" place="3" resultid="100955" />
                    <RANKING order="4" place="4" resultid="101438" />
                    <RANKING order="5" place="-1" resultid="100671" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99911" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101842" />
                    <RANKING order="2" place="2" resultid="103386" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99912" agemax="74" agemin="70" name="KAT.J, 70-74 lat" />
                <AGEGROUP agegroupid="99913" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101470" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99914" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99915" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99916" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105289" daytime="17:49" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105290" daytime="17:55" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105291" daytime="17:59" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105292" daytime="18:04" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="105293" daytime="18:07" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="105294" daytime="18:11" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99218" daytime="18:14" gender="M" number="25" order="10" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99917" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102905" />
                    <RANKING order="2" place="2" resultid="100800" />
                    <RANKING order="3" place="3" resultid="100682" />
                    <RANKING order="4" place="-1" resultid="102809" />
                    <RANKING order="5" place="-1" resultid="103031" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99918" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101153" />
                    <RANKING order="2" place="2" resultid="102280" />
                    <RANKING order="3" place="3" resultid="103458" />
                    <RANKING order="4" place="4" resultid="101859" />
                    <RANKING order="5" place="5" resultid="103369" />
                    <RANKING order="6" place="6" resultid="101174" />
                    <RANKING order="7" place="-1" resultid="101230" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99919" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102066" />
                    <RANKING order="2" place="2" resultid="101010" />
                    <RANKING order="3" place="3" resultid="102378" />
                    <RANKING order="4" place="4" resultid="100280" />
                    <RANKING order="5" place="4" resultid="100868" />
                    <RANKING order="6" place="6" resultid="102894" />
                    <RANKING order="7" place="7" resultid="101053" />
                    <RANKING order="8" place="8" resultid="101654" />
                    <RANKING order="9" place="9" resultid="102992" />
                    <RANKING order="10" place="10" resultid="102148" />
                    <RANKING order="11" place="11" resultid="101808" />
                    <RANKING order="12" place="-1" resultid="101795" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99920" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102158" />
                    <RANKING order="2" place="2" resultid="102883" />
                    <RANKING order="3" place="3" resultid="101923" />
                    <RANKING order="4" place="4" resultid="101812" />
                    <RANKING order="5" place="5" resultid="100756" />
                    <RANKING order="6" place="6" resultid="101134" />
                    <RANKING order="7" place="7" resultid="102494" />
                    <RANKING order="8" place="8" resultid="101069" />
                    <RANKING order="9" place="-1" resultid="100109" />
                    <RANKING order="10" place="-1" resultid="100223" />
                    <RANKING order="11" place="-1" resultid="101601" />
                    <RANKING order="12" place="-1" resultid="102008" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99921" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101216" />
                    <RANKING order="2" place="2" resultid="103253" />
                    <RANKING order="3" place="3" resultid="103514" />
                    <RANKING order="4" place="4" resultid="101410" />
                    <RANKING order="5" place="5" resultid="101191" />
                    <RANKING order="6" place="6" resultid="105036" />
                    <RANKING order="7" place="7" resultid="100473" />
                    <RANKING order="8" place="8" resultid="100215" />
                    <RANKING order="9" place="9" resultid="103593" />
                    <RANKING order="10" place="10" resultid="102514" />
                    <RANKING order="11" place="11" resultid="100202" />
                    <RANKING order="12" place="12" resultid="101758" />
                    <RANKING order="13" place="13" resultid="101605" />
                    <RANKING order="14" place="14" resultid="103584" />
                    <RANKING order="15" place="-1" resultid="101108" />
                    <RANKING order="16" place="-1" resultid="101342" />
                    <RANKING order="17" place="-1" resultid="102984" />
                    <RANKING order="18" place="-1" resultid="101945" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99922" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101834" />
                    <RANKING order="2" place="2" resultid="104975" />
                    <RANKING order="3" place="3" resultid="100454" />
                    <RANKING order="4" place="4" resultid="105004" />
                    <RANKING order="5" place="5" resultid="103248" />
                    <RANKING order="6" place="6" resultid="101693" />
                    <RANKING order="7" place="7" resultid="102842" />
                    <RANKING order="8" place="8" resultid="101562" />
                    <RANKING order="9" place="9" resultid="103237" />
                    <RANKING order="10" place="10" resultid="102576" />
                    <RANKING order="11" place="11" resultid="103569" />
                    <RANKING order="12" place="12" resultid="101083" />
                    <RANKING order="13" place="-1" resultid="100723" />
                    <RANKING order="14" place="-1" resultid="101425" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99923" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101612" />
                    <RANKING order="2" place="2" resultid="102385" />
                    <RANKING order="3" place="3" resultid="105046" />
                    <RANKING order="4" place="4" resultid="104389" />
                    <RANKING order="5" place="5" resultid="103018" />
                    <RANKING order="6" place="6" resultid="103326" />
                    <RANKING order="7" place="-1" resultid="101737" />
                    <RANKING order="8" place="-1" resultid="100123" />
                    <RANKING order="9" place="-1" resultid="101254" />
                    <RANKING order="10" place="-1" resultid="101636" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99924" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103506" />
                    <RANKING order="2" place="2" resultid="100947" />
                    <RANKING order="3" place="3" resultid="101671" />
                    <RANKING order="4" place="4" resultid="103196" />
                    <RANKING order="5" place="-1" resultid="100625" />
                    <RANKING order="6" place="-1" resultid="100992" />
                    <RANKING order="7" place="-1" resultid="102015" />
                    <RANKING order="8" place="-1" resultid="102267" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99925" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100273" />
                    <RANKING order="2" place="2" resultid="101774" />
                    <RANKING order="3" place="3" resultid="102197" />
                    <RANKING order="4" place="4" resultid="101032" />
                    <RANKING order="5" place="5" resultid="102639" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99926" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102529" />
                    <RANKING order="2" place="2" resultid="103166" />
                    <RANKING order="3" place="3" resultid="103376" />
                    <RANKING order="4" place="4" resultid="105057" />
                    <RANKING order="5" place="5" resultid="100088" />
                    <RANKING order="6" place="6" resultid="103551" />
                    <RANKING order="7" place="-1" resultid="103159" />
                    <RANKING order="8" place="-1" resultid="102970" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99927" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101681" />
                    <RANKING order="2" place="2" resultid="102978" />
                    <RANKING order="3" place="-1" resultid="103410" />
                    <RANKING order="4" place="-1" resultid="102521" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99928" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100692" />
                    <RANKING order="2" place="2" resultid="104385" />
                    <RANKING order="3" place="3" resultid="100407" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99929" agemax="84" agemin="80" name="KAT.L, 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100998" />
                    <RANKING order="2" place="2" resultid="104994" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99930" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99931" agemax="94" agemin="90" name="KAT.N, 90-94 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100617" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105295" daytime="18:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105296" daytime="18:21" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105297" daytime="18:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105298" daytime="18:29" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="105299" daytime="18:33" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="105300" daytime="18:37" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="105301" daytime="18:40" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="105302" daytime="18:44" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="105303" daytime="18:47" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="105304" daytime="18:51" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="105305" daytime="18:54" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99234" daytime="18:57" gender="F" number="26" order="11" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99526" agemax="96" agemin="80" name="KAT.0, 80-96 lat" calculate="TOTAL" />
                <AGEGROUP agegroupid="99527" agemax="119" agemin="100" name="KAT.A, 100-119 lat" calculate="TOTAL" />
                <AGEGROUP agegroupid="99528" agemax="159" agemin="120" name="KAT.B, 120-159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101875" />
                    <RANKING order="2" place="2" resultid="100253" />
                    <RANKING order="3" place="-1" resultid="104103" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99529" agemax="199" agemin="160" name="KAT.C,160-199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103271" />
                    <RANKING order="2" place="2" resultid="100639" />
                    <RANKING order="3" place="-1" resultid="101372" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99530" agemax="239" agemin="200" name="KAT.D, 200-239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103423" />
                    <RANKING order="2" place="2" resultid="103277" />
                    <RANKING order="3" place="3" resultid="101374" />
                    <RANKING order="4" place="-1" resultid="102763" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99531" agemax="279" agemin="240" name="KAT.E, 240-279 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100734" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99532" agemax="-1" agemin="280" name="KAT.F, 280+ lat" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105306" daytime="18:57" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105307" daytime="19:01" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99250" daytime="19:04" gender="M" number="27" order="12" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99533" agemax="96" agemin="80" name="KAT.0, 80-96 lat" calculate="TOTAL" />
                <AGEGROUP agegroupid="99534" agemax="119" agemin="100" name="KAT.A, 100-119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101876" />
                    <RANKING order="2" place="2" resultid="100328" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99535" agemax="159" agemin="120" name="KAT.B, 120-159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103479" />
                    <RANKING order="2" place="2" resultid="100256" />
                    <RANKING order="3" place="3" resultid="100330" />
                    <RANKING order="4" place="4" resultid="103430" />
                    <RANKING order="5" place="5" resultid="103424" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99536" agemax="199" agemin="160" name="KAT.C,160-199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101428" />
                    <RANKING order="2" place="2" resultid="101877" />
                    <RANKING order="3" place="3" resultid="102221" />
                    <RANKING order="4" place="4" resultid="104105" />
                    <RANKING order="5" place="5" resultid="101112" />
                    <RANKING order="6" place="6" resultid="102870" />
                    <RANKING order="7" place="7" resultid="100257" />
                    <RANKING order="8" place="8" resultid="103283" />
                    <RANKING order="9" place="9" resultid="104106" />
                    <RANKING order="10" place="10" resultid="101114" />
                    <RANKING order="11" place="-1" resultid="101368" />
                    <RANKING order="12" place="-1" resultid="101948" />
                    <RANKING order="13" place="-1" resultid="102223" />
                    <RANKING order="14" place="-1" resultid="102296" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99537" agemax="239" agemin="200" name="KAT.D, 200-239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="104104" />
                    <RANKING order="2" place="2" resultid="103276" />
                    <RANKING order="3" place="3" resultid="100838" />
                    <RANKING order="4" place="4" resultid="101370" />
                    <RANKING order="5" place="5" resultid="102399" />
                    <RANKING order="6" place="-1" resultid="101878" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99538" agemax="279" agemin="240" name="KAT.E, 240-279 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103274" />
                    <RANKING order="2" place="2" resultid="100735" />
                    <RANKING order="3" place="3" resultid="100641" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99539" agemax="-1" agemin="280" name="KAT.F, 280+ lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102219" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105308" daytime="19:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105309" daytime="19:07" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105310" daytime="19:11" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105311" daytime="19:14" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99266" daytime="19:17" gender="F" number="28" order="13" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99932" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102110" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99933" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103563" />
                    <RANKING order="2" place="2" resultid="102176" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99934" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="102959" />
                    <RANKING order="2" place="-1" resultid="103357" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99935" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="105052" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99936" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100703" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99937" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103498" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99938" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100439" />
                    <RANKING order="2" place="2" resultid="102759" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99939" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101995" />
                    <RANKING order="2" place="2" resultid="102702" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99940" agemax="64" agemin="60" name="KAT.H, 60-64 lat" />
                <AGEGROUP agegroupid="99941" agemax="69" agemin="65" name="KAT.I, 65-69 lat" />
                <AGEGROUP agegroupid="99942" agemax="74" agemin="70" name="KAT.J, 70-74 lat" />
                <AGEGROUP agegroupid="99943" agemax="79" agemin="75" name="KAT.K, 75-79 lat" />
                <AGEGROUP agegroupid="99944" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99945" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99946" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="106045" daytime="19:17" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="106046" daytime="19:26" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99282" daytime="19:35" gender="M" number="29" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99947" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100801" />
                    <RANKING order="2" place="2" resultid="104959" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99948" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101147" />
                    <RANKING order="2" place="2" resultid="100288" />
                    <RANKING order="3" place="3" resultid="104384" />
                    <RANKING order="4" place="4" resultid="103025" />
                    <RANKING order="5" place="-1" resultid="105092" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99949" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101011" />
                    <RANKING order="2" place="2" resultid="102379" />
                    <RANKING order="3" place="3" resultid="100281" />
                    <RANKING order="4" place="4" resultid="103540" />
                    <RANKING order="5" place="-1" resultid="102149" />
                    <RANKING order="6" place="-1" resultid="102185" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99950" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102167" />
                    <RANKING order="2" place="2" resultid="101924" />
                    <RANKING order="3" place="3" resultid="100835" />
                    <RANKING order="4" place="4" resultid="101715" />
                    <RANKING order="5" place="5" resultid="101198" />
                    <RANKING order="6" place="6" resultid="100810" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99951" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100765" />
                    <RANKING order="2" place="2" resultid="101182" />
                    <RANKING order="3" place="3" resultid="103399" />
                    <RANKING order="4" place="4" resultid="100783" />
                    <RANKING order="5" place="-1" resultid="101237" />
                    <RANKING order="6" place="-1" resultid="101938" />
                    <RANKING order="7" place="-1" resultid="102985" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99952" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103578" />
                    <RANKING order="2" place="2" resultid="105082" />
                    <RANKING order="3" place="3" resultid="100862" />
                    <RANKING order="4" place="4" resultid="101258" />
                    <RANKING order="5" place="5" resultid="100919" />
                    <RANKING order="6" place="6" resultid="102851" />
                    <RANKING order="7" place="7" resultid="101783" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99953" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103200" />
                    <RANKING order="2" place="2" resultid="104980" />
                    <RANKING order="3" place="3" resultid="100792" />
                    <RANKING order="4" place="4" resultid="103545" />
                    <RANKING order="5" place="5" resultid="102396" />
                    <RANKING order="6" place="6" resultid="102351" />
                    <RANKING order="7" place="-1" resultid="101444" />
                    <RANKING order="8" place="-1" resultid="101662" />
                    <RANKING order="9" place="-1" resultid="103019" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99954" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100559" />
                    <RANKING order="2" place="2" resultid="102571" />
                    <RANKING order="3" place="3" resultid="102016" />
                    <RANKING order="4" place="4" resultid="102031" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99955" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102507" />
                    <RANKING order="2" place="2" resultid="101062" />
                    <RANKING order="3" place="3" resultid="102737" />
                    <RANKING order="4" place="4" resultid="102117" />
                    <RANKING order="5" place="5" resultid="102024" />
                    <RANKING order="6" place="6" resultid="100390" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99956" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100774" />
                    <RANKING order="2" place="2" resultid="101489" />
                    <RANKING order="3" place="3" resultid="100354" />
                    <RANKING order="4" place="4" resultid="101291" />
                    <RANKING order="5" place="5" resultid="105058" />
                    <RANKING order="6" place="6" resultid="102951" />
                    <RANKING order="7" place="7" resultid="103377" />
                    <RANKING order="8" place="8" resultid="101019" />
                    <RANKING order="9" place="-1" resultid="102971" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99957" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100372" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99958" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="101587" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99959" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99960" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99961" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="106047" daytime="19:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="106048" daytime="19:47" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="106049" daytime="19:57" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="106050" daytime="20:06" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="106051" daytime="20:14" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="106052" daytime="20:22" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="106053" daytime="20:29" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99314" daytime="17:16" gender="F" number="22" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99872" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100314" />
                    <RANKING order="2" place="2" resultid="100889" />
                    <RANKING order="3" place="3" resultid="100910" />
                    <RANKING order="4" place="-1" resultid="104380" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99873" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103392" />
                    <RANKING order="2" place="2" resultid="102943" />
                    <RANKING order="3" place="3" resultid="101168" />
                    <RANKING order="4" place="4" resultid="101789" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99874" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103520" />
                    <RANKING order="2" place="2" resultid="100584" />
                    <RANKING order="3" place="-1" resultid="102958" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99875" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100168" />
                    <RANKING order="2" place="2" resultid="101688" />
                    <RANKING order="3" place="-1" resultid="101705" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99876" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100612" />
                    <RANKING order="2" place="2" resultid="100236" />
                    <RANKING order="3" place="3" resultid="103127" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99877" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100728" />
                    <RANKING order="2" place="2" resultid="103428" />
                    <RANKING order="3" place="3" resultid="101075" />
                    <RANKING order="4" place="4" resultid="100875" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99878" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101461" />
                    <RANKING order="2" place="2" resultid="100591" />
                    <RANKING order="3" place="3" resultid="103116" />
                    <RANKING order="4" place="-1" resultid="101329" />
                    <RANKING order="5" place="-1" resultid="103102" />
                    <RANKING order="6" place="-1" resultid="103108" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99879" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101994" />
                    <RANKING order="2" place="2" resultid="105023" />
                    <RANKING order="3" place="-1" resultid="100937" />
                    <RANKING order="4" place="-1" resultid="101295" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99880" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100448" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99881" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101570" />
                    <RANKING order="2" place="2" resultid="101496" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99882" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100688" />
                    <RANKING order="2" place="2" resultid="102743" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99883" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101574" />
                    <RANKING order="2" place="-1" resultid="100465" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99884" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99885" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99886" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105277" daytime="17:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105278" daytime="17:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105279" daytime="17:23" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105280" daytime="17:26" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2014-06-29" daytime="09:00" number="4" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="99344" daytime="09:00" gender="F" number="30" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99962" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100197" />
                    <RANKING order="2" place="2" resultid="100911" />
                    <RANKING order="3" place="-1" resultid="103063" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99963" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103140" />
                    <RANKING order="2" place="2" resultid="103564" />
                    <RANKING order="3" place="3" resultid="102177" />
                    <RANKING order="4" place="4" resultid="101595" />
                    <RANKING order="5" place="5" resultid="101628" />
                    <RANKING order="6" place="6" resultid="101620" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99964" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101710" />
                    <RANKING order="2" place="2" resultid="103528" />
                    <RANKING order="3" place="-1" resultid="102293" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99965" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="101307" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99966" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100613" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99967" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100820" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99968" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100592" />
                    <RANKING order="2" place="2" resultid="100440" />
                    <RANKING order="3" place="-1" resultid="101450" />
                    <RANKING order="4" place="-1" resultid="102552" />
                    <RANKING order="5" place="-1" resultid="102760" />
                    <RANKING order="6" place="-1" resultid="103109" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99969" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102724" />
                    <RANKING order="2" place="2" resultid="105103" />
                    <RANKING order="3" place="3" resultid="102784" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99970" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102716" />
                    <RANKING order="2" place="2" resultid="101439" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99971" agemax="69" agemin="65" name="KAT.I, 65-69 lat" />
                <AGEGROUP agegroupid="99972" agemax="74" agemin="70" name="KAT.J, 70-74 lat" />
                <AGEGROUP agegroupid="99973" agemax="79" agemin="75" name="KAT.K, 75-79 lat" />
                <AGEGROUP agegroupid="99974" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99975" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99976" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105321" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105322" daytime="09:03" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105323" daytime="09:06" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99361" daytime="09:08" gender="M" number="31" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99977" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100902" />
                    <RANKING order="2" place="2" resultid="104960" />
                    <RANKING order="3" place="-1" resultid="103032" />
                    <RANKING order="4" place="-1" resultid="103045" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99978" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102281" />
                    <RANKING order="2" place="2" resultid="101005" />
                    <RANKING order="3" place="3" resultid="101728" />
                    <RANKING order="4" place="4" resultid="100321" />
                    <RANKING order="5" place="5" resultid="101826" />
                    <RANKING order="6" place="-1" resultid="103013" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99979" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102067" />
                    <RANKING order="2" place="2" resultid="102993" />
                    <RANKING order="3" place="3" resultid="101054" />
                    <RANKING order="4" place="4" resultid="102210" />
                    <RANKING order="5" place="-1" resultid="102150" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99980" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102824" />
                    <RANKING order="2" place="2" resultid="101925" />
                    <RANKING order="3" place="3" resultid="101716" />
                    <RANKING order="4" place="4" resultid="104404" />
                    <RANKING order="5" place="5" resultid="100293" />
                    <RANKING order="6" place="6" resultid="101819" />
                    <RANKING order="7" place="7" resultid="102250" />
                    <RANKING order="8" place="8" resultid="100110" />
                    <RANKING order="9" place="-1" resultid="100224" />
                    <RANKING order="10" place="-1" resultid="102168" />
                    <RANKING order="11" place="-1" resultid="102966" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99981" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100766" />
                    <RANKING order="2" place="2" resultid="101406" />
                    <RANKING order="3" place="3" resultid="103515" />
                    <RANKING order="4" place="4" resultid="100474" />
                    <RANKING order="5" place="5" resultid="103400" />
                    <RANKING order="6" place="6" resultid="100216" />
                    <RANKING order="7" place="7" resultid="102515" />
                    <RANKING order="8" place="-1" resultid="100246" />
                    <RANKING order="9" place="-1" resultid="101939" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99982" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="105005" />
                    <RANKING order="2" place="2" resultid="101835" />
                    <RANKING order="3" place="3" resultid="101468" />
                    <RANKING order="4" place="4" resultid="102843" />
                    <RANKING order="5" place="5" resultid="100828" />
                    <RANKING order="6" place="6" resultid="103570" />
                    <RANKING order="7" place="7" resultid="101257" />
                    <RANKING order="8" place="8" resultid="100863" />
                    <RANKING order="9" place="9" resultid="101784" />
                    <RANKING order="10" place="-1" resultid="100455" />
                    <RANKING order="11" place="-1" resultid="100480" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99983" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103201" />
                    <RANKING order="2" place="2" resultid="100132" />
                    <RANKING order="3" place="3" resultid="104981" />
                    <RANKING order="4" place="4" resultid="102352" />
                    <RANKING order="5" place="-1" resultid="100124" />
                    <RANKING order="6" place="-1" resultid="101663" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99984" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102262" />
                    <RANKING order="2" place="2" resultid="100626" />
                    <RANKING order="3" place="3" resultid="100560" />
                    <RANKING order="4" place="4" resultid="102017" />
                    <RANKING order="5" place="5" resultid="102049" />
                    <RANKING order="6" place="6" resultid="101091" />
                    <RANKING order="7" place="-1" resultid="100605" />
                    <RANKING order="8" place="-1" resultid="100931" />
                    <RANKING order="9" place="-1" resultid="100948" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99985" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102198" />
                    <RANKING order="2" place="2" resultid="100382" />
                    <RANKING order="3" place="3" resultid="102118" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99986" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102530" />
                    <RANKING order="2" place="2" resultid="100355" />
                    <RANKING order="3" place="3" resultid="100577" />
                    <RANKING order="4" place="4" resultid="101292" />
                    <RANKING order="5" place="5" resultid="103378" />
                    <RANKING order="6" place="6" resultid="102952" />
                    <RANKING order="7" place="7" resultid="105059" />
                    <RANKING order="8" place="8" resultid="101020" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99987" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100140" />
                    <RANKING order="2" place="2" resultid="100373" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99988" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="101588" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99989" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="99990" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="99991" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105324" daytime="09:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105325" daytime="09:12" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105326" daytime="09:16" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105327" daytime="09:18" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="105328" daytime="09:21" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="105329" daytime="09:23" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="105330" daytime="09:26" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="105331" daytime="09:28" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99377" daytime="09:30" gender="F" number="32" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99992" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100890" />
                    <RANKING order="2" place="2" resultid="102111" />
                    <RANKING order="3" place="3" resultid="104381" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99993" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103393" />
                    <RANKING order="2" place="2" resultid="101170" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99994" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103521" />
                    <RANKING order="2" place="-1" resultid="102960" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99995" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100169" />
                    <RANKING order="2" place="2" resultid="101706" />
                    <RANKING order="3" place="3" resultid="101690" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99996" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100238" />
                    <RANKING order="2" place="2" resultid="103128" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99997" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="105017" />
                    <RANKING order="2" place="2" resultid="100729" />
                    <RANKING order="3" place="3" resultid="103429" />
                    <RANKING order="4" place="4" resultid="101077" />
                    <RANKING order="5" place="5" resultid="100876" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99998" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101463" />
                    <RANKING order="2" place="2" resultid="100593" />
                    <RANKING order="3" place="-1" resultid="101330" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99999" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="105024" />
                    <RANKING order="2" place="2" resultid="101996" />
                    <RANKING order="3" place="3" resultid="102703" />
                    <RANKING order="4" place="4" resultid="102793" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100000" agemax="64" agemin="60" name="KAT.H, 60-64 lat" />
                <AGEGROUP agegroupid="100001" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101497" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100002" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100689" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100003" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101575" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100004" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="100005" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="100006" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105332" daytime="09:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105333" daytime="09:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105334" daytime="09:41" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99393" daytime="09:45" gender="M" number="33" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="100007" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100973" />
                    <RANKING order="2" place="2" resultid="104961" />
                    <RANKING order="3" place="3" resultid="100802" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100008" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103444" />
                    <RANKING order="2" place="2" resultid="101148" />
                    <RANKING order="3" place="3" resultid="101006" />
                    <RANKING order="4" place="4" resultid="101647" />
                    <RANKING order="5" place="-1" resultid="102868" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100009" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101012" />
                    <RANKING order="2" place="2" resultid="102372" />
                    <RANKING order="3" place="3" resultid="102889" />
                    <RANKING order="4" place="-1" resultid="101043" />
                    <RANKING order="5" place="-1" resultid="102068" />
                    <RANKING order="6" place="-1" resultid="102186" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100010" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102825" />
                    <RANKING order="2" place="2" resultid="100757" />
                    <RANKING order="3" place="3" resultid="101199" />
                    <RANKING order="4" place="4" resultid="103053" />
                    <RANKING order="5" place="5" resultid="103449" />
                    <RANKING order="6" place="6" resultid="102191" />
                    <RANKING order="7" place="7" resultid="101717" />
                    <RANKING order="8" place="8" resultid="100811" />
                    <RANKING order="9" place="9" resultid="102103" />
                    <RANKING order="10" place="10" resultid="104405" />
                    <RANKING order="11" place="11" resultid="100111" />
                    <RANKING order="12" place="-1" resultid="102169" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100011" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101192" />
                    <RANKING order="2" place="2" resultid="100767" />
                    <RANKING order="3" place="3" resultid="101476" />
                    <RANKING order="4" place="4" resultid="101183" />
                    <RANKING order="5" place="5" resultid="101416" />
                    <RANKING order="6" place="6" resultid="100784" />
                    <RANKING order="7" place="-1" resultid="101933" />
                    <RANKING order="8" place="-1" resultid="102042" />
                    <RANKING order="9" place="-1" resultid="105037" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100012" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100724" />
                    <RANKING order="2" place="2" resultid="102359" />
                    <RANKING order="3" place="3" resultid="101701" />
                    <RANKING order="4" place="4" resultid="100399" />
                    <RANKING order="5" place="5" resultid="103579" />
                    <RANKING order="6" place="6" resultid="100829" />
                    <RANKING order="7" place="7" resultid="101426" />
                    <RANKING order="8" place="8" resultid="100920" />
                    <RANKING order="9" place="9" resultid="102852" />
                    <RANKING order="10" place="-1" resultid="104969" />
                    <RANKING order="11" place="-1" resultid="100461" />
                    <RANKING order="12" place="-1" resultid="103244" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100013" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100133" />
                    <RANKING order="2" place="2" resultid="100793" />
                    <RANKING order="3" place="3" resultid="104390" />
                    <RANKING order="4" place="-1" resultid="100661" />
                    <RANKING order="5" place="-1" resultid="101664" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100014" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103507" />
                    <RANKING order="2" place="2" resultid="102572" />
                    <RANKING order="3" place="3" resultid="101161" />
                    <RANKING order="4" place="4" resultid="105392" />
                    <RANKING order="5" place="-1" resultid="100627" />
                    <RANKING order="6" place="-1" resultid="100675" />
                    <RANKING order="7" place="-1" resultid="102832" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100015" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101580" />
                    <RANKING order="2" place="2" resultid="101775" />
                    <RANKING order="3" place="3" resultid="100383" />
                    <RANKING order="4" place="4" resultid="101033" />
                    <RANKING order="5" place="5" resultid="101063" />
                    <RANKING order="6" place="6" resultid="102565" />
                    <RANKING order="7" place="7" resultid="102025" />
                    <RANKING order="8" place="8" resultid="100391" />
                    <RANKING order="9" place="9" resultid="100895" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100016" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101490" />
                    <RANKING order="2" place="2" resultid="100775" />
                    <RANKING order="3" place="3" resultid="100679" />
                    <RANKING order="4" place="4" resultid="102953" />
                    <RANKING order="5" place="5" resultid="103404" />
                    <RANKING order="6" place="6" resultid="101337" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100017" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102560" />
                    <RANKING order="2" place="2" resultid="102979" />
                    <RANKING order="3" place="3" resultid="100374" />
                    <RANKING order="4" place="-1" resultid="101682" />
                    <RANKING order="5" place="-1" resultid="102143" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100018" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102750" />
                    <RANKING order="2" place="2" resultid="100408" />
                    <RANKING order="3" place="-1" resultid="101589" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100019" agemax="84" agemin="80" name="KAT.L, 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100999" />
                    <RANKING order="2" place="2" resultid="104991" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100020" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="100021" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105335" daytime="09:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105336" daytime="09:52" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105337" daytime="09:59" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105338" daytime="10:04" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="105339" daytime="10:08" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="105340" daytime="10:13" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="105341" daytime="10:17" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="105342" daytime="10:20" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="105343" daytime="10:24" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99409" daytime="10:27" gender="F" number="34" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="100022" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103002" />
                    <RANKING order="2" place="2" resultid="103473" />
                    <RANKING order="3" place="3" resultid="100912" />
                    <RANKING order="4" place="-1" resultid="103064" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100023" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102178" />
                    <RANKING order="2" place="2" resultid="102945" />
                    <RANKING order="3" place="3" resultid="103565" />
                    <RANKING order="4" place="4" resultid="102501" />
                    <RANKING order="5" place="-1" resultid="102391" />
                    <RANKING order="6" place="-1" resultid="102910" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100024" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="105094" />
                    <RANKING order="2" place="2" resultid="103358" />
                    <RANKING order="3" place="-1" resultid="102961" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100025" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101244" />
                    <RANKING order="2" place="2" resultid="100170" />
                    <RANKING order="3" place="3" resultid="100186" />
                    <RANKING order="4" place="4" resultid="102096" />
                    <RANKING order="5" place="5" resultid="100884" />
                    <RANKING order="6" place="6" resultid="102799" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100026" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102055" />
                    <RANKING order="2" place="2" resultid="101803" />
                    <RANKING order="3" place="3" resultid="101359" />
                    <RANKING order="4" place="4" resultid="103335" />
                    <RANKING order="5" place="5" resultid="100117" />
                    <RANKING order="6" place="-1" resultid="103067" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100027" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103352" />
                    <RANKING order="2" place="2" resultid="105032" />
                    <RANKING order="3" place="3" resultid="100821" />
                    <RANKING order="4" place="4" resultid="103499" />
                    <RANKING order="5" place="5" resultid="100877" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100028" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100633" />
                    <RANKING order="2" place="2" resultid="101748" />
                    <RANKING order="3" place="3" resultid="103467" />
                    <RANKING order="4" place="4" resultid="103117" />
                    <RANKING order="5" place="5" resultid="102459" />
                    <RANKING order="6" place="6" resultid="102761" />
                    <RANKING order="7" place="7" resultid="100429" />
                    <RANKING order="8" place="-1" resultid="103103" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100029" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103415" />
                    <RANKING order="2" place="2" resultid="102546" />
                    <RANKING order="3" place="3" resultid="103085" />
                    <RANKING order="4" place="4" resultid="102725" />
                    <RANKING order="5" place="5" resultid="103091" />
                    <RANKING order="6" place="6" resultid="105064" />
                    <RANKING order="7" place="7" resultid="102794" />
                    <RANKING order="8" place="8" resultid="102785" />
                    <RANKING order="9" place="-1" resultid="100939" />
                    <RANKING order="10" place="-1" resultid="101298" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100030" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102717" />
                    <RANKING order="2" place="2" resultid="102538" />
                    <RANKING order="3" place="3" resultid="102464" />
                    <RANKING order="4" place="4" resultid="101440" />
                    <RANKING order="5" place="5" resultid="100449" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100031" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101455" />
                    <RANKING order="2" place="2" resultid="101286" />
                    <RANKING order="3" place="3" resultid="103387" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100032" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100714" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100033" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="105028" />
                    <RANKING order="2" place="2" resultid="103080" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100034" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="100035" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="100036" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105344" daytime="10:27" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105345" daytime="10:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105346" daytime="10:31" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105347" daytime="10:33" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="105348" daytime="10:35" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="105349" daytime="10:37" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99425" daytime="10:38" gender="M" number="35" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="100037" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102906" />
                    <RANKING order="2" place="2" resultid="103033" />
                    <RANKING order="3" place="-1" resultid="103046" />
                    <RANKING order="4" place="-1" resultid="102810" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100038" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100162" />
                    <RANKING order="2" place="2" resultid="101764" />
                    <RANKING order="3" place="3" resultid="101175" />
                    <RANKING order="4" place="4" resultid="101827" />
                    <RANKING order="5" place="5" resultid="100302" />
                    <RANKING order="6" place="6" resultid="102487" />
                    <RANKING order="7" place="-1" resultid="101302" />
                    <RANKING order="8" place="-1" resultid="102485" />
                    <RANKING order="9" place="-1" resultid="103014" />
                    <RANKING order="10" place="-1" resultid="103440" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100039" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103454" />
                    <RANKING order="2" place="2" resultid="101733" />
                    <RANKING order="3" place="3" resultid="103541" />
                    <RANKING order="4" place="4" resultid="102380" />
                    <RANKING order="5" place="5" resultid="100155" />
                    <RANKING order="6" place="6" resultid="101252" />
                    <RANKING order="7" place="7" resultid="102994" />
                    <RANKING order="8" place="8" resultid="103602" />
                    <RANKING order="9" place="9" resultid="100327" />
                    <RANKING order="10" place="10" resultid="102215" />
                    <RANKING order="11" place="11" resultid="100308" />
                    <RANKING order="12" place="-1" resultid="101222" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100040" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102074" />
                    <RANKING order="2" place="2" resultid="102159" />
                    <RANKING order="3" place="3" resultid="100836" />
                    <RANKING order="4" place="4" resultid="101267" />
                    <RANKING order="5" place="5" resultid="100598" />
                    <RANKING order="6" place="6" resultid="101602" />
                    <RANKING order="7" place="7" resultid="102584" />
                    <RANKING order="8" place="8" resultid="103054" />
                    <RANKING order="9" place="9" resultid="100758" />
                    <RANKING order="10" place="10" resultid="102479" />
                    <RANKING order="11" place="11" resultid="102256" />
                    <RANKING order="12" place="-1" resultid="102916" />
                    <RANKING order="13" place="-1" resultid="103260" />
                    <RANKING order="14" place="-1" resultid="103265" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100041" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101354" />
                    <RANKING order="2" place="2" resultid="101238" />
                    <RANKING order="3" place="3" resultid="100191" />
                    <RANKING order="4" place="4" resultid="100987" />
                    <RANKING order="5" place="5" resultid="100247" />
                    <RANKING order="6" place="6" resultid="100785" />
                    <RANKING order="7" place="-1" resultid="102482" />
                    <RANKING order="8" place="-1" resultid="100657" />
                    <RANKING order="9" place="-1" resultid="100962" />
                    <RANKING order="10" place="-1" resultid="101205" />
                    <RANKING order="11" place="-1" resultid="101217" />
                    <RANKING order="12" place="-1" resultid="102043" />
                    <RANKING order="13" place="-1" resultid="105086" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100042" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101039" />
                    <RANKING order="2" place="2" resultid="101754" />
                    <RANKING order="3" place="3" resultid="105006" />
                    <RANKING order="4" place="4" resultid="103615" />
                    <RANKING order="5" place="5" resultid="101421" />
                    <RANKING order="6" place="6" resultid="101643" />
                    <RANKING order="7" place="7" resultid="100864" />
                    <RANKING order="8" place="8" resultid="100921" />
                    <RANKING order="9" place="9" resultid="103557" />
                    <RANKING order="10" place="10" resultid="101785" />
                    <RANKING order="11" place="11" resultid="100468" />
                    <RANKING order="12" place="-1" resultid="101333" />
                    <RANKING order="13" place="-1" resultid="101563" />
                    <RANKING order="14" place="-1" resultid="102004" />
                    <RANKING order="15" place="-1" resultid="102469" />
                    <RANKING order="16" place="-1" resultid="102577" />
                    <RANKING order="17" place="-1" resultid="102848" />
                    <RANKING order="18" place="-1" resultid="103074" />
                    <RANKING order="19" place="-1" resultid="103231" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100043" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101613" />
                    <RANKING order="2" place="2" resultid="101501" />
                    <RANKING order="3" place="3" resultid="101482" />
                    <RANKING order="4" place="4" resultid="102860" />
                    <RANKING order="5" place="5" resultid="102365" />
                    <RANKING order="6" place="6" resultid="104982" />
                    <RANKING order="7" place="7" resultid="103208" />
                    <RANKING order="8" place="8" resultid="103215" />
                    <RANKING order="9" place="9" resultid="103327" />
                    <RANKING order="10" place="10" resultid="103221" />
                    <RANKING order="11" place="-1" resultid="103020" />
                    <RANKING order="12" place="-1" resultid="103226" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100044" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102268" />
                    <RANKING order="2" place="2" resultid="100561" />
                    <RANKING order="3" place="3" resultid="103191" />
                    <RANKING order="4" place="4" resultid="100606" />
                    <RANKING order="5" place="5" resultid="102038" />
                    <RANKING order="6" place="6" resultid="102050" />
                    <RANKING order="7" place="7" resultid="103364" />
                    <RANKING order="8" place="-1" resultid="100932" />
                    <RANKING order="9" place="-1" resultid="106116" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100045" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102508" />
                    <RANKING order="2" place="2" resultid="101276" />
                    <RANKING order="3" place="3" resultid="102204" />
                    <RANKING order="4" place="4" resultid="105011" />
                    <RANKING order="5" place="5" resultid="104374" />
                    <RANKING order="6" place="6" resultid="102640" />
                    <RANKING order="7" place="7" resultid="102124" />
                    <RANKING order="8" place="8" resultid="102738" />
                    <RANKING order="9" place="9" resultid="103588" />
                    <RANKING order="10" place="10" resultid="102119" />
                    <RANKING order="11" place="-1" resultid="101325" />
                    <RANKING order="12" place="-1" resultid="103174" />
                    <RANKING order="13" place="-1" resultid="103179" />
                    <RANKING order="14" place="-1" resultid="103185" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100046" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102466" />
                    <RANKING order="2" place="2" resultid="100567" />
                    <RANKING order="3" place="3" resultid="100571" />
                    <RANKING order="4" place="4" resultid="100356" />
                    <RANKING order="5" place="5" resultid="103167" />
                    <RANKING order="6" place="6" resultid="102132" />
                    <RANKING order="7" place="7" resultid="101021" />
                    <RANKING order="8" place="8" resultid="101743" />
                    <RANKING order="9" place="-1" resultid="103152" />
                    <RANKING order="10" place="-1" resultid="103160" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100047" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100141" />
                    <RANKING order="2" place="2" resultid="100709" />
                    <RANKING order="3" place="3" resultid="102522" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100048" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102751" />
                    <RANKING order="2" place="2" resultid="100409" />
                    <RANKING order="3" place="3" resultid="102137" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100049" agemax="84" agemin="80" name="KAT.L, 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102709" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100050" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="100051" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105350" daytime="10:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105351" daytime="10:41" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105352" daytime="10:44" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="105353" daytime="10:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="105354" daytime="10:47" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="105355" daytime="10:49" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="105356" daytime="10:51" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="105357" daytime="10:52" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="105358" daytime="10:54" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="105359" daytime="10:56" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="105360" daytime="10:57" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="105361" daytime="10:59" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="105362" daytime="11:00" number="13" order="13" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99441" daytime="11:02" gender="X" number="36" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="99540" agemax="96" agemin="80" name="KAT.0, 80-96 lat" calculate="TOTAL" />
                <AGEGROUP agegroupid="99541" agemax="119" agemin="100" name="KAT.A, 100-119 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101880" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99542" agemax="159" agemin="120" name="KAT.B, 120-159 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101879" />
                    <RANKING order="2" place="2" resultid="104107" />
                    <RANKING order="3" place="3" resultid="100250" />
                    <RANKING order="4" place="4" resultid="103421" />
                    <RANKING order="5" place="5" resultid="106117" />
                    <RANKING order="6" place="-1" resultid="101362" />
                    <RANKING order="7" place="-1" resultid="102217" />
                    <RANKING order="8" place="-1" resultid="103282" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99543" agemax="199" agemin="160" name="KAT.C,160-199 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101375" />
                    <RANKING order="2" place="2" resultid="100635" />
                    <RANKING order="3" place="3" resultid="103419" />
                    <RANKING order="4" place="4" resultid="103267" />
                    <RANKING order="5" place="5" resultid="100251" />
                    <RANKING order="6" place="6" resultid="102489" />
                    <RANKING order="7" place="7" resultid="104108" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99544" agemax="239" agemin="200" name="KAT.D, 200-239 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103280" />
                    <RANKING order="2" place="2" resultid="102586" />
                    <RANKING order="3" place="3" resultid="100637" />
                    <RANKING order="4" place="4" resultid="105066" />
                    <RANKING order="5" place="-1" resultid="101364" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99545" agemax="279" agemin="240" name="KAT.E, 240-279 lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103269" />
                    <RANKING order="2" place="2" resultid="105040" />
                    <RANKING order="3" place="3" resultid="101366" />
                    <RANKING order="4" place="4" resultid="103417" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="99546" agemax="-1" agemin="280" name="KAT.F, 280+ lat" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100736" />
                    <RANKING order="2" place="2" resultid="102764" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="105363" daytime="11:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="105364" daytime="11:06" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="105365" daytime="11:10" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99457" daytime="11:13" gender="F" number="37" order="8" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="100052" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103003" />
                    <RANKING order="2" place="2" resultid="103612" />
                    <RANKING order="3" place="3" resultid="100315" />
                    <RANKING order="4" place="4" resultid="105071" />
                    <RANKING order="5" place="-1" resultid="101723" />
                    <RANKING order="6" place="-1" resultid="102112" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100053" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102288" />
                    <RANKING order="2" place="2" resultid="101142" />
                    <RANKING order="3" place="3" resultid="103394" />
                    <RANKING order="4" place="4" resultid="101596" />
                    <RANKING order="5" place="5" resultid="102502" />
                    <RANKING order="6" place="6" resultid="101629" />
                    <RANKING order="7" place="7" resultid="101621" />
                    <RANKING order="8" place="8" resultid="101790" />
                    <RANKING order="9" place="9" resultid="100435" />
                    <RANKING order="10" place="-1" resultid="101349" />
                    <RANKING order="11" place="-1" resultid="103146" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100054" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103535" />
                    <RANKING order="2" place="2" resultid="103529" />
                    <RANKING order="3" place="3" resultid="101853" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100055" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100926" />
                    <RANKING order="2" place="2" resultid="100182" />
                    <RANKING order="3" place="3" resultid="100176" />
                    <RANKING order="4" place="4" resultid="100885" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100056" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100704" />
                    <RANKING order="2" place="2" resultid="103135" />
                    <RANKING order="3" place="3" resultid="100239" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100057" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="105018" />
                    <RANKING order="2" place="2" resultid="103500" />
                    <RANKING order="3" place="-1" resultid="100552" />
                    <RANKING order="4" place="-1" resultid="101078" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100058" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101464" />
                    <RANKING order="2" place="2" resultid="102732" />
                    <RANKING order="3" place="3" resultid="100441" />
                    <RANKING order="4" place="-1" resultid="100543" />
                    <RANKING order="5" place="-1" resultid="102553" />
                    <RANKING order="6" place="-1" resultid="103097" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100059" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103092" />
                    <RANKING order="2" place="2" resultid="101997" />
                    <RANKING order="3" place="3" resultid="100940" />
                    <RANKING order="4" place="-1" resultid="102704" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100060" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100956" />
                    <RANKING order="2" place="2" resultid="100450" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100061" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101843" />
                    <RANKING order="2" place="2" resultid="103388" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100062" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100715" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100063" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101471" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100064" agemax="84" agemin="80" name="KAT.L, 80-84 lat" />
                <AGEGROUP agegroupid="100065" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="100066" agemax="94" agemin="90" name="KAT.N, 90-94 lat" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="106054" daytime="11:13" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="106055" daytime="11:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="106056" daytime="11:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="106057" daytime="11:41" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="99473" daytime="11:54" gender="M" number="38" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="100067" agemax="24" agemin="20" name="KAT.0, 20-24 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100903" />
                    <RANKING order="2" place="2" resultid="102907" />
                    <RANKING order="3" place="3" resultid="100803" />
                    <RANKING order="4" place="4" resultid="100683" />
                    <RANKING order="5" place="-1" resultid="102811" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100068" agemax="29" agemin="25" name="KAT.A, 25-29 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102282" />
                    <RANKING order="2" place="2" resultid="101154" />
                    <RANKING order="3" place="3" resultid="105093" />
                    <RANKING order="4" place="4" resultid="100289" />
                    <RANKING order="5" place="5" resultid="103459" />
                    <RANKING order="6" place="6" resultid="101860" />
                    <RANKING order="7" place="7" resultid="100322" />
                    <RANKING order="8" place="-1" resultid="101104" />
                    <RANKING order="9" place="-1" resultid="101231" />
                    <RANKING order="10" place="-1" resultid="103370" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100069" agemax="34" agemin="30" name="KAT.B, 30-34 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101013" />
                    <RANKING order="2" place="2" resultid="102381" />
                    <RANKING order="3" place="3" resultid="100282" />
                    <RANKING order="4" place="4" resultid="100869" />
                    <RANKING order="5" place="5" resultid="101055" />
                    <RANKING order="6" place="6" resultid="101655" />
                    <RANKING order="7" place="-1" resultid="105391" />
                    <RANKING order="8" place="-1" resultid="101796" />
                    <RANKING order="9" place="-1" resultid="102151" />
                    <RANKING order="10" place="-1" resultid="102187" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100070" agemax="39" agemin="35" name="KAT.C, 35-39 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102160" />
                    <RANKING order="2" place="2" resultid="102884" />
                    <RANKING order="3" place="3" resultid="101926" />
                    <RANKING order="4" place="4" resultid="100415" />
                    <RANKING order="5" place="5" resultid="101135" />
                    <RANKING order="6" place="-1" resultid="100812" />
                    <RANKING order="7" place="-1" resultid="101200" />
                    <RANKING order="8" place="-1" resultid="101813" />
                    <RANKING order="9" place="-1" resultid="102009" />
                    <RANKING order="10" place="-1" resultid="102967" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100071" agemax="44" agemin="40" name="KAT.D, 40-44 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101218" />
                    <RANKING order="2" place="2" resultid="101239" />
                    <RANKING order="3" place="3" resultid="103254" />
                    <RANKING order="4" place="4" resultid="103516" />
                    <RANKING order="5" place="5" resultid="101411" />
                    <RANKING order="6" place="6" resultid="101184" />
                    <RANKING order="7" place="7" resultid="100217" />
                    <RANKING order="8" place="8" resultid="103594" />
                    <RANKING order="9" place="9" resultid="100203" />
                    <RANKING order="10" place="10" resultid="102516" />
                    <RANKING order="11" place="11" resultid="101606" />
                    <RANKING order="12" place="-1" resultid="105038" />
                    <RANKING order="13" place="-1" resultid="101193" />
                    <RANKING order="14" place="-1" resultid="101343" />
                    <RANKING order="15" place="-1" resultid="101946" />
                    <RANKING order="16" place="-1" resultid="102986" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100072" agemax="49" agemin="45" name="KAT.E, 45-49 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100456" />
                    <RANKING order="2" place="2" resultid="104976" />
                    <RANKING order="3" place="3" resultid="101694" />
                    <RANKING order="4" place="4" resultid="103249" />
                    <RANKING order="5" place="5" resultid="105083" />
                    <RANKING order="6" place="6" resultid="103580" />
                    <RANKING order="7" place="7" resultid="103238" />
                    <RANKING order="8" place="8" resultid="102853" />
                    <RANKING order="9" place="9" resultid="103571" />
                    <RANKING order="10" place="-1" resultid="101564" />
                    <RANKING order="11" place="-1" resultid="101836" />
                    <RANKING order="12" place="-1" resultid="101256" />
                    <RANKING order="13" place="-1" resultid="104970" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100073" agemax="54" agemin="50" name="KAT.F, 50-54 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101614" />
                    <RANKING order="2" place="2" resultid="102386" />
                    <RANKING order="3" place="3" resultid="103202" />
                    <RANKING order="4" place="4" resultid="105047" />
                    <RANKING order="5" place="5" resultid="103546" />
                    <RANKING order="6" place="6" resultid="102397" />
                    <RANKING order="7" place="7" resultid="102353" />
                    <RANKING order="8" place="-1" resultid="100794" />
                    <RANKING order="9" place="-1" resultid="101255" />
                    <RANKING order="10" place="-1" resultid="103021" />
                    <RANKING order="11" place="-1" resultid="103328" />
                    <RANKING order="12" place="-1" resultid="104391" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100074" agemax="59" agemin="55" name="KAT.G, 55-59 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103508" />
                    <RANKING order="2" place="2" resultid="100949" />
                    <RANKING order="3" place="3" resultid="102018" />
                    <RANKING order="4" place="4" resultid="101162" />
                    <RANKING order="5" place="5" resultid="101672" />
                    <RANKING order="6" place="6" resultid="103197" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100075" agemax="64" agemin="60" name="KAT.H, 60-64 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101776" />
                    <RANKING order="2" place="2" resultid="102199" />
                    <RANKING order="3" place="3" resultid="101064" />
                    <RANKING order="4" place="4" resultid="101034" />
                    <RANKING order="5" place="5" resultid="100392" />
                    <RANKING order="6" place="6" resultid="102641" />
                    <RANKING order="7" place="-1" resultid="100274" />
                    <RANKING order="8" place="-1" resultid="102566" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100076" agemax="69" agemin="65" name="KAT.I, 65-69 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="103168" />
                    <RANKING order="2" place="2" resultid="100776" />
                    <RANKING order="3" place="3" resultid="101491" />
                    <RANKING order="4" place="4" resultid="103379" />
                    <RANKING order="5" place="5" resultid="105060" />
                    <RANKING order="6" place="6" resultid="100089" />
                    <RANKING order="7" place="7" resultid="103552" />
                    <RANKING order="8" place="-1" resultid="103405" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100077" agemax="74" agemin="70" name="KAT.J, 70-74 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="102972" />
                    <RANKING order="2" place="2" resultid="101683" />
                    <RANKING order="3" place="3" resultid="103411" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100078" agemax="79" agemin="75" name="KAT.K, 75-79 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="100693" />
                    <RANKING order="2" place="2" resultid="100982" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100079" agemax="84" agemin="80" name="KAT.L, 80-84 lat">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="101000" />
                    <RANKING order="2" place="2" resultid="104995" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="100080" agemax="89" agemin="85" name="KAT.M, 85-89 lat" />
                <AGEGROUP agegroupid="100081" agemax="94" agemin="90" name="KAT.N, 90-94 lat">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="100618" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="106059" daytime="11:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="106060" daytime="12:08" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="106061" daytime="12:17" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="106062" daytime="12:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="106063" daytime="12:33" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="106064" daytime="12:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="106065" daytime="12:46" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="106066" daytime="12:53" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="106067" daytime="12:59" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" nation="POL" clubid="101201" name="10 Brygada Kawalerii Panc. Świętoszów" shortname="10 BK Panc. Świętoszów">
          <CONTACT city="Świdnica" email="horbacz.marcin@wp.pl" name="Horbacz Marcin" state="LBS" street="Buchałów 12c" zip="66-008" />
          <ATHLETES>
            <ATHLETE birthdate="1974-12-15" firstname="Oskar" gender="M" lastname="BOGUCKI" nation="POL" athleteid="101202">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="101203" heatid="105132" lane="9" entrytime="00:00:31.00" entrycourse="LCM" />
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="101204" heatid="105255" lane="2" entrytime="00:01:22.00" entrycourse="LCM" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="101205" heatid="105357" lane="3" entrytime="00:00:38.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-03-14" firstname="Jarosław" gender="M" lastname="DRUCIAREK" nation="POL" swrid="4992762" athleteid="101206">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="101207" heatid="105136" lane="0" entrytime="00:00:29.00" entrycourse="LCM" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="101208" heatid="105219" lane="3" entrytime="00:01:10.00" entrycourse="LCM" />
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="101209" heatid="105267" lane="6" entrytime="00:00:39.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-06-16" firstname="Marcin" gender="M" lastname="Horbacz" nation="POL" swrid="4992761" athleteid="101210">
              <RESULTS>
                <RESULT eventid="98798" points="442" reactiontime="+90" swimtime="00:00:27.43" resultid="101211" heatid="105123" lane="3" entrytime="00:01:00.00" entrycourse="LCM" />
                <RESULT eventid="98830" points="494" reactiontime="+91" swimtime="00:02:24.14" resultid="101212" heatid="105158" lane="0" entrytime="00:02:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                    <SPLIT distance="100" swimtime="00:01:09.29" />
                    <SPLIT distance="150" swimtime="00:01:49.66" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="98956" points="451" reactiontime="+88" swimtime="00:02:45.52" resultid="101213" heatid="105199" lane="9" entrytime="00:03:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.58" />
                    <SPLIT distance="100" swimtime="00:01:18.00" />
                    <SPLIT distance="150" swimtime="00:02:01.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="485" reactiontime="+93" swimtime="00:00:59.67" resultid="101214" heatid="105227" lane="1" entrytime="00:00:58.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="101215" heatid="105249" lane="2" entrytime="00:02:00.00" entrycourse="LCM" />
                <RESULT eventid="99218" points="500" reactiontime="+76" swimtime="00:02:08.44" resultid="101216" heatid="105305" lane="7" entrytime="00:02:08.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.28" />
                    <SPLIT distance="100" swimtime="00:01:02.55" />
                    <SPLIT distance="150" swimtime="00:01:35.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="101217" heatid="105351" lane="7" entrytime="00:01:00.00" entrycourse="LCM" />
                <RESULT eventid="99473" points="508" reactiontime="+76" swimtime="00:04:35.63" resultid="101218" heatid="106059" lane="8" entrytime="00:04:35.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.04" />
                    <SPLIT distance="100" swimtime="00:01:04.49" />
                    <SPLIT distance="150" swimtime="00:01:39.10" />
                    <SPLIT distance="200" swimtime="00:02:14.19" />
                    <SPLIT distance="250" swimtime="00:02:49.42" />
                    <SPLIT distance="300" swimtime="00:03:24.95" />
                    <SPLIT distance="350" swimtime="00:04:00.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-09-29" firstname="Radosław" gender="M" lastname="STĘPIEŃ" nation="POL" swrid="4992764" athleteid="101219">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="101220" heatid="105137" lane="9" entrytime="00:00:28.70" entrycourse="LCM" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="101221" heatid="105221" lane="2" entrytime="00:01:07.00" entrycourse="LCM" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="101222" heatid="105357" lane="7" entrytime="00:00:39.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-07-27" firstname="Natalia" gender="F" lastname="SZCZĘSNOWICZ" nation="POL" swrid="4992766" athleteid="101223">
              <RESULTS>
                <RESULT eventid="98777" status="DNS" swimtime="00:00:00.00" resultid="101224" heatid="105118" lane="5" entrytime="00:00:32.88" entrycourse="SCM" />
                <RESULT eventid="98972" status="DNS" swimtime="00:00:00.00" resultid="101225" heatid="105210" lane="3" entrytime="00:01:12.00" entrycourse="LCM" />
                <RESULT eventid="99154" status="DNS" swimtime="00:00:00.00" resultid="101226" heatid="105262" lane="9" entrytime="00:00:37.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-05-13" firstname="Łukasz" gender="M" lastname="KLEKOT" nation="POL" swrid="4071663" athleteid="101227">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="101228" heatid="105140" lane="2" entrytime="00:00:27.00" entrycourse="LCM" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="101229" heatid="105228" lane="9" entrytime="00:00:57.00" entrycourse="LCM" />
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="101230" heatid="105305" lane="1" entrytime="00:02:08.00" entrycourse="LCM" />
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="101231" entrytime="00:04:40.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="OCSUC" nation="POL" region="WIE" clubid="105087" name="4SM Octopus Suchy Las">
          <CONTACT city="Suchy Las" email="uksoctopus.suchylas@gmail.com" name="Łukasz Kolendowicz" phone="608098108" state="WLKP" street="Szkolna 18" zip="62-002" />
          <ATHLETES>
            <ATHLETE birthdate="1988-05-16" firstname="Łukasz" gender="M" lastname="KOLENDOWICZ" nation="POL" athleteid="105088">
              <RESULTS>
                <RESULT eventid="98891" points="460" swimtime="00:18:48.32" resultid="105089" heatid="105420" lane="5" entrytime="00:18:40.00" />
                <RESULT eventid="98924" points="520" reactiontime="+70" swimtime="00:00:29.89" resultid="105090" heatid="105190" lane="6" entrytime="00:00:29.00" />
                <RESULT eventid="99186" points="489" reactiontime="+78" swimtime="00:01:05.92" resultid="105091" heatid="105288" lane="5" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" status="DNS" swimtime="00:00:00.00" resultid="105092" heatid="106053" lane="5" entrytime="00:05:10.00" />
                <RESULT eventid="99473" points="514" reactiontime="+90" swimtime="00:04:34.64" resultid="105093" heatid="106059" lane="5" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                    <SPLIT distance="100" swimtime="00:01:03.19" />
                    <SPLIT distance="150" swimtime="00:01:37.49" />
                    <SPLIT distance="200" swimtime="00:02:12.30" />
                    <SPLIT distance="250" swimtime="00:02:47.78" />
                    <SPLIT distance="300" swimtime="00:03:23.93" />
                    <SPLIT distance="350" swimtime="00:04:00.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="ŚL" clubid="100553" name="AZS PWSZ Racibórz">
          <CONTACT city="Racibórz" email="adip45@poczta.onet.pl" name="kunicki marcin" phone="606 114286" state="ŚL" street="słowackiego 55" zip="47-400" />
          <ATHLETES>
            <ATHLETE birthdate="1957-04-11" firstname="Adolf" gender="M" lastname="PIECHULA" nation="POL" swrid="4992724" athleteid="100554">
              <RESULTS>
                <RESULT eventid="98830" points="244" reactiontime="+81" swimtime="00:03:02.23" resultid="100555" heatid="105152" lane="6" entrytime="00:03:01.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                    <SPLIT distance="100" swimtime="00:01:24.77" />
                    <SPLIT distance="150" swimtime="00:02:18.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="246" reactiontime="+84" swimtime="00:03:22.44" resultid="100556" heatid="105201" lane="9" entrytime="00:03:11.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.48" />
                    <SPLIT distance="100" swimtime="00:01:36.24" />
                    <SPLIT distance="150" swimtime="00:02:29.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="194" reactiontime="+102" swimtime="00:03:12.51" resultid="100557" heatid="105234" lane="3" entrytime="00:03:09.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.26" />
                    <SPLIT distance="100" swimtime="00:01:32.23" />
                    <SPLIT distance="150" swimtime="00:02:23.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="267" reactiontime="+85" swimtime="00:01:30.68" resultid="100558" heatid="105253" lane="7" entrytime="00:01:27.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="231" reactiontime="+94" swimtime="00:06:37.14" resultid="100559" heatid="106051" lane="8" entrytime="00:06:28.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.30" />
                    <SPLIT distance="100" swimtime="00:01:35.75" />
                    <SPLIT distance="150" swimtime="00:02:27.51" />
                    <SPLIT distance="200" swimtime="00:03:18.29" />
                    <SPLIT distance="250" swimtime="00:04:13.63" />
                    <SPLIT distance="300" swimtime="00:05:08.65" />
                    <SPLIT distance="350" swimtime="00:05:53.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="200" reactiontime="+90" swimtime="00:01:25.17" resultid="100560" heatid="105328" lane="8" entrytime="00:01:23.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="293" reactiontime="+81" swimtime="00:00:40.12" resultid="100561" heatid="105358" lane="0" entrytime="00:00:37.89" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="102933" name="AZS UW Warszawa">
          <ATHLETES>
            <ATHLETE birthdate="1992-02-14" firstname="Hubert" gender="M" lastname="BIGDOWSKI" nation="POL" swrid="4992714" athleteid="102934">
              <RESULTS>
                <RESULT eventid="98798" points="481" reactiontime="+81" swimtime="00:00:26.67" resultid="103028" heatid="105143" lane="4" entrytime="00:00:22.50" />
                <RESULT eventid="98988" points="433" reactiontime="+90" swimtime="00:01:01.99" resultid="103029" heatid="105226" lane="4" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="446" reactiontime="+89" swimtime="00:00:29.34" resultid="103030" heatid="105273" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="103031" heatid="105302" lane="6" entrytime="00:02:20.00" />
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="103032" heatid="105330" lane="9" entrytime="00:01:10.00" />
                <RESULT eventid="99425" points="437" reactiontime="+81" swimtime="00:00:35.13" resultid="103033" heatid="105361" lane="6" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="103481" name="AZS UWM Masters Olsztyn" shortname="AZS UWM Mrs Olsztyn">
          <CONTACT email="gozdzik@uwm.edu.pl" name="Goździejewska Anna" phone="501372846" />
          <ATHLETES>
            <ATHLETE birthdate="1965-02-14" firstname="Dariusz" gender="M" lastname="POZIEMSKI" nation="POL" athleteid="103489">
              <RESULTS>
                <RESULT eventid="98924" points="341" reactiontime="+74" swimtime="00:00:34.39" resultid="103490" heatid="105188" lane="9" entrytime="00:00:33.00" />
                <RESULT eventid="99170" points="351" reactiontime="+68" swimtime="00:00:31.79" resultid="103491" heatid="105274" lane="9" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-03-18" firstname="Anna" gender="F" lastname="GOŹDZIEJEWSKA" nation="POL" swrid="4313183" athleteid="103492">
              <RESULTS>
                <RESULT eventid="98814" points="281" reactiontime="+82" swimtime="00:03:12.54" resultid="103493" heatid="105145" lane="7" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.83" />
                    <SPLIT distance="100" swimtime="00:01:34.13" />
                    <SPLIT distance="150" swimtime="00:02:29.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98863" points="320" swimtime="00:12:01.46" resultid="103494" heatid="105405" lane="5" entrytime="00:12:00.00" />
                <RESULT eventid="98940" points="274" swimtime="00:03:34.00" resultid="103495" heatid="105193" lane="7" entrytime="00:03:30.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.63" />
                    <SPLIT distance="100" swimtime="00:01:44.94" />
                    <SPLIT distance="150" swimtime="00:02:39.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="343" reactiontime="+96" swimtime="00:01:14.37" resultid="103496" heatid="105209" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="306" swimtime="00:02:47.60" resultid="103497" heatid="105292" lane="1" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.03" />
                    <SPLIT distance="100" swimtime="00:01:21.92" />
                    <SPLIT distance="150" swimtime="00:02:05.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" points="278" reactiontime="+101" swimtime="00:06:50.85" resultid="103498" heatid="106046" lane="6" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.54" />
                    <SPLIT distance="100" swimtime="00:01:45.44" />
                    <SPLIT distance="150" swimtime="00:02:40.26" />
                    <SPLIT distance="200" swimtime="00:03:33.24" />
                    <SPLIT distance="250" swimtime="00:04:28.58" />
                    <SPLIT distance="300" swimtime="00:05:23.78" />
                    <SPLIT distance="350" swimtime="00:06:08.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="248" reactiontime="+88" swimtime="00:00:46.90" resultid="103499" heatid="105346" lane="5" entrytime="00:00:45.80" />
                <RESULT eventid="99457" points="312" swimtime="00:05:52.25" resultid="103500" heatid="106055" lane="8" entrytime="00:05:55.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.18" />
                    <SPLIT distance="100" swimtime="00:01:24.24" />
                    <SPLIT distance="150" swimtime="00:02:09.42" />
                    <SPLIT distance="200" swimtime="00:02:54.70" />
                    <SPLIT distance="250" swimtime="00:03:39.58" />
                    <SPLIT distance="300" swimtime="00:04:24.37" />
                    <SPLIT distance="350" swimtime="00:05:09.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-01-29" firstname="Mariusz" gender="M" lastname="GABIEC" nation="POL" swrid="4754711" athleteid="103501">
              <RESULTS>
                <RESULT eventid="98798" points="377" reactiontime="+95" swimtime="00:00:28.94" resultid="103502" heatid="105123" lane="1" />
                <RESULT eventid="98830" points="342" reactiontime="+99" swimtime="00:02:43.01" resultid="103503" heatid="105155" lane="0" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                    <SPLIT distance="100" swimtime="00:01:15.50" />
                    <SPLIT distance="150" swimtime="00:02:05.46" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="98924" points="356" reactiontime="+137" swimtime="00:00:33.90" resultid="103504" heatid="105180" lane="2" />
                <RESULT eventid="98988" points="383" reactiontime="+82" swimtime="00:01:04.57" resultid="103505" heatid="105222" lane="8" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="367" reactiontime="+91" swimtime="00:02:22.43" resultid="103506" heatid="105300" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                    <SPLIT distance="100" swimtime="00:01:10.24" />
                    <SPLIT distance="150" swimtime="00:01:46.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="294" reactiontime="+85" swimtime="00:02:48.27" resultid="103507" heatid="105335" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.58" />
                    <SPLIT distance="100" swimtime="00:01:22.49" />
                    <SPLIT distance="150" swimtime="00:02:05.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="367" reactiontime="+90" swimtime="00:05:07.24" resultid="103508" heatid="106063" lane="2" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                    <SPLIT distance="100" swimtime="00:01:14.57" />
                    <SPLIT distance="150" swimtime="00:01:53.67" />
                    <SPLIT distance="200" swimtime="00:02:32.93" />
                    <SPLIT distance="250" swimtime="00:03:12.37" />
                    <SPLIT distance="300" swimtime="00:03:52.05" />
                    <SPLIT distance="350" swimtime="00:04:31.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-30" firstname="Paweł" gender="M" lastname="GREGOROWICZ" nation="POL" swrid="4992729" athleteid="103509">
              <RESULTS>
                <RESULT eventid="98798" points="477" reactiontime="+79" swimtime="00:00:26.76" resultid="103510" heatid="105127" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="98830" points="419" reactiontime="+72" swimtime="00:02:32.27" resultid="103511" heatid="105156" lane="8" entrytime="00:02:36.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.51" />
                    <SPLIT distance="100" swimtime="00:01:12.49" />
                    <SPLIT distance="150" swimtime="00:01:57.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="505" reactiontime="+74" swimtime="00:00:58.87" resultid="103512" heatid="105226" lane="9" entrytime="00:00:59.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="462" reactiontime="+88" swimtime="00:00:29.00" resultid="103513" heatid="105274" lane="2" entrytime="00:00:29.04" />
                <RESULT eventid="99218" points="452" reactiontime="+88" swimtime="00:02:12.82" resultid="103514" heatid="105304" lane="1" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.80" />
                    <SPLIT distance="100" swimtime="00:01:04.66" />
                    <SPLIT distance="150" swimtime="00:01:39.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="439" reactiontime="+87" swimtime="00:01:05.55" resultid="103515" heatid="105329" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="410" reactiontime="+88" swimtime="00:04:56.05" resultid="103516" heatid="106062" lane="5" entrytime="00:05:05.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                    <SPLIT distance="100" swimtime="00:01:11.80" />
                    <SPLIT distance="150" swimtime="00:01:50.35" />
                    <SPLIT distance="200" swimtime="00:02:28.68" />
                    <SPLIT distance="250" swimtime="00:03:06.40" />
                    <SPLIT distance="300" swimtime="00:03:44.27" />
                    <SPLIT distance="350" swimtime="00:04:21.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-02-15" firstname="Jowita" gender="F" lastname="KUCHARSKA" nation="POL" swrid="4313184" athleteid="103517">
              <RESULTS>
                <RESULT eventid="98777" points="407" reactiontime="+88" swimtime="00:00:32.01" resultid="103518" heatid="105119" lane="2" entrytime="00:00:31.79" entrycourse="SCM" />
                <RESULT eventid="98907" points="316" reactiontime="+87" swimtime="00:00:39.71" resultid="103519" heatid="105176" lane="3" entrytime="00:00:39.00" />
                <RESULT eventid="99314" points="326" reactiontime="+77" swimtime="00:01:24.44" resultid="103520" heatid="105279" lane="6" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="290" reactiontime="+90" swimtime="00:03:07.32" resultid="103521" heatid="105334" lane="1" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.41" />
                    <SPLIT distance="100" swimtime="00:01:31.91" />
                    <SPLIT distance="150" swimtime="00:02:20.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="367" reactiontime="+110" swimtime="00:00:35.01" resultid="105084" heatid="105262" lane="4" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-26" firstname="Aleksandra" gender="F" lastname="PRZYBYSZ" nation="POL" swrid="4992725" athleteid="103522">
              <RESULTS>
                <RESULT eventid="98863" points="295" swimtime="00:12:21.10" resultid="103523" heatid="105405" lane="2" entrytime="00:12:20.00" />
                <RESULT eventid="98972" status="DNS" swimtime="00:00:00.00" resultid="103524" heatid="105208" lane="7" entrytime="00:01:19.00" />
                <RESULT eventid="99004" points="201" reactiontime="+108" swimtime="00:03:27.86" resultid="103525" heatid="105230" lane="7" entrytime="00:03:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.22" />
                    <SPLIT distance="100" swimtime="00:01:39.73" />
                    <SPLIT distance="150" swimtime="00:02:34.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="232" reactiontime="+106" swimtime="00:00:40.75" resultid="103526" heatid="105260" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="99202" points="295" reactiontime="+103" swimtime="00:02:49.59" resultid="103527" heatid="105292" lane="0" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                    <SPLIT distance="100" swimtime="00:01:23.57" />
                    <SPLIT distance="150" swimtime="00:02:07.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="211" reactiontime="+106" swimtime="00:01:33.94" resultid="103528" heatid="105322" lane="1" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="285" reactiontime="+104" swimtime="00:06:03.00" resultid="103529" heatid="106056" lane="5" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.43" />
                    <SPLIT distance="100" swimtime="00:01:28.97" />
                    <SPLIT distance="150" swimtime="00:02:15.74" />
                    <SPLIT distance="200" swimtime="00:03:02.48" />
                    <SPLIT distance="250" swimtime="00:03:49.45" />
                    <SPLIT distance="300" swimtime="00:04:35.48" />
                    <SPLIT distance="350" swimtime="00:05:21.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-08-01" firstname="Małgorzata" gender="F" lastname="POLITO" nation="POL" athleteid="103530">
              <RESULTS>
                <RESULT eventid="98863" points="310" swimtime="00:12:09.62" resultid="103531" heatid="105405" lane="6" entrytime="00:12:20.00" />
                <RESULT eventid="98940" points="345" reactiontime="+86" swimtime="00:03:18.25" resultid="103532" heatid="105193" lane="5" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.78" />
                    <SPLIT distance="100" swimtime="00:01:37.11" />
                    <SPLIT distance="150" swimtime="00:02:28.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="333" reactiontime="+86" swimtime="00:01:32.83" resultid="103533" heatid="105246" lane="5" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="311" reactiontime="+94" swimtime="00:02:46.66" resultid="103534" heatid="105292" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.96" />
                    <SPLIT distance="100" swimtime="00:01:21.60" />
                    <SPLIT distance="150" swimtime="00:02:05.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="307" reactiontime="+99" swimtime="00:05:54.45" resultid="103535" heatid="106055" lane="2" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.49" />
                    <SPLIT distance="100" swimtime="00:01:24.92" />
                    <SPLIT distance="150" swimtime="00:02:10.63" />
                    <SPLIT distance="200" swimtime="00:02:57.16" />
                    <SPLIT distance="250" swimtime="00:03:42.17" />
                    <SPLIT distance="300" swimtime="00:04:28.14" />
                    <SPLIT distance="350" swimtime="00:05:13.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="335" reactiontime="+87" swimtime="00:00:42.42" resultid="105094" heatid="105348" lane="3" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-13" firstname="Michał" gender="M" lastname="KOZIKOWSKI" nation="POL" swrid="4992728" athleteid="103536">
              <RESULTS>
                <RESULT eventid="98830" points="417" reactiontime="+81" swimtime="00:02:32.53" resultid="103537" heatid="105155" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                    <SPLIT distance="100" swimtime="00:01:12.78" />
                    <SPLIT distance="150" swimtime="00:01:55.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="459" reactiontime="+86" swimtime="00:02:44.65" resultid="103538" heatid="105204" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.62" />
                    <SPLIT distance="100" swimtime="00:01:17.20" />
                    <SPLIT distance="150" swimtime="00:01:59.89" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="04" eventid="99091" reactiontime="+67" status="DSQ" swimtime="00:00:00.00" resultid="103539" heatid="105257" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="354" reactiontime="+88" swimtime="00:05:44.49" resultid="103540" heatid="106052" lane="3" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                    <SPLIT distance="100" swimtime="00:01:24.92" />
                    <SPLIT distance="150" swimtime="00:02:10.57" />
                    <SPLIT distance="200" swimtime="00:02:54.47" />
                    <SPLIT distance="250" swimtime="00:03:39.73" />
                    <SPLIT distance="300" swimtime="00:04:24.35" />
                    <SPLIT distance="350" swimtime="00:05:06.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="459" reactiontime="+87" swimtime="00:00:34.56" resultid="103541" heatid="105361" lane="3" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-09-01" firstname="Marek" gender="M" lastname="KOŹLIKOWSKI" nation="POL" swrid="4992727" athleteid="103542">
              <RESULTS>
                <RESULT eventid="98830" points="230" reactiontime="+99" swimtime="00:03:06.06" resultid="103543" heatid="105151" lane="1" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                    <SPLIT distance="100" swimtime="00:01:31.28" />
                    <SPLIT distance="150" swimtime="00:02:24.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="275" reactiontime="+92" swimtime="00:01:12.11" resultid="103544" heatid="105216" lane="9" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="192" reactiontime="+97" swimtime="00:07:02.10" resultid="103545" heatid="106049" lane="6" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.70" />
                    <SPLIT distance="100" swimtime="00:01:41.96" />
                    <SPLIT distance="150" swimtime="00:02:41.04" />
                    <SPLIT distance="200" swimtime="00:03:39.65" />
                    <SPLIT distance="250" swimtime="00:04:34.69" />
                    <SPLIT distance="300" swimtime="00:05:30.94" />
                    <SPLIT distance="350" swimtime="00:06:16.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="221" reactiontime="+108" swimtime="00:06:03.80" resultid="103546" heatid="106065" lane="1" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.74" />
                    <SPLIT distance="100" swimtime="00:01:23.71" />
                    <SPLIT distance="150" swimtime="00:02:10.23" />
                    <SPLIT distance="200" swimtime="00:02:57.88" />
                    <SPLIT distance="250" swimtime="00:03:45.53" />
                    <SPLIT distance="300" swimtime="00:04:33.00" />
                    <SPLIT distance="350" swimtime="00:05:19.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-12-31" firstname="Marek" gender="M" lastname="HASSO-AGOPSOWICZ" nation="POL" athleteid="103547">
              <RESULTS>
                <RESULT eventid="98798" points="126" reactiontime="+108" swimtime="00:00:41.65" resultid="103548" heatid="105124" lane="6" entrytime="00:00:42.00" />
                <RESULT eventid="98988" points="104" reactiontime="+108" swimtime="00:01:39.58" resultid="103550" heatid="105213" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="78" reactiontime="+109" swimtime="00:03:58.41" resultid="103551" heatid="105295" lane="6" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.16" />
                    <SPLIT distance="100" swimtime="00:01:49.78" />
                    <SPLIT distance="150" swimtime="00:02:56.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="72" reactiontime="+115" swimtime="00:08:48.03" resultid="103552" heatid="106066" lane="9" entrytime="00:08:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.04" />
                    <SPLIT distance="100" swimtime="00:01:56.73" />
                    <SPLIT distance="150" swimtime="00:03:04.04" />
                    <SPLIT distance="200" swimtime="00:04:14.42" />
                    <SPLIT distance="250" swimtime="00:05:23.65" />
                    <SPLIT distance="300" swimtime="00:06:35.44" />
                    <SPLIT distance="350" swimtime="00:07:46.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-06-10" firstname="Dariusz" gender="M" lastname="ONICHIMOWSKI" nation="POL" athleteid="103553">
              <RESULTS>
                <RESULT eventid="98798" points="270" reactiontime="+96" swimtime="00:00:32.34" resultid="103554" heatid="105130" lane="8" entrytime="00:00:32.00" />
                <RESULT eventid="98924" points="236" reactiontime="+67" swimtime="00:00:38.88" resultid="103555" heatid="105185" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="99186" points="48" reactiontime="+125" swimtime="00:02:22.03" resultid="103556" heatid="105281" lane="9" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="240" reactiontime="+80" swimtime="00:00:42.86" resultid="103557" heatid="105357" lane="9" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-17" firstname="Anna" gender="F" lastname="PIEKUT" nation="POL" swrid="4072764" athleteid="103558">
              <RESULTS>
                <RESULT eventid="98814" points="365" reactiontime="+89" swimtime="00:02:56.39" resultid="103559" heatid="105147" lane="0" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.37" />
                    <SPLIT distance="100" swimtime="00:01:20.55" />
                    <SPLIT distance="150" swimtime="00:02:13.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="288" reactiontime="+78" swimtime="00:03:30.53" resultid="103560" heatid="105191" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.49" />
                    <SPLIT distance="100" swimtime="00:01:41.94" />
                    <SPLIT distance="150" swimtime="00:02:36.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99004" points="388" reactiontime="+84" swimtime="00:02:46.89" resultid="103561" heatid="105230" lane="5" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                    <SPLIT distance="100" swimtime="00:01:20.30" />
                    <SPLIT distance="150" swimtime="00:02:03.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="387" swimtime="00:00:34.40" resultid="103562" heatid="105263" lane="7" entrytime="00:00:34.05" />
                <RESULT eventid="99266" points="379" reactiontime="+90" swimtime="00:06:10.65" resultid="103563" heatid="106046" lane="4" entrytime="00:06:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.14" />
                    <SPLIT distance="100" swimtime="00:01:20.87" />
                    <SPLIT distance="150" swimtime="00:02:11.36" />
                    <SPLIT distance="200" swimtime="00:02:59.92" />
                    <SPLIT distance="250" swimtime="00:03:52.32" />
                    <SPLIT distance="300" swimtime="00:04:45.47" />
                    <SPLIT distance="350" swimtime="00:05:28.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="381" reactiontime="+88" swimtime="00:01:17.16" resultid="103564" heatid="105323" lane="2" entrytime="00:01:15.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="295" reactiontime="+85" swimtime="00:00:44.26" resultid="103565" heatid="105348" lane="0" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-09-01" firstname="Grzegorz" gender="M" lastname="MÓWIŃSKI" nation="POL" swrid="4992726" athleteid="103566">
              <RESULTS>
                <RESULT eventid="98891" status="WDR" swimtime="00:00:00.00" resultid="103567" entrytime="00:24:00.00" />
                <RESULT eventid="99020" points="192" reactiontime="+89" swimtime="00:03:13.05" resultid="103568" heatid="105234" lane="9" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.36" />
                    <SPLIT distance="100" swimtime="00:01:32.17" />
                    <SPLIT distance="150" swimtime="00:02:24.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="210" reactiontime="+79" swimtime="00:02:51.55" resultid="103569" heatid="105298" lane="8" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.42" />
                    <SPLIT distance="100" swimtime="00:01:23.48" />
                    <SPLIT distance="150" swimtime="00:02:08.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="212" reactiontime="+91" swimtime="00:01:23.55" resultid="103570" heatid="105327" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="209" reactiontime="+86" swimtime="00:06:10.72" resultid="103571" heatid="106064" lane="8" entrytime="00:06:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.82" />
                    <SPLIT distance="100" swimtime="00:01:25.91" />
                    <SPLIT distance="150" swimtime="00:02:13.29" />
                    <SPLIT distance="200" swimtime="00:03:01.02" />
                    <SPLIT distance="250" swimtime="00:03:49.69" />
                    <SPLIT distance="300" swimtime="00:04:37.77" />
                    <SPLIT distance="350" swimtime="00:05:25.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-11-25" firstname="Piotr" gender="M" lastname="MARKOWICZ" nation="POL" swrid="4992730" athleteid="103572">
              <RESULTS>
                <RESULT eventid="98798" points="340" reactiontime="+88" swimtime="00:00:29.95" resultid="103573" heatid="105131" lane="6" entrytime="00:00:31.20" />
                <RESULT eventid="98830" points="332" reactiontime="+102" swimtime="00:02:44.62" resultid="103574" heatid="105154" lane="1" entrytime="00:02:51.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.93" />
                    <SPLIT distance="100" swimtime="00:01:17.84" />
                    <SPLIT distance="150" swimtime="00:02:05.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="301" reactiontime="+73" swimtime="00:00:35.85" resultid="103575" heatid="105186" lane="7" entrytime="00:00:36.00" />
                <RESULT eventid="98988" points="361" reactiontime="+83" swimtime="00:01:05.86" resultid="103576" heatid="105218" lane="7" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" status="DNS" swimtime="00:00:00.00" resultid="103577" heatid="105284" lane="4" entrytime="00:01:18.70" />
                <RESULT eventid="99282" points="292" reactiontime="+92" swimtime="00:06:07.43" resultid="103578" heatid="106051" lane="6" entrytime="00:06:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.58" />
                    <SPLIT distance="100" swimtime="00:01:20.18" />
                    <SPLIT distance="150" swimtime="00:02:08.26" />
                    <SPLIT distance="200" swimtime="00:02:56.31" />
                    <SPLIT distance="250" swimtime="00:03:51.39" />
                    <SPLIT distance="300" swimtime="00:04:46.31" />
                    <SPLIT distance="350" swimtime="00:05:27.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="258" reactiontime="+77" swimtime="00:02:55.60" resultid="103579" heatid="105340" lane="7" entrytime="00:02:51.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.44" />
                    <SPLIT distance="100" swimtime="00:01:25.75" />
                    <SPLIT distance="150" swimtime="00:02:11.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="301" reactiontime="+88" swimtime="00:05:28.02" resultid="103580" heatid="106062" lane="9" entrytime="00:05:25.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                    <SPLIT distance="100" swimtime="00:01:18.65" />
                    <SPLIT distance="150" swimtime="00:02:00.87" />
                    <SPLIT distance="200" swimtime="00:02:43.66" />
                    <SPLIT distance="250" swimtime="00:03:26.02" />
                    <SPLIT distance="300" swimtime="00:04:08.33" />
                    <SPLIT distance="350" swimtime="00:04:49.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-09-30" firstname="Karol" gender="M" lastname="DZIEMIAN" nation="POL" athleteid="103581">
              <RESULTS>
                <RESULT eventid="98798" points="211" reactiontime="+96" swimtime="00:00:35.09" resultid="103582" heatid="105128" lane="0" entrytime="00:00:34.88" />
                <RESULT eventid="98988" points="211" reactiontime="+114" swimtime="00:01:18.73" resultid="103583" heatid="105215" lane="3" entrytime="00:01:20.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="165" reactiontime="+117" swimtime="00:03:05.95" resultid="103584" heatid="105297" lane="0" entrytime="00:03:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.01" />
                    <SPLIT distance="100" swimtime="00:01:30.12" />
                    <SPLIT distance="150" swimtime="00:02:20.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-09-21" firstname="Tomasz" gender="M" lastname="KOZŁOWSKI" nation="POL" athleteid="103585">
              <RESULTS>
                <RESULT eventid="98956" points="153" reactiontime="+96" swimtime="00:03:56.96" resultid="103586" heatid="105200" lane="5" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.26" />
                    <SPLIT distance="100" swimtime="00:01:55.09" />
                    <SPLIT distance="150" swimtime="00:02:57.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="164" reactiontime="+76" swimtime="00:01:46.79" resultid="103587" heatid="105252" lane="8" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="159" reactiontime="+107" swimtime="00:00:49.21" resultid="103588" heatid="105354" lane="4" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-04-24" firstname="Przemysław" gender="M" lastname="BIELSKI" nation="POL" athleteid="103589">
              <RESULTS>
                <RESULT eventid="98798" points="316" reactiontime="+93" swimtime="00:00:30.67" resultid="103590" heatid="105130" lane="9" entrytime="00:00:32.40" />
                <RESULT eventid="98988" points="344" reactiontime="+103" swimtime="00:01:06.89" resultid="103591" heatid="105220" lane="2" entrytime="00:01:08.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="274" reactiontime="+120" swimtime="00:00:34.50" resultid="103592" heatid="105269" lane="1" entrytime="00:00:35.40" />
                <RESULT eventid="99218" points="294" reactiontime="+113" swimtime="00:02:33.26" resultid="103593" heatid="105298" lane="1" entrytime="00:02:50.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                    <SPLIT distance="100" swimtime="00:01:12.04" />
                    <SPLIT distance="150" swimtime="00:01:52.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="273" reactiontime="+103" swimtime="00:05:39.05" resultid="103594" heatid="106064" lane="7" entrytime="00:06:01.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                    <SPLIT distance="100" swimtime="00:01:15.84" />
                    <SPLIT distance="150" swimtime="00:01:58.42" />
                    <SPLIT distance="200" swimtime="00:02:42.13" />
                    <SPLIT distance="250" swimtime="00:03:26.57" />
                    <SPLIT distance="300" swimtime="00:04:11.28" />
                    <SPLIT distance="350" swimtime="00:04:56.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-03-04" firstname="Tomasz" gender="M" lastname="KLAMRA" nation="POL" athleteid="103595">
              <RESULTS>
                <RESULT eventid="98830" points="173" reactiontime="+98" swimtime="00:03:24.27" resultid="103596" heatid="105148" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.66" />
                    <SPLIT distance="100" swimtime="00:01:30.76" />
                    <SPLIT distance="150" swimtime="00:02:36.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="167" reactiontime="+77" swimtime="00:00:43.62" resultid="103597" heatid="105185" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="99170" points="217" reactiontime="+83" swimtime="00:00:37.28" resultid="103598" heatid="105269" lane="9" entrytime="00:00:35.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-05-30" firstname="Piotr" gender="M" lastname="KOZŁOWSKI" nation="POL" athleteid="103599">
              <RESULTS>
                <RESULT eventid="98956" status="DNS" swimtime="00:00:00.00" resultid="103600" heatid="105202" lane="9" entrytime="00:03:05.00" />
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="103601" heatid="105256" lane="0" entrytime="00:01:21.00" />
                <RESULT eventid="99425" points="356" reactiontime="+77" swimtime="00:00:37.63" resultid="103602" heatid="105358" lane="8" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-03-26" firstname="Grzegorz" gender="M" lastname="KALINOWSKI" nation="POL" athleteid="103603">
              <RESULTS>
                <RESULT eventid="98798" points="307" reactiontime="+70" swimtime="00:00:30.97" resultid="103604" heatid="105129" lane="8" entrytime="00:00:33.00" />
                <RESULT eventid="98924" points="223" reactiontime="+75" swimtime="00:00:39.60" resultid="103605" heatid="105185" lane="8" entrytime="00:00:39.00" />
                <RESULT eventid="98988" points="299" reactiontime="+84" swimtime="00:01:10.10" resultid="103606" heatid="105219" lane="5" entrytime="00:01:09.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-21" firstname="Monika" gender="F" lastname="CHODYNA" nation="POL" swrid="4072155" athleteid="103607">
              <RESULTS>
                <RESULT eventid="98777" points="561" reactiontime="+79" swimtime="00:00:28.76" resultid="103609" heatid="105121" lane="6" entrytime="00:00:28.80" entrycourse="LCM" />
                <RESULT eventid="98972" points="572" reactiontime="+86" swimtime="00:01:02.71" resultid="103610" heatid="105212" lane="2" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="566" reactiontime="+83" swimtime="00:02:16.52" resultid="103611" heatid="105294" lane="4" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                    <SPLIT distance="100" swimtime="00:01:05.88" />
                    <SPLIT distance="150" swimtime="00:01:41.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="566" reactiontime="+82" swimtime="00:04:48.99" resultid="103612" heatid="106054" lane="4" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                    <SPLIT distance="100" swimtime="00:01:08.54" />
                    <SPLIT distance="150" swimtime="00:01:45.37" />
                    <SPLIT distance="200" swimtime="00:02:22.53" />
                    <SPLIT distance="250" swimtime="00:03:00.12" />
                    <SPLIT distance="300" swimtime="00:03:37.79" />
                    <SPLIT distance="350" swimtime="00:04:14.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98863" points="548" reactiontime="+86" swimtime="00:10:03.41" resultid="103613" heatid="105404" lane="4" entrytime="00:09:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                    <SPLIT distance="100" swimtime="00:01:09.63" />
                    <SPLIT distance="150" swimtime="00:01:47.31" />
                    <SPLIT distance="200" swimtime="00:02:24.83" />
                    <SPLIT distance="250" swimtime="00:03:02.49" />
                    <SPLIT distance="300" swimtime="00:03:40.38" />
                    <SPLIT distance="350" swimtime="00:04:18.62" />
                    <SPLIT distance="400" swimtime="00:04:56.85" />
                    <SPLIT distance="450" swimtime="00:05:35.14" />
                    <SPLIT distance="500" swimtime="00:06:13.61" />
                    <SPLIT distance="550" swimtime="00:06:52.49" />
                    <SPLIT distance="600" swimtime="00:07:31.50" />
                    <SPLIT distance="650" swimtime="00:08:09.79" />
                    <SPLIT distance="700" swimtime="00:08:48.46" />
                    <SPLIT distance="750" swimtime="00:09:26.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="502" reactiontime="+81" swimtime="00:00:31.53" resultid="103614" heatid="105264" lane="5" entrytime="00:00:30.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-11-25" firstname="Janusz" gender="M" lastname="CHODYNA" nation="POL" athleteid="103608">
              <RESULTS>
                <RESULT eventid="99425" points="409" reactiontime="+75" swimtime="00:00:35.92" resultid="103615" heatid="105361" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="99091" points="357" reactiontime="+77" swimtime="00:01:22.35" resultid="103616" heatid="105255" lane="3" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" status="DNS" swimtime="00:00:00.00" resultid="103617" heatid="105202" lane="0" entrytime="00:03:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-09-29" firstname="Jakub" gender="M" lastname="STĘPIEŃ" nation="POL" athleteid="104371">
              <RESULTS>
                <RESULT eventid="98798" points="327" reactiontime="+78" swimtime="00:00:30.33" resultid="104372" heatid="105136" lane="7" entrytime="00:00:29.00" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="104373" heatid="105219" lane="6" entrytime="00:01:10.00" />
                <RESULT comment="04" eventid="99473" reactiontime="+77" status="DSQ" swimtime="00:00:00.00" resultid="105391" heatid="106063" lane="6" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.70" />
                    <SPLIT distance="100" swimtime="00:01:16.84" />
                    <SPLIT distance="150" swimtime="00:02:01.47" />
                    <SPLIT distance="200" swimtime="00:02:48.49" />
                    <SPLIT distance="250" swimtime="00:03:35.50" />
                    <SPLIT distance="300" swimtime="00:04:22.25" />
                    <SPLIT distance="350" swimtime="00:05:09.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99059" points="356" reactiontime="+85" swimtime="00:02:11.79" resultid="104100" heatid="105241" lane="7" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.51" />
                    <SPLIT distance="100" swimtime="00:01:12.41" />
                    <SPLIT distance="150" swimtime="00:01:41.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103501" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="103509" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="103608" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="103603" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99250" points="387" reactiontime="+97" swimtime="00:01:56.43" resultid="104104" heatid="105310" lane="2" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                    <SPLIT distance="100" swimtime="00:01:00.49" />
                    <SPLIT distance="150" swimtime="00:01:27.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103603" number="1" reactiontime="+97" />
                    <RELAYPOSITION athleteid="103489" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="103509" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="103501" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="99059" points="288" reactiontime="+78" swimtime="00:02:21.36" resultid="104101" heatid="105241" lane="9" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.67" />
                    <SPLIT distance="100" swimtime="00:01:10.64" />
                    <SPLIT distance="150" swimtime="00:01:46.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103572" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="103536" number="2" />
                    <RELAYPOSITION athleteid="103595" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="103599" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="99250" points="398" reactiontime="+87" swimtime="00:01:55.34" resultid="104105" heatid="105310" lane="9" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.08" />
                    <SPLIT distance="100" swimtime="00:00:58.28" />
                    <SPLIT distance="150" swimtime="00:01:28.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103572" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="103608" number="2" />
                    <RELAYPOSITION athleteid="103589" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="103536" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="99059" points="257" reactiontime="+83" swimtime="00:02:26.91" resultid="104102" heatid="105240" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.10" />
                    <SPLIT distance="100" swimtime="00:01:20.50" />
                    <SPLIT distance="150" swimtime="00:01:57.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103553" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="103566" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="103589" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="103542" number="4" reactiontime="+63" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" points="270" reactiontime="+97" swimtime="00:02:11.13" resultid="104106" heatid="105309" lane="3" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                    <SPLIT distance="100" swimtime="00:01:08.05" />
                    <SPLIT distance="150" swimtime="00:01:39.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103553" number="1" reactiontime="+97" />
                    <RELAYPOSITION athleteid="103581" number="2" reactiontime="+74" />
                    <RELAYPOSITION athleteid="103542" number="3" reactiontime="+18" />
                    <RELAYPOSITION athleteid="103595" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="99036" points="361" reactiontime="+83" swimtime="00:02:28.91" resultid="104099" heatid="105238" lane="2" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                    <SPLIT distance="100" swimtime="00:01:20.73" />
                    <SPLIT distance="150" swimtime="00:01:54.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103517" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="103530" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="103558" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="103522" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="S 4/ 4 zmiana" eventid="99234" reactiontime="+100" status="DSQ" swimtime="00:00:00.00" resultid="104103" heatid="105307" lane="3" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                    <SPLIT distance="100" swimtime="00:01:06.89" />
                    <SPLIT distance="150" swimtime="00:01:40.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103517" number="1" reactiontime="+100" status="DSQ" />
                    <RELAYPOSITION athleteid="103522" number="2" reactiontime="+16" status="DSQ" />
                    <RELAYPOSITION athleteid="103530" number="3" reactiontime="+46" status="DSQ" />
                    <RELAYPOSITION athleteid="103558" number="4" reactiontime="-4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="307" reactiontime="+97" swimtime="00:02:05.73" resultid="104098" heatid="105160" lane="5" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.43" />
                    <SPLIT distance="100" swimtime="00:01:05.27" />
                    <SPLIT distance="150" swimtime="00:01:38.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103542" number="1" reactiontime="+97" />
                    <RELAYPOSITION athleteid="103558" number="2" reactiontime="+24" />
                    <RELAYPOSITION athleteid="103530" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="103509" number="4" reactiontime="+63" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" points="338" reactiontime="+78" swimtime="00:02:14.00" resultid="104107" heatid="105365" lane="7" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.20" />
                    <SPLIT distance="100" swimtime="00:01:13.86" />
                    <SPLIT distance="150" swimtime="00:01:47.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103517" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="103536" number="2" reactiontime="+38" />
                    <RELAYPOSITION athleteid="103558" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="103509" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="98846" points="245" reactiontime="+82" swimtime="00:02:15.56" resultid="104097" heatid="105160" lane="8" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                    <SPLIT distance="100" swimtime="00:01:12.92" />
                    <SPLIT distance="150" swimtime="00:01:46.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103517" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="103547" number="2" reactiontime="+82" />
                    <RELAYPOSITION athleteid="103492" number="3" />
                    <RELAYPOSITION athleteid="103501" number="4" reactiontime="+10" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="99441" points="155" reactiontime="+78" swimtime="00:02:53.78" resultid="104108" heatid="105364" lane="7" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.14" />
                    <SPLIT distance="100" swimtime="00:01:31.02" />
                    <SPLIT distance="150" swimtime="00:02:12.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103530" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="103599" number="2" reactiontime="+54" />
                    <RELAYPOSITION athleteid="103522" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="103547" number="4" reactiontime="+64" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="LOD" clubid="102060" name="AZS UŁ Pł Łódź">
          <CONTACT name="AZS UŁ PŁ ŁÓDŹ" state="LOD" street="Styrska 20" />
          <ATHLETES>
            <ATHLETE birthdate="1984-06-08" firstname="Marcin" gender="M" lastname="BABUCHOWSKI" nation="POL" swrid="4037687" athleteid="102061">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski Masters" eventid="98830" points="603" reactiontime="+77" swimtime="00:02:14.89" resultid="102062" heatid="105158" lane="4" entrytime="00:02:11.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.47" />
                    <SPLIT distance="100" swimtime="00:01:01.06" />
                    <SPLIT distance="150" swimtime="00:01:43.59" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="98924" points="603" reactiontime="+67" swimtime="00:00:28.44" resultid="102063" heatid="105190" lane="5" entrytime="00:00:27.60" entrycourse="LCM" />
                <RESULT comment="Rekord Polski Masters" eventid="98988" points="664" reactiontime="+76" swimtime="00:00:53.75" resultid="102064" heatid="105228" lane="4" entrytime="00:00:52.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="682" reactiontime="+77" swimtime="00:00:25.48" resultid="102065" heatid="105276" lane="4" entrytime="00:00:24.80" entrycourse="LCM" />
                <RESULT comment="Rekord Polski Masters" eventid="99218" points="589" reactiontime="+83" swimtime="00:02:01.62" resultid="102066" heatid="105305" lane="3" entrytime="00:02:05.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.52" />
                    <SPLIT distance="100" swimtime="00:01:00.66" />
                    <SPLIT distance="150" swimtime="00:01:31.85" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99361" points="683" reactiontime="+75" swimtime="00:00:56.56" resultid="102067" heatid="105331" lane="4" entrytime="00:00:55.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="102068" heatid="105343" lane="4" entrytime="00:02:14.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZSDG" nation="POL" region="SLA" clubid="102802" name="AZS WSB Dąbrowa Górnicza">
          <CONTACT email="kacperkapron@wp.pl" name="Kaproń Kacper" phone="791-512-012" state="ŚLĄSK" street="Mickiewicza 9/21a" zip="41-300" />
          <ATHLETES>
            <ATHLETE birthdate="1993-02-05" firstname="Kacper" gender="M" lastname="KAPROŃ" nation="POL" license="S02711200035" swrid="4086800" athleteid="102803">
              <RESULTS>
                <RESULT eventid="98924" points="356" reactiontime="+67" swimtime="00:00:33.90" resultid="102806" heatid="105187" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="102808" heatid="105275" lane="7" entrytime="00:00:28.00" />
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="102809" heatid="105303" lane="4" entrytime="00:02:14.00" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="102810" heatid="105362" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="102811" entrytime="00:04:50.00" />
                <RESULT eventid="98956" points="322" reactiontime="+76" swimtime="00:03:05.29" resultid="104383" heatid="105203" lane="5" entrytime="00:02:52.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.30" />
                    <SPLIT distance="100" swimtime="00:01:27.28" />
                    <SPLIT distance="150" swimtime="00:02:15.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="102938" name="AquaStars Gdynia">
          <ATHLETES>
            <ATHLETE birthdate="1978-01-01" firstname="Mariusz" gender="M" lastname="GOLON" nation="POL" athleteid="102939">
              <RESULTS>
                <RESULT eventid="98798" points="412" reactiontime="+83" swimtime="00:00:28.08" resultid="103047" heatid="105136" lane="6" entrytime="00:00:29.00" />
                <RESULT eventid="98830" points="324" reactiontime="+98" swimtime="00:02:45.89" resultid="103048" heatid="105153" lane="6" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                    <SPLIT distance="100" swimtime="00:01:15.27" />
                    <SPLIT distance="150" swimtime="00:02:05.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="355" reactiontime="+76" swimtime="00:00:33.93" resultid="103049" heatid="105188" lane="7" entrytime="00:00:33.00" />
                <RESULT eventid="98956" status="DNS" swimtime="00:00:00.00" resultid="103050" heatid="105201" lane="6" entrytime="00:03:10.00" />
                <RESULT eventid="99170" points="439" reactiontime="+87" swimtime="00:00:29.50" resultid="103051" heatid="105273" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="99186" points="329" reactiontime="+78" swimtime="00:01:15.17" resultid="103052" heatid="105285" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="293" reactiontime="+87" swimtime="00:02:48.45" resultid="103053" heatid="105340" lane="8" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.13" />
                    <SPLIT distance="100" swimtime="00:01:19.96" />
                    <SPLIT distance="150" swimtime="00:02:04.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="407" reactiontime="+83" swimtime="00:00:35.97" resultid="103054" heatid="105358" lane="6" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="102642" name="Aquapark Wrocław">
          <CONTACT name="Dudek" phone="665103411" />
          <ATHLETES>
            <ATHLETE birthdate="1988-07-21" firstname="Mateusz" gender="M" lastname="DUDEK" nation="POL" swrid="4072803" athleteid="103436">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="103437" heatid="105142" lane="7" entrytime="00:00:26.00" entrycourse="LCM" />
                <RESULT eventid="98956" points="492" reactiontime="+80" swimtime="00:02:40.85" resultid="103438" heatid="105204" lane="3" entrytime="00:02:34.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.49" />
                    <SPLIT distance="100" swimtime="00:01:16.06" />
                    <SPLIT distance="150" swimtime="00:01:57.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="570" reactiontime="+79" swimtime="00:01:10.50" resultid="103439" heatid="105258" lane="6" entrytime="00:01:09.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="103440" heatid="105362" lane="2" entrytime="00:00:31.66" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-07-05" firstname="Sebastian" gender="M" lastname="FIGARSKI" nation="POL" swrid="4754698" athleteid="103441">
              <RESULTS>
                <RESULT eventid="98924" points="490" reactiontime="+81" swimtime="00:00:30.49" resultid="103442" heatid="105190" lane="2" entrytime="00:00:29.50" entrycourse="LCM" />
                <RESULT eventid="99186" points="497" reactiontime="+75" swimtime="00:01:05.57" resultid="103443" heatid="105288" lane="6" entrytime="00:01:03.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="473" reactiontime="+77" swimtime="00:02:23.60" resultid="103444" heatid="105343" lane="3" entrytime="00:02:19.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                    <SPLIT distance="100" swimtime="00:01:08.58" />
                    <SPLIT distance="150" swimtime="00:01:46.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-04-06" firstname="Andrzej" gender="M" lastname="PERZ" nation="POL" athleteid="103445">
              <RESULTS>
                <RESULT eventid="98798" points="379" reactiontime="+94" swimtime="00:00:28.87" resultid="103446" heatid="105137" lane="5" entrytime="00:00:28.40" />
                <RESULT eventid="98988" points="346" reactiontime="+104" swimtime="00:01:06.78" resultid="103447" heatid="105222" lane="0" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="300" reactiontime="+89" swimtime="00:01:17.51" resultid="103448" heatid="105286" lane="0" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="274" reactiontime="+77" swimtime="00:02:52.13" resultid="103449" heatid="105341" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                    <SPLIT distance="100" swimtime="00:01:21.09" />
                    <SPLIT distance="150" swimtime="00:02:07.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-11-17" firstname="Michał" gender="M" lastname="STASIACZEK" nation="POL" swrid="4292725" athleteid="103450">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="103451" heatid="105141" lane="4" entrytime="00:00:26.50" />
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="103452" heatid="105157" lane="4" entrytime="00:02:29.00" />
                <RESULT eventid="99091" points="553" reactiontime="+83" swimtime="00:01:11.19" resultid="103453" heatid="105258" lane="2" entrytime="00:01:09.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="567" reactiontime="+73" swimtime="00:00:32.22" resultid="103454" heatid="105362" lane="7" entrytime="00:00:31.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-04-14" firstname="Mateusz" gender="M" lastname="KWAŚNIEWSKI" nation="POL" swrid="4382042" athleteid="103455">
              <RESULTS>
                <RESULT eventid="99170" points="516" reactiontime="+69" swimtime="00:00:27.95" resultid="103457" heatid="105276" lane="7" entrytime="00:00:26.90" />
                <RESULT eventid="99218" points="462" reactiontime="+73" swimtime="00:02:11.86" resultid="103458" heatid="105305" lane="4" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.31" />
                    <SPLIT distance="100" swimtime="00:01:02.21" />
                    <SPLIT distance="150" swimtime="00:01:36.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="439" reactiontime="+90" swimtime="00:04:49.54" resultid="103459" heatid="106059" lane="3" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                    <SPLIT distance="100" swimtime="00:01:08.43" />
                    <SPLIT distance="150" swimtime="00:01:45.91" />
                    <SPLIT distance="200" swimtime="00:02:23.23" />
                    <SPLIT distance="250" swimtime="00:03:00.42" />
                    <SPLIT distance="300" swimtime="00:03:37.59" />
                    <SPLIT distance="350" swimtime="00:04:14.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="569" reactiontime="+62" swimtime="00:00:56.61" resultid="104370" heatid="105228" lane="7" entrytime="00:00:54.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-05-11" firstname="Joanna" gender="F" lastname="KROWICKA" nation="POL" athleteid="103460">
              <RESULTS>
                <RESULT eventid="98777" points="227" reactiontime="+101" swimtime="00:00:38.88" resultid="103461" heatid="105116" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="98814" points="159" reactiontime="+113" swimtime="00:03:52.71" resultid="103462" heatid="105145" lane="1" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.11" />
                    <SPLIT distance="100" swimtime="00:01:52.17" />
                    <SPLIT distance="150" swimtime="00:02:57.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="213" reactiontime="+95" swimtime="00:03:52.72" resultid="103463" heatid="105193" lane="2" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.73" />
                    <SPLIT distance="100" swimtime="00:01:51.77" />
                    <SPLIT distance="150" swimtime="00:02:54.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="166" reactiontime="+110" swimtime="00:01:34.62" resultid="103464" heatid="105208" lane="1" entrytime="00:01:19.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="232" reactiontime="+100" swimtime="00:01:44.58" resultid="103465" heatid="105245" lane="7" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="136" reactiontime="+93" swimtime="00:00:48.65" resultid="103466" heatid="105261" lane="8" entrytime="00:00:39.99" />
                <RESULT eventid="99409" points="256" reactiontime="+102" swimtime="00:00:46.38" resultid="103467" heatid="105348" lane="9" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-11-20" firstname="Katarzyna" gender="F" lastname="STASZKIEWICZ" nation="POL" swrid="4071838" athleteid="103468">
              <RESULTS>
                <RESULT eventid="98777" status="DNS" swimtime="00:00:00.00" resultid="103469" heatid="105121" lane="7" entrytime="00:00:28.85" entrycourse="LCM" />
                <RESULT eventid="98907" points="564" reactiontime="+73" swimtime="00:00:32.74" resultid="103470" heatid="105177" lane="8" entrytime="00:00:38.00" />
                <RESULT eventid="98972" points="710" reactiontime="+81" swimtime="00:00:58.34" resultid="103471" heatid="105212" lane="5" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="633" reactiontime="+81" swimtime="00:00:29.19" resultid="103472" heatid="105263" lane="3" entrytime="00:00:34.00" />
                <RESULT eventid="99409" points="540" reactiontime="+84" swimtime="00:00:36.19" resultid="103473" heatid="105349" lane="0" entrytime="00:00:39.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-12-04" firstname="Karolina" gender="F" lastname="WCISŁO" nation="POL" athleteid="103474">
              <RESULTS>
                <RESULT eventid="98777" status="DNS" swimtime="00:00:00.00" resultid="103475" heatid="105117" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="98907" points="229" reactiontime="+76" swimtime="00:00:44.17" resultid="103476" heatid="105177" lane="7" entrytime="00:00:38.00" />
                <RESULT eventid="98972" status="DNS" swimtime="00:00:00.00" resultid="103477" heatid="105210" lane="5" entrytime="00:01:12.00" />
                <RESULT eventid="99154" status="DNS" swimtime="00:00:00.00" resultid="103478" heatid="105262" lane="0" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99250" points="501" reactiontime="+80" swimtime="00:01:46.80" resultid="103479" heatid="105308" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.52" />
                    <SPLIT distance="100" swimtime="00:00:53.00" />
                    <SPLIT distance="150" swimtime="00:01:18.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103450" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="103436" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="103455" number="3" reactiontime="+30" />
                    <RELAYPOSITION athleteid="103445" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="99059" points="529" reactiontime="+69" swimtime="00:01:55.52" resultid="103480" heatid="105240" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.96" />
                    <SPLIT distance="100" swimtime="00:01:02.14" />
                    <SPLIT distance="150" swimtime="00:01:29.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103441" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="103436" number="2" />
                    <RELAYPOSITION athleteid="103455" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="103450" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="104375" name="Białystok">
          <ATHLETES>
            <ATHLETE birthdate="1963-01-16" firstname="Wojciech" gender="M" lastname="ŻMIEJKO" nation="POL" swrid="4186249" athleteid="100126">
              <RESULTS>
                <RESULT eventid="98798" points="399" reactiontime="+87" swimtime="00:00:28.38" resultid="100127" heatid="105137" lane="2" entrytime="00:00:28.50" />
                <RESULT eventid="98830" points="366" reactiontime="+80" swimtime="00:02:39.24" resultid="100128" heatid="105155" lane="8" entrytime="00:02:41.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.97" />
                    <SPLIT distance="100" swimtime="00:01:15.33" />
                    <SPLIT distance="150" swimtime="00:02:02.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="418" reactiontime="+86" swimtime="00:01:02.70" resultid="100129" heatid="105223" lane="4" entrytime="00:01:02.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="408" reactiontime="+84" swimtime="00:00:30.22" resultid="100130" heatid="105272" lane="4" entrytime="00:00:30.85" />
                <RESULT eventid="99186" points="314" reactiontime="+85" swimtime="00:01:16.39" resultid="100131" heatid="105285" lane="5" entrytime="00:01:15.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="354" reactiontime="+90" swimtime="00:01:10.39" resultid="100132" heatid="105329" lane="5" entrytime="00:01:10.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="268" reactiontime="+72" swimtime="00:02:53.40" resultid="100133" heatid="105341" lane="9" entrytime="00:02:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.24" />
                    <SPLIT distance="100" swimtime="00:01:24.15" />
                    <SPLIT distance="150" swimtime="00:02:09.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CM UJ MAST" nation="POL" region="MAL" clubid="100475" name="Collegium Medicum UJ Mrs Kraków" shortname="Collegium Medicum UJ Masters K">
          <CONTACT city="Kraków" email="MariuszBaranik@gmail.com" name="Mariusz Baranik" street="Białoprądnicka 32c/3" zip="31-221" />
          <ATHLETES>
            <ATHLETE birthdate="1969-06-29" firstname="Mariusz" gender="M" lastname="BARANIK" nation="POL" swrid="4992740" athleteid="100476">
              <RESULTS>
                <RESULT eventid="98798" points="450" reactiontime="+85" swimtime="00:00:27.27" resultid="100477" heatid="105140" lane="5" entrytime="00:00:27.00" />
                <RESULT eventid="98988" points="435" reactiontime="+79" swimtime="00:01:01.89" resultid="100478" heatid="105224" lane="6" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="462" reactiontime="+76" swimtime="00:00:29.01" resultid="100479" heatid="105273" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="100480" heatid="105329" lane="3" entrytime="00:01:11.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="CYP" clubid="102838" name="Cyprus Masters Swimming Federation" shortname="Cyprus Mrs Swiim. Fed.">
          <CONTACT email="p.koush@cytanet.com.cy" name="Pavlos Koushappas" />
          <ATHLETES>
            <ATHLETE birthdate="1965-12-27" firstname="Costas" gender="M" lastname="CHRISTOFOROU" nation="CYP" swrid="4877693" athleteid="102839">
              <RESULTS>
                <RESULT eventid="98830" points="331" reactiontime="+89" swimtime="00:02:44.75" resultid="102840" heatid="105156" lane="0" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                    <SPLIT distance="100" swimtime="00:01:17.22" />
                    <SPLIT distance="150" swimtime="00:02:08.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" reactiontime="+83" status="DNF" swimtime="00:00:00.00" resultid="102841" heatid="105234" lane="4" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                    <SPLIT distance="100" swimtime="00:01:23.41" />
                    <SPLIT distance="150" swimtime="00:02:17.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="354" reactiontime="+85" swimtime="00:02:24.08" resultid="102842" heatid="105301" lane="5" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.14" />
                    <SPLIT distance="100" swimtime="00:01:09.71" />
                    <SPLIT distance="150" swimtime="00:01:47.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="246" reactiontime="+84" swimtime="00:01:19.45" resultid="102843" heatid="105329" lane="1" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-08-11" firstname="Costas" gender="M" lastname="KOUSHAPPAS" nation="CYP" swrid="4967112" athleteid="102844">
              <RESULTS>
                <RESULT eventid="98891" points="199" swimtime="00:24:51.31" resultid="102845" heatid="105423" lane="7" entrytime="00:23:59.00" />
                <RESULT eventid="98956" points="216" reactiontime="+108" swimtime="00:03:31.55" resultid="102846" heatid="105198" lane="8" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.18" />
                    <SPLIT distance="100" swimtime="00:01:41.08" />
                    <SPLIT distance="150" swimtime="00:02:37.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="102847" heatid="105250" lane="9" entrytime="00:01:53.00" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="102848" heatid="105355" lane="1" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-08-11" firstname="Pavlos" gender="M" lastname="KOUSHAPPAS" nation="CYP" swrid="4877694" athleteid="102849">
              <RESULTS>
                <RESULT eventid="98798" points="339" reactiontime="+92" swimtime="00:00:29.96" resultid="102850" heatid="105135" lane="4" entrytime="00:00:29.10" />
                <RESULT eventid="99282" points="170" reactiontime="+115" swimtime="00:07:19.49" resultid="102851" heatid="106050" lane="3" entrytime="00:06:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.54" />
                    <SPLIT distance="100" swimtime="00:01:49.67" />
                    <SPLIT distance="150" swimtime="00:02:47.59" />
                    <SPLIT distance="200" swimtime="00:03:42.81" />
                    <SPLIT distance="250" swimtime="00:04:48.23" />
                    <SPLIT distance="300" swimtime="00:05:51.37" />
                    <SPLIT distance="350" swimtime="00:06:36.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="172" reactiontime="+104" swimtime="00:03:21.18" resultid="102852" heatid="105338" lane="0" entrytime="00:03:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.78" />
                    <SPLIT distance="100" swimtime="00:01:42.40" />
                    <SPLIT distance="150" swimtime="00:02:35.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="230" reactiontime="+94" swimtime="00:05:58.76" resultid="102853" heatid="106064" lane="4" entrytime="00:05:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.13" />
                    <SPLIT distance="100" swimtime="00:01:22.34" />
                    <SPLIT distance="150" swimtime="00:02:08.50" />
                    <SPLIT distance="200" swimtime="00:02:55.31" />
                    <SPLIT distance="250" swimtime="00:03:42.53" />
                    <SPLIT distance="300" swimtime="00:04:28.75" />
                    <SPLIT distance="350" swimtime="00:05:14.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-01-28" firstname="Larrys" gender="M" lastname="FYLACTOU" nation="CYP" athleteid="102854">
              <RESULTS>
                <RESULT eventid="98798" points="432" reactiontime="+91" swimtime="00:00:27.65" resultid="102855" heatid="105141" lane="6" entrytime="00:00:26.50" />
                <RESULT eventid="98924" points="339" reactiontime="+100" swimtime="00:00:34.45" resultid="102856" heatid="105188" lane="1" entrytime="00:00:33.00" />
                <RESULT eventid="98988" points="423" reactiontime="+80" swimtime="00:01:02.46" resultid="102857" heatid="105225" lane="5" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="335" reactiontime="+80" swimtime="00:00:32.28" resultid="102858" heatid="105272" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="99186" points="258" reactiontime="+91" swimtime="00:01:21.56" resultid="102859" heatid="105286" lane="2" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="348" reactiontime="+79" swimtime="00:00:37.90" resultid="102860" heatid="105357" lane="1" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-01-15" firstname="Costas" gender="M" lastname="HAILIS" nation="CYP" athleteid="102861">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="102862" heatid="105142" lane="3" entrytime="00:00:25.60" />
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="102863" heatid="105158" lane="1" entrytime="00:02:22.00" />
                <RESULT eventid="98924" status="DNS" swimtime="00:00:00.00" resultid="102864" heatid="105190" lane="9" entrytime="00:00:30.01" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="102865" heatid="105228" lane="0" entrytime="00:00:56.90" />
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="102866" heatid="105275" lane="4" entrytime="00:00:27.50" />
                <RESULT eventid="99186" status="DNS" swimtime="00:00:00.00" resultid="102867" heatid="105288" lane="1" entrytime="00:01:05.00" />
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="102868" heatid="105343" lane="7" entrytime="00:02:25.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Cyprus Masters Swimmin Federation" number="1">
              <RESULTS>
                <RESULT eventid="99059" points="296" reactiontime="+72" swimtime="00:02:20.10" resultid="102869" heatid="105240" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.92" />
                    <SPLIT distance="100" swimtime="00:01:19.03" />
                    <SPLIT distance="150" swimtime="00:01:49.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102854" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="102839" number="2" reactiontime="+84" />
                    <RELAYPOSITION athleteid="102844" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="102849" number="4" reactiontime="+70" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" points="371" reactiontime="+75" swimtime="00:01:58.01" resultid="102870" heatid="105308" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.57" />
                    <SPLIT distance="100" swimtime="00:00:56.85" />
                    <SPLIT distance="150" swimtime="00:01:30.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102839" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="102854" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="102849" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="102844" number="4" reactiontime="+70" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="LOD" clubid="101079" name="Delfin Masters Łódz">
          <CONTACT city="ŁÓDZ" email="roman.wiczel@gmail.com" name="WICZEL" phone="691-928-922" state="ŁÓDZK" street="FLORECISTÓW 3 B" zip="94-042" />
          <ATHLETES>
            <ATHLETE birthdate="1969-06-03" firstname="Tomasz" gender="M" lastname="WIADERNY" nation="POL" athleteid="101080">
              <RESULTS>
                <RESULT eventid="98988" points="205" reactiontime="+95" swimtime="00:01:19.52" resultid="101081" heatid="105216" lane="4" entrytime="00:01:15.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="186" reactiontime="+92" swimtime="00:00:39.23" resultid="101082" heatid="105266" lane="6" entrytime="00:00:42.50" entrycourse="LCM" />
                <RESULT eventid="99218" points="155" reactiontime="+103" swimtime="00:03:09.80" resultid="101083" heatid="105301" lane="1" entrytime="00:02:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.23" />
                    <SPLIT distance="100" swimtime="00:01:27.54" />
                    <SPLIT distance="150" swimtime="00:02:20.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-05-26" firstname="Ewa" gender="F" lastname="CIEPLUCHA" nation="POL" athleteid="101084">
              <RESULTS>
                <RESULT eventid="98907" points="357" reactiontime="+71" swimtime="00:00:38.12" resultid="101085" heatid="105177" lane="5" entrytime="00:00:36.20" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-03-16" firstname="Janusz" gender="M" lastname="BŁASIAK" nation="POL" athleteid="101086">
              <RESULTS>
                <RESULT eventid="98830" points="76" reactiontime="+113" swimtime="00:04:28.60" resultid="101087" heatid="105148" lane="4" entrytime="00:04:36.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.06" />
                    <SPLIT distance="100" swimtime="00:02:13.82" />
                    <SPLIT distance="150" swimtime="00:03:32.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="69" reactiontime="+107" swimtime="00:00:58.53" resultid="101088" heatid="105180" lane="4" entrytime="00:00:58.30" entrycourse="LCM" />
                <RESULT eventid="99020" points="49" reactiontime="+111" swimtime="00:05:04.30" resultid="101089" heatid="105234" lane="0" entrytime="00:03:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.97" />
                    <SPLIT distance="100" swimtime="00:02:23.29" />
                    <SPLIT distance="150" swimtime="00:03:45.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="67" reactiontime="+114" swimtime="00:00:55.00" resultid="101090" heatid="105265" lane="3" entrytime="00:00:56.74" entrycourse="LCM" />
                <RESULT eventid="99361" points="49" reactiontime="+111" swimtime="00:02:16.13" resultid="101091" heatid="105325" lane="1" entrytime="00:02:07.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="106116" heatid="105350" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-05-15" firstname="Grzegorz" gender="M" lastname="KĘDZIORA" nation="POL" athleteid="101092">
              <RESULTS>
                <RESULT eventid="99020" reactiontime="+108" status="DNF" swimtime="00:00:00.00" resultid="101093" heatid="105236" lane="5" entrytime="00:02:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                    <SPLIT distance="100" swimtime="00:01:13.96" />
                    <SPLIT distance="150" swimtime="00:02:33.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="444" reactiontime="+78" swimtime="00:00:29.39" resultid="101094" heatid="105274" lane="5" entrytime="00:00:28.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-04-11" firstname="Rafał" gender="M" lastname="MACIEJEWSKI" nation="POL" athleteid="101095">
              <RESULTS>
                <RESULT eventid="98988" points="234" reactiontime="+95" swimtime="00:01:16.09" resultid="101096" heatid="105221" lane="0" entrytime="00:01:07.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="162" reactiontime="+72" swimtime="00:01:35.09" resultid="101097" heatid="105286" lane="8" entrytime="00:01:14.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-14" firstname="Wojciech" gender="M" lastname="URBAŃSKI" nation="POL" athleteid="101098">
              <RESULTS>
                <RESULT eventid="98988" points="373" reactiontime="+101" swimtime="00:01:05.14" resultid="101099" heatid="105222" lane="7" entrytime="00:01:04.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="399" reactiontime="+103" swimtime="00:00:30.45" resultid="101100" heatid="105272" lane="0" entrytime="00:00:31.20" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-03-05" firstname="Adam" gender="M" lastname="JERZYKOWSKI" nation="POL" athleteid="101101">
              <RESULTS>
                <RESULT eventid="98798" points="272" reactiontime="+88" swimtime="00:00:32.25" resultid="101102" heatid="105124" lane="3" entrytime="00:00:41.80" entrycourse="LCM" />
                <RESULT eventid="98988" points="272" reactiontime="+68" swimtime="00:01:12.40" resultid="101103" heatid="105215" lane="9" entrytime="00:01:25.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="101104" heatid="106064" lane="0" entrytime="00:06:15.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-04-10" firstname="Grzegorz" gender="M" lastname="ROGALSKI" nation="POL" athleteid="101105">
              <RESULTS>
                <RESULT eventid="98988" points="419" reactiontime="+95" swimtime="00:01:02.66" resultid="101106" heatid="105223" lane="0" entrytime="00:01:03.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="383" reactiontime="+94" swimtime="00:00:30.88" resultid="101107" heatid="105273" lane="2" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="101108" heatid="105303" lane="7" entrytime="00:02:15.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-24" firstname="Piotr" gender="M" lastname="GEADE" nation="POL" athleteid="101109">
              <RESULTS>
                <RESULT eventid="99091" points="319" reactiontime="+74" swimtime="00:01:25.51" resultid="101110" heatid="105255" lane="8" entrytime="00:01:22.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99059" points="308" reactiontime="+77" swimtime="00:02:18.26" resultid="101111" heatid="105241" lane="4" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                    <SPLIT distance="100" swimtime="00:01:19.61" />
                    <SPLIT distance="150" swimtime="00:01:50.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101095" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="101109" number="2" reactiontime="+33" />
                    <RELAYPOSITION athleteid="101105" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="101092" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" points="391" reactiontime="+101" swimtime="00:01:56.00" resultid="101112" heatid="105311" lane="0" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.20" />
                    <SPLIT distance="100" swimtime="00:01:01.08" />
                    <SPLIT distance="150" swimtime="00:01:28.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101095" number="1" reactiontime="+101" />
                    <RELAYPOSITION athleteid="101098" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="101105" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="101092" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="99059" points="171" reactiontime="+73" swimtime="00:02:48.08" resultid="101113" heatid="105241" lane="6" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.20" />
                    <SPLIT distance="100" swimtime="00:01:45.69" />
                    <SPLIT distance="150" swimtime="00:01:54.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101086" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="101080" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="101098" number="3" reactiontime="+74" />
                    <RELAYPOSITION athleteid="101101" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" points="229" reactiontime="+109" swimtime="00:02:18.66" resultid="101114" heatid="105310" lane="7" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.12" />
                    <SPLIT distance="100" swimtime="00:01:14.42" />
                    <SPLIT distance="150" swimtime="00:01:46.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101086" number="1" reactiontime="+109" />
                    <RELAYPOSITION athleteid="101080" number="2" reactiontime="+85" />
                    <RELAYPOSITION athleteid="101109" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="101101" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="DEOSIE" nation="POL" region="KUJ" clubid="104952" name="Dęby Osielsko">
          <CONTACT city="Osielsko" email="wfadrian@gmail.com" name="Chwaliszewski" phone="694273582" state="KUJ-P" street="Centralna 7" zip="86-031" />
          <ATHLETES>
            <ATHLETE birthdate="1976-11-02" firstname="Tomasz" gender="M" lastname="CHWALISZEWSKI" nation="POL" athleteid="102800">
              <RESULTS>
                <RESULT eventid="98891" points="131" swimtime="00:28:32.85" resultid="102801" heatid="105422" lane="3" entrytime="00:22:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-09-12" firstname="Adrian" gender="M" lastname="TEODORSKI" nation="POL" swrid="4071733" athleteid="104953">
              <RESULTS>
                <RESULT eventid="98830" points="396" reactiontime="+93" swimtime="00:02:35.22" resultid="104954" heatid="105157" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.23" />
                    <SPLIT distance="100" swimtime="00:01:10.28" />
                    <SPLIT distance="150" swimtime="00:01:59.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="332" swimtime="00:20:57.62" resultid="104955" heatid="105421" lane="1" entrytime="00:21:12.00" />
                <RESULT eventid="98956" points="281" reactiontime="+97" swimtime="00:03:13.69" resultid="104956" heatid="105202" lane="5" entrytime="00:03:00.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.62" />
                    <SPLIT distance="100" swimtime="00:01:32.75" />
                    <SPLIT distance="150" swimtime="00:02:23.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="345" reactiontime="+111" swimtime="00:02:38.85" resultid="104957" heatid="105236" lane="0" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.28" />
                    <SPLIT distance="100" swimtime="00:01:13.95" />
                    <SPLIT distance="150" swimtime="00:01:55.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="310" reactiontime="+85" swimtime="00:01:26.32" resultid="104958" heatid="105257" lane="8" entrytime="00:01:17.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="364" reactiontime="+106" swimtime="00:05:41.24" resultid="104959" heatid="106051" lane="2" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.28" />
                    <SPLIT distance="100" swimtime="00:01:08.41" />
                    <SPLIT distance="150" swimtime="00:01:56.77" />
                    <SPLIT distance="200" swimtime="00:02:43.29" />
                    <SPLIT distance="250" swimtime="00:03:34.54" />
                    <SPLIT distance="300" swimtime="00:04:26.31" />
                    <SPLIT distance="350" swimtime="00:05:04.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="478" reactiontime="+86" swimtime="00:01:03.70" resultid="104960" heatid="105331" lane="8" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="341" reactiontime="+94" swimtime="00:02:40.14" resultid="104961" heatid="105343" lane="9" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.55" />
                    <SPLIT distance="100" swimtime="00:01:18.74" />
                    <SPLIT distance="150" swimtime="00:02:00.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="102688" name="Gdynia Masters">
          <CONTACT email="k.mysiak@wpit.am.gdynia.pl" name="Mysiak Katarzyna" />
          <ATHLETES>
            <ATHLETE birthdate="1959-01-01" firstname="Renata" gender="F" lastname="POLAŃCZYK" nation="POL" swrid="4754664" athleteid="102696">
              <RESULTS>
                <RESULT eventid="98814" status="DNS" swimtime="00:00:00.00" resultid="102697" heatid="105144" lane="3" entrytime="00:03:46.65" />
                <RESULT eventid="98863" points="209" swimtime="00:13:52.03" resultid="102698" heatid="105405" lane="9" entrytime="00:13:49.65" />
                <RESULT eventid="99004" status="DNS" swimtime="00:00:00.00" resultid="102700" heatid="105229" lane="5" entrytime="00:04:10.53" />
                <RESULT eventid="99266" points="166" reactiontime="+127" swimtime="00:08:07.65" resultid="102702" heatid="106046" lane="0" entrytime="00:07:59.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.89" />
                    <SPLIT distance="100" swimtime="00:01:59.04" />
                    <SPLIT distance="150" swimtime="00:02:57.87" />
                    <SPLIT distance="200" swimtime="00:03:53.85" />
                    <SPLIT distance="250" swimtime="00:05:10.82" />
                    <SPLIT distance="300" swimtime="00:06:28.03" />
                    <SPLIT distance="350" swimtime="00:07:21.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="177" reactiontime="+82" swimtime="00:03:40.92" resultid="102703" heatid="105332" lane="4" entrytime="00:03:30.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.47" />
                    <SPLIT distance="100" swimtime="00:01:48.99" />
                    <SPLIT distance="150" swimtime="00:02:47.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" status="DNS" swimtime="00:00:00.00" resultid="102704" heatid="106056" lane="7" entrytime="00:06:48.96" />
                <RESULT eventid="99202" status="DNS" swimtime="00:00:00.00" resultid="105102" heatid="105290" lane="0" entrytime="00:03:30.00" />
                <RESULT eventid="99344" points="99" reactiontime="+109" swimtime="00:02:00.74" resultid="105103" heatid="105321" lane="7" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1934-01-01" firstname="Bogdan" gender="M" lastname="CIUNDZIEWCKI" nation="POL" athleteid="102705">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski Masters" eventid="98924" points="126" reactiontime="+74" swimtime="00:00:47.91" resultid="102706" heatid="105182" lane="6" entrytime="00:00:48.00" />
                <RESULT eventid="98956" status="DNS" swimtime="00:00:00.00" resultid="102707" heatid="105197" lane="2" entrytime="00:03:55.00" />
                <RESULT comment="Rekord Polski Masters" eventid="99091" points="154" swimtime="00:01:48.92" resultid="102708" heatid="105250" lane="0" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="161" swimtime="00:00:48.98" resultid="102709" heatid="105352" lane="6" entrytime="00:00:47.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-01-01" firstname="Hanka" gender="F" lastname="KANIA" nation="POL" swrid="4754667" athleteid="102710">
              <RESULTS>
                <RESULT eventid="98814" points="166" reactiontime="+114" swimtime="00:03:49.08" resultid="102711" heatid="105144" lane="6" entrytime="00:03:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.74" />
                    <SPLIT distance="100" swimtime="00:01:56.41" />
                    <SPLIT distance="150" swimtime="00:02:57.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="200" reactiontime="+103" swimtime="00:03:57.76" resultid="102712" heatid="105192" lane="8" entrytime="00:04:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.65" />
                    <SPLIT distance="100" swimtime="00:01:53.86" />
                    <SPLIT distance="150" swimtime="00:02:56.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="196" reactiontime="+86" swimtime="00:01:29.49" resultid="102713" heatid="105206" lane="3" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="186" reactiontime="+121" swimtime="00:01:52.67" resultid="102714" heatid="105244" lane="4" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="160" reactiontime="+123" swimtime="00:03:27.78" resultid="102715" heatid="105290" lane="2" entrytime="00:03:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.38" />
                    <SPLIT distance="100" swimtime="00:01:39.36" />
                    <SPLIT distance="150" swimtime="00:02:34.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="103" reactiontime="+118" swimtime="00:01:59.18" resultid="102716" heatid="105321" lane="3" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="196" reactiontime="+112" swimtime="00:00:50.69" resultid="102717" heatid="105345" lane="2" entrytime="00:00:52.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Katarzyna" gender="F" lastname="MAZUREK" nation="POL" swrid="4191116" athleteid="102718">
              <RESULTS>
                <RESULT eventid="98777" points="271" reactiontime="+95" swimtime="00:00:36.66" resultid="102719" heatid="105116" lane="2" entrytime="00:00:36.37" entrycourse="SCM" />
                <RESULT eventid="98972" points="222" reactiontime="+108" swimtime="00:01:25.91" resultid="102720" heatid="105207" lane="6" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99004" status="DNS" swimtime="00:00:00.00" resultid="102721" heatid="105229" lane="4" entrytime="00:04:10.00" />
                <RESULT eventid="99089" points="233" reactiontime="+99" swimtime="00:01:44.48" resultid="102722" heatid="105246" lane="6" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="190" reactiontime="+99" swimtime="00:00:43.55" resultid="102723" heatid="105260" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="99344" points="157" reactiontime="+107" swimtime="00:01:43.63" resultid="102724" heatid="105322" lane="2" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="283" reactiontime="+93" swimtime="00:00:44.90" resultid="102725" heatid="105348" lane="6" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-01-01" firstname="Katarzyna" gender="F" lastname="MYSIAK" nation="POL" swrid="4754669" athleteid="102726">
              <RESULTS>
                <RESULT eventid="98777" points="223" reactiontime="+110" swimtime="00:00:39.10" resultid="102727" heatid="105115" lane="4" entrytime="00:00:37.64" entrycourse="SCM" />
                <RESULT eventid="98907" points="205" reactiontime="+79" swimtime="00:00:45.83" resultid="102728" heatid="105174" lane="5" entrytime="00:00:44.00" />
                <RESULT eventid="98972" points="192" reactiontime="+101" swimtime="00:01:30.21" resultid="102729" heatid="105207" lane="9" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" status="DNS" swimtime="00:00:00.00" resultid="102730" heatid="105260" lane="0" entrytime="00:00:44.00" />
                <RESULT eventid="99202" points="174" swimtime="00:03:22.05" resultid="102731" heatid="105290" lane="8" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.90" />
                    <SPLIT distance="100" swimtime="00:01:37.06" />
                    <SPLIT distance="150" swimtime="00:02:30.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="180" swimtime="00:07:02.78" resultid="102732" heatid="106056" lane="8" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.59" />
                    <SPLIT distance="100" swimtime="00:01:34.99" />
                    <SPLIT distance="150" swimtime="00:02:29.70" />
                    <SPLIT distance="200" swimtime="00:03:24.07" />
                    <SPLIT distance="250" swimtime="00:04:19.80" />
                    <SPLIT distance="300" swimtime="00:05:15.22" />
                    <SPLIT distance="350" swimtime="00:06:11.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Czesław" gender="M" lastname="MIKOŁAJCZYK" nation="POL" swrid="4754640" athleteid="102733">
              <RESULTS>
                <RESULT eventid="98830" points="146" reactiontime="+99" swimtime="00:03:36.13" resultid="102734" heatid="105150" lane="4" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.75" />
                    <SPLIT distance="100" swimtime="00:01:49.60" />
                    <SPLIT distance="150" swimtime="00:02:46.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" status="DNS" swimtime="00:00:00.00" resultid="102735" heatid="105199" lane="0" entrytime="00:03:40.00" />
                <RESULT eventid="99091" points="174" reactiontime="+99" swimtime="00:01:44.57" resultid="102736" heatid="105251" lane="6" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="141" reactiontime="+107" swimtime="00:07:47.46" resultid="102737" heatid="106049" lane="2" entrytime="00:07:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.88" />
                    <SPLIT distance="100" swimtime="00:01:56.35" />
                    <SPLIT distance="150" swimtime="00:03:00.58" />
                    <SPLIT distance="200" swimtime="00:04:03.10" />
                    <SPLIT distance="250" swimtime="00:05:01.89" />
                    <SPLIT distance="300" swimtime="00:06:01.55" />
                    <SPLIT distance="350" swimtime="00:06:55.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="202" reactiontime="+99" swimtime="00:00:45.39" resultid="102738" heatid="105353" lane="2" entrytime="00:00:45.00" />
                <RESULT eventid="99020" points="98" reactiontime="+102" swimtime="00:04:01.63" resultid="105096" heatid="105233" lane="7" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.80" />
                    <SPLIT distance="100" swimtime="00:01:53.34" />
                    <SPLIT distance="150" swimtime="00:02:57.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-01-01" firstname="Anna" gender="F" lastname="WALCZAK" nation="POL" swrid="4754666" athleteid="102739">
              <RESULTS>
                <RESULT eventid="98777" points="122" reactiontime="+108" swimtime="00:00:47.77" resultid="102740" heatid="105113" lane="6" entrytime="00:00:46.66" entrycourse="SCM" />
                <RESULT eventid="98907" points="149" reactiontime="+70" swimtime="00:00:50.96" resultid="102741" heatid="105173" lane="7" entrytime="00:00:52.00" />
                <RESULT eventid="98972" status="DNS" swimtime="00:00:00.00" resultid="102742" heatid="105206" lane="8" entrytime="00:01:52.00" />
                <RESULT eventid="99314" points="120" reactiontime="+71" swimtime="00:01:57.53" resultid="102743" heatid="105277" lane="5" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-01-01" firstname="Andrzej" gender="M" lastname="SKWARŁO" nation="POL" swrid="4302086" athleteid="102744">
              <RESULTS>
                <RESULT eventid="98830" points="102" reactiontime="+106" swimtime="00:04:03.84" resultid="102745" heatid="105150" lane="9" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.29" />
                    <SPLIT distance="100" swimtime="00:01:59.53" />
                    <SPLIT distance="150" swimtime="00:03:07.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="113" reactiontime="+96" swimtime="00:00:49.61" resultid="102746" heatid="105182" lane="5" entrytime="00:00:47.50" />
                <RESULT eventid="98956" status="DNS" swimtime="00:00:00.00" resultid="102747" heatid="105197" lane="1" entrytime="00:03:56.00" />
                <RESULT eventid="99091" points="150" reactiontime="+114" swimtime="00:01:49.87" resultid="102748" heatid="105250" lane="5" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="96" reactiontime="+106" swimtime="00:01:53.28" resultid="102749" heatid="105282" lane="1" entrytime="00:01:50.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="92" reactiontime="+94" swimtime="00:04:07.38" resultid="102750" heatid="105337" lane="8" entrytime="00:04:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.63" />
                    <SPLIT distance="100" swimtime="00:01:56.29" />
                    <SPLIT distance="150" swimtime="00:03:01.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="174" reactiontime="+107" swimtime="00:00:47.74" resultid="102751" heatid="105354" lane="8" entrytime="00:00:43.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-24" firstname="Andrzej" gender="M" lastname="JACASZEK" nation="POL" swrid="4992743" athleteid="102752">
              <RESULTS>
                <RESULT eventid="98798" points="196" reactiontime="+87" swimtime="00:00:35.94" resultid="103034" heatid="105127" lane="9" entrytime="00:00:36.00" />
                <RESULT eventid="98956" points="183" swimtime="00:03:43.40" resultid="103035" heatid="105199" lane="7" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.24" />
                    <SPLIT distance="100" swimtime="00:01:44.62" />
                    <SPLIT distance="150" swimtime="00:02:45.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="231" reactiontime="+104" swimtime="00:01:35.19" resultid="103036" heatid="105251" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="262" reactiontime="+92" swimtime="00:00:41.65" resultid="104374" heatid="105355" lane="7" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-01" firstname="Danuta" gender="F" lastname="RADKOWIAK" nation="POL" swrid="4992757" athleteid="102753">
              <RESULTS>
                <RESULT eventid="98777" reactiontime="+94" status="DNS" swimtime="00:00:00.00" resultid="102754" heatid="105116" lane="3" entrytime="00:00:36.00" />
                <RESULT eventid="98814" status="DNS" swimtime="00:00:00.00" resultid="102755" heatid="105144" lane="2" entrytime="00:04:00.00" />
                <RESULT eventid="98940" status="DNS" swimtime="00:00:00.00" resultid="102756" heatid="105192" lane="7" entrytime="00:04:00.00" />
                <RESULT eventid="99004" status="DNS" swimtime="00:00:00.00" resultid="102757" heatid="105230" lane="0" entrytime="00:04:00.00" />
                <RESULT eventid="99154" status="DNS" swimtime="00:00:00.00" resultid="102758" heatid="105259" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="99266" points="117" reactiontime="+115" swimtime="00:09:07.41" resultid="102759" heatid="106045" lane="4" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.52" />
                    <SPLIT distance="100" swimtime="00:02:04.88" />
                    <SPLIT distance="150" swimtime="00:03:25.52" />
                    <SPLIT distance="200" swimtime="00:04:45.20" />
                    <SPLIT distance="250" swimtime="00:05:53.82" />
                    <SPLIT distance="300" swimtime="00:07:03.79" />
                    <SPLIT distance="350" swimtime="00:08:05.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" status="DNS" swimtime="00:00:00.00" resultid="102760" heatid="105322" lane="9" entrytime="00:01:50.00" />
                <RESULT eventid="99409" points="168" reactiontime="+101" swimtime="00:00:53.37" resultid="102761" heatid="105346" lane="9" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="99059" points="132" reactiontime="+90" swimtime="00:03:03.44" resultid="102765" heatid="105239" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.72" />
                    <SPLIT distance="100" swimtime="00:01:40.44" />
                    <SPLIT distance="150" swimtime="00:02:27.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102752" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="102733" number="2" reactiontime="+67" />
                    <RELAYPOSITION athleteid="102744" number="3" reactiontime="+80" />
                    <RELAYPOSITION athleteid="102705" number="4" reactiontime="+73" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="99036" points="168" reactiontime="+72" swimtime="00:03:11.87" resultid="102762" heatid="105237" lane="3" entrytime="00:34:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.08" />
                    <SPLIT distance="100" swimtime="00:01:39.19" />
                    <SPLIT distance="150" swimtime="00:02:23.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102696" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="102718" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="102710" number="3" reactiontime="+76" />
                    <RELAYPOSITION athleteid="102739" number="4" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="99234" status="DNS" swimtime="00:00:00.00" resultid="102763" heatid="105306" lane="3" entrytime="00:02:40.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102718" number="1" />
                    <RELAYPOSITION athleteid="102726" number="2" />
                    <RELAYPOSITION athleteid="102696" number="3" />
                    <RELAYPOSITION athleteid="102753" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="99441" points="126" reactiontime="+80" swimtime="00:03:06.34" resultid="102764" heatid="105363" lane="2" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.83" />
                    <SPLIT distance="100" swimtime="00:01:38.68" />
                    <SPLIT distance="150" swimtime="00:02:21.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102739" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="102705" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="102718" number="3" reactiontime="+100" />
                    <RELAYPOSITION athleteid="102744" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" status="DNS" swimtime="00:00:00.00" resultid="102766" heatid="105159" lane="1" entrytime="00:03:40.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102710" number="1" />
                    <RELAYPOSITION athleteid="102744" number="2" />
                    <RELAYPOSITION athleteid="102752" number="3" />
                    <RELAYPOSITION athleteid="102739" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="BLR" clubid="102454" name="Grodnomk.team">
          <CONTACT email="laricheva.ira@mail.ru" name="Laricheva Irina" />
          <ATHLETES>
            <ATHLETE birthdate="1963-07-22" firstname="Irina" gender="F" lastname="LARICHEVA" nation="BLR" swrid="4875830" athleteid="102455">
              <RESULTS>
                <RESULT eventid="98777" points="347" reactiontime="+98" swimtime="00:00:33.76" resultid="102456" heatid="105119" lane="4" entrytime="00:00:31.08" entrycourse="LCM" />
                <RESULT eventid="98907" points="271" reactiontime="+92" swimtime="00:00:41.81" resultid="102457" heatid="105175" lane="7" entrytime="00:00:42.00" />
                <RESULT eventid="99154" points="238" reactiontime="+98" swimtime="00:00:40.42" resultid="102458" heatid="105260" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="99409" points="249" reactiontime="+94" swimtime="00:00:46.85" resultid="102459" heatid="105345" lane="6" entrytime="00:00:52.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-06-07" firstname="Nadzeya" gender="F" lastname="KUZMINA" nation="BLR" swrid="4776833" athleteid="102460">
              <RESULTS>
                <RESULT eventid="98777" points="170" reactiontime="+113" swimtime="00:00:42.78" resultid="102461" heatid="105114" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="98907" points="171" reactiontime="+121" swimtime="00:00:48.75" resultid="102462" heatid="105173" lane="5" entrytime="00:00:50.00" />
                <RESULT eventid="99154" points="99" reactiontime="+115" swimtime="00:00:54.08" resultid="102463" heatid="105259" lane="6" entrytime="00:00:50.00" />
                <RESULT eventid="99409" points="130" reactiontime="+88" swimtime="00:00:58.19" resultid="102464" heatid="105345" lane="8" entrytime="00:00:53.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-02-02" firstname="Yuri" gender="M" lastname="KOMOU" nation="BLR" athleteid="102465">
              <RESULTS>
                <RESULT eventid="99425" points="330" reactiontime="+99" swimtime="00:00:38.57" resultid="102466" heatid="105355" lane="8" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-09-05" firstname="Sergey" gender="M" lastname="POMELOV" nation="BLR" athleteid="102467">
              <RESULTS>
                <RESULT eventid="98798" points="304" reactiontime="+104" swimtime="00:00:31.08" resultid="102468" heatid="105134" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="102469" heatid="105356" lane="7" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-12-21" firstname="Mikhail" gender="M" lastname="BARYSEVICH" nation="BLR" swrid="4875833" athleteid="102470">
              <RESULTS>
                <RESULT eventid="98798" points="398" reactiontime="+84" swimtime="00:00:28.42" resultid="102471" heatid="105138" lane="7" entrytime="00:00:28.00" />
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="102472" heatid="105271" lane="1" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-04-02" firstname="Yauheni" gender="M" lastname="SHCHEPEL" nation="BLR" swrid="4875831" athleteid="102473">
              <RESULTS>
                <RESULT eventid="98798" points="385" reactiontime="+84" swimtime="00:00:28.74" resultid="102474" heatid="105138" lane="2" entrytime="00:00:28.00" />
                <RESULT eventid="98924" points="359" reactiontime="+87" swimtime="00:00:33.80" resultid="102475" heatid="105188" lane="5" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-04-04" firstname="Dzmitry" gender="M" lastname="CHALY" nation="BLR" swrid="4967037" athleteid="102476">
              <RESULTS>
                <RESULT eventid="98798" points="361" reactiontime="+105" swimtime="00:00:29.35" resultid="102477" heatid="105138" lane="1" entrytime="00:00:28.00" />
                <RESULT eventid="98988" points="348" reactiontime="+110" swimtime="00:01:06.66" resultid="102478" heatid="105220" lane="5" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="293" reactiontime="+108" swimtime="00:00:40.11" resultid="102479" heatid="105357" lane="0" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-05-05" firstname="Vladimir" gender="M" lastname="MISHENKO" nation="BLR" athleteid="102480">
              <RESULTS>
                <RESULT eventid="98798" points="245" reactiontime="+119" swimtime="00:00:33.41" resultid="102481" heatid="105131" lane="9" entrytime="00:00:32.00" />
                <RESULT comment="K 15" eventid="99425" reactiontime="+107" status="DSQ" swimtime="00:00:00.00" resultid="102482" heatid="105356" lane="6" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-11-24" firstname="Vadim" gender="M" lastname="DUBROUSKI" nation="BLR" athleteid="102483">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="102484" heatid="105130" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="102485" heatid="105355" lane="9" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-10-27" firstname="Pavel" gender="M" lastname="TARASHCYK" nation="BLR" athleteid="102486">
              <RESULTS>
                <RESULT eventid="99425" points="234" reactiontime="+114" swimtime="00:00:43.27" resultid="102487" heatid="105354" lane="3" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M">
              <RESULTS>
                <RESULT eventid="99250" points="388" reactiontime="+96" swimtime="00:01:56.28" resultid="103430" heatid="105308" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.00" />
                    <SPLIT distance="100" swimtime="00:01:00.28" />
                    <SPLIT distance="150" swimtime="00:01:28.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102467" number="1" reactiontime="+96" />
                    <RELAYPOSITION athleteid="102476" number="2" reactiontime="+84" />
                    <RELAYPOSITION athleteid="102473" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="102470" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99059" points="329" reactiontime="+78" swimtime="00:02:15.24" resultid="103431" heatid="105240" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                    <SPLIT distance="100" swimtime="00:01:14.26" />
                    <SPLIT distance="150" swimtime="00:01:46.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102473" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="102467" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="102470" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="102476" number="4" reactiontime="+72" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Grodno.team">
              <RESULTS>
                <RESULT eventid="98846" points="255" reactiontime="+106" swimtime="00:02:13.65" resultid="102488" heatid="105159" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                    <SPLIT distance="100" swimtime="00:01:12.28" />
                    <SPLIT distance="150" swimtime="00:01:45.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102467" number="1" reactiontime="+106" />
                    <RELAYPOSITION athleteid="102460" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="102455" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="102470" number="4" reactiontime="+63" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" points="208" reactiontime="+115" swimtime="00:02:37.55" resultid="102489" heatid="105363" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.50" />
                    <SPLIT distance="100" swimtime="00:01:30.47" />
                    <SPLIT distance="150" swimtime="00:02:10.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102460" number="1" reactiontime="+115" />
                    <RELAYPOSITION athleteid="102467" number="2" reactiontime="+80" />
                    <RELAYPOSITION athleteid="102455" number="3" reactiontime="+69" />
                    <RELAYPOSITION athleteid="102470" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MŁA" nation="POL" region="WAR" clubid="102051" name="IGAN Mława">
          <CONTACT city="Mława" name="Szlagor" phone="09621127" state="MAZ" street="Żwirki" />
          <ATHLETES>
            <ATHLETE birthdate="1971-12-24" firstname="Ewa" gender="F" lastname="SZLAGOR" nation="POL" swrid="4992760" athleteid="102052">
              <RESULTS>
                <RESULT eventid="98777" points="478" reactiontime="+87" swimtime="00:00:30.33" resultid="102053" heatid="105120" lane="4" entrytime="00:00:29.30" entrycourse="SCM" />
                <RESULT eventid="99154" status="DNS" swimtime="00:00:00.00" resultid="102054" heatid="105264" lane="2" entrytime="00:00:31.00" entrycourse="LCM" />
                <RESULT eventid="99409" points="488" reactiontime="+89" swimtime="00:00:37.44" resultid="102055" heatid="105349" lane="3" entrytime="00:00:36.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="101551" name="IKS Konstancin">
          <CONTACT name="Juchno" phone="691440213" />
          <ATHLETES>
            <ATHLETE birthdate="1969-04-11" firstname="Paweł" gender="M" lastname="OBIEDZIŃSKI" nation="POL" athleteid="101557">
              <RESULTS>
                <RESULT eventid="98798" points="419" reactiontime="+73" swimtime="00:00:27.93" resultid="101558" heatid="105138" lane="3" entrytime="00:00:28.00" />
                <RESULT eventid="98830" points="345" reactiontime="+84" swimtime="00:02:42.41" resultid="101559" heatid="105154" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                    <SPLIT distance="100" swimtime="00:01:17.06" />
                    <SPLIT distance="150" swimtime="00:02:05.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="427" reactiontime="+88" swimtime="00:01:02.25" resultid="101560" heatid="105225" lane="0" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="348" reactiontime="+76" swimtime="00:01:23.10" resultid="101561" heatid="105254" lane="1" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="352" reactiontime="+83" swimtime="00:02:24.39" resultid="101562" heatid="105302" lane="0" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                    <SPLIT distance="100" swimtime="00:01:10.24" />
                    <SPLIT distance="150" swimtime="00:01:48.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="101563" heatid="105357" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="101564" heatid="106062" lane="8" entrytime="00:05:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-10-03" firstname="Rafal" gender="M" lastname="JUCHNO" nation="POL" swrid="4992759" athleteid="102490">
              <RESULTS>
                <RESULT eventid="98798" points="340" reactiontime="+92" swimtime="00:00:29.93" resultid="102491" heatid="105133" lane="2" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT eventid="98988" points="332" reactiontime="+105" swimtime="00:01:07.71" resultid="102492" heatid="105220" lane="1" entrytime="00:01:09.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="267" reactiontime="+99" swimtime="00:01:30.69" resultid="102493" heatid="105252" lane="7" entrytime="00:01:31.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="257" reactiontime="+119" swimtime="00:02:40.29" resultid="102494" heatid="105297" lane="3" entrytime="00:03:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                    <SPLIT distance="100" swimtime="00:01:16.65" />
                    <SPLIT distance="150" swimtime="00:02:00.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="RUS" clubid="103065" name="Individualno">
          <CONTACT email="a.tervinsky@gov39.ru" name="Kaliningrad" />
          <ATHLETES>
            <ATHLETE birthdate="1962-08-02" firstname="Aida" gender="F" lastname="VILIMIENE" nation="LTU" athleteid="100090">
              <RESULTS>
                <RESULT eventid="98863" status="WDR" swimtime="00:00:00.00" resultid="100540" entrytime="00:11:56.71" />
                <RESULT eventid="99202" status="DNS" swimtime="00:00:00.00" resultid="100541" heatid="105293" lane="1" entrytime="00:02:39.68" />
                <RESULT eventid="98972" status="DNS" swimtime="00:00:00.00" resultid="100542" heatid="105210" lane="0" entrytime="00:01:13.44" />
                <RESULT eventid="99457" status="WDR" swimtime="00:00:00.00" resultid="100543" entrytime="00:05:43.01" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-01-01" firstname="Svetlana" gender="F" lastname="SMIRNOVA" nation="RUS" swrid="4992860" athleteid="103066">
              <RESULTS>
                <RESULT eventid="99409" status="DNS" swimtime="00:00:00.00" resultid="103067" heatid="105346" lane="0" entrytime="00:00:49.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-01-01" firstname="Igor" gender="M" lastname="ERSHOV" nation="RUS" athleteid="103068">
              <RESULTS>
                <RESULT eventid="98798" points="189" reactiontime="+107" swimtime="00:00:36.38" resultid="103069" heatid="105126" lane="7" entrytime="00:00:36.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-01-01" firstname="Evgeniy" gender="M" lastname="NOVIKOV" nation="RUS" athleteid="103070">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="103071" heatid="105133" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="98956" points="260" reactiontime="+91" swimtime="00:03:18.89" resultid="103072" heatid="105200" lane="4" entrytime="00:03:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.29" />
                    <SPLIT distance="100" swimtime="00:01:32.03" />
                    <SPLIT distance="150" swimtime="00:02:25.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="103073" heatid="105253" lane="5" entrytime="00:01:26.50" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="103074" heatid="105358" lane="5" entrytime="00:00:36.80" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="LAT" clubid="100547" name="KIPSALA Swimming Club Riga">
          <CONTACT email="ilse.aigare@gmail.com" name="Aigare Ilse" />
          <ATHLETES>
            <ATHLETE birthdate="1965-09-07" firstname="Ilse" gender="F" lastname="AIGARE" nation="LAT" athleteid="100548">
              <RESULTS>
                <RESULT eventid="98814" points="409" reactiontime="+90" swimtime="00:02:49.92" resultid="100549" heatid="105147" lane="9" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.20" />
                    <SPLIT distance="100" swimtime="00:01:22.62" />
                    <SPLIT distance="150" swimtime="00:02:11.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98863" points="403" reactiontime="+106" swimtime="00:11:08.07" resultid="100550" heatid="105404" lane="0" entrytime="00:11:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.16" />
                    <SPLIT distance="100" swimtime="00:01:17.85" />
                    <SPLIT distance="150" swimtime="00:02:00.12" />
                    <SPLIT distance="200" swimtime="00:02:42.73" />
                    <SPLIT distance="250" swimtime="00:03:25.35" />
                    <SPLIT distance="300" swimtime="00:04:08.38" />
                    <SPLIT distance="350" swimtime="00:04:50.99" />
                    <SPLIT distance="400" swimtime="00:05:33.83" />
                    <SPLIT distance="450" swimtime="00:06:16.46" />
                    <SPLIT distance="500" swimtime="00:06:59.03" />
                    <SPLIT distance="550" swimtime="00:07:41.38" />
                    <SPLIT distance="600" swimtime="00:08:23.78" />
                    <SPLIT distance="650" swimtime="00:09:05.73" />
                    <SPLIT distance="700" swimtime="00:09:47.78" />
                    <SPLIT distance="750" swimtime="00:10:28.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="413" reactiontime="+85" swimtime="00:02:31.59" resultid="100551" heatid="105293" lane="3" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                    <SPLIT distance="100" swimtime="00:01:13.30" />
                    <SPLIT distance="150" swimtime="00:01:53.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" status="WDR" swimtime="00:00:00.00" resultid="100552" entrytime="00:05:24.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="WIE" clubid="101988" name="KP Koziegłowy">
          <CONTACT city="Koziegłowy" email="ewaszala59@wp.pl" name="Ewa Szała" street="Osiedle Leśne 13/21" zip="62-028" />
          <ATHLETES>
            <ATHLETE birthdate="1959-03-19" firstname="Ewa" gender="F" lastname="SZAŁA" nation="POL" swrid="4302573" athleteid="101989">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters,  200 zm, 50 mot" eventid="98814" points="310" reactiontime="+98" swimtime="00:03:06.25" resultid="101990" heatid="105146" lane="0" entrytime="00:03:06.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                    <SPLIT distance="100" swimtime="00:01:26.85" />
                    <SPLIT distance="150" swimtime="00:02:22.36" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters,  200,400,800 m" eventid="98863" points="311" swimtime="00:12:08.16" resultid="101991" heatid="105405" lane="3" entrytime="00:12:25.30">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.34" />
                    <SPLIT distance="200" swimtime="00:02:57.77" />
                    <SPLIT distance="300" swimtime="00:04:30.43" />
                    <SPLIT distance="400" swimtime="00:06:02.15" />
                    <SPLIT distance="500" swimtime="00:07:32.32" />
                    <SPLIT distance="600" swimtime="00:09:04.56" />
                    <SPLIT distance="700" swimtime="00:10:36.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="291" reactiontime="+91" swimtime="00:00:40.83" resultid="101992" heatid="105175" lane="4" entrytime="00:00:40.25" />
                <RESULT comment="Rekord Polski Masters,  100,200 mot" eventid="99004" points="193" reactiontime="+107" swimtime="00:03:30.71" resultid="101993" heatid="105230" lane="2" entrytime="00:03:20.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.78" />
                    <SPLIT distance="100" swimtime="00:01:40.97" />
                    <SPLIT distance="150" swimtime="00:02:36.28" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99314" points="288" reactiontime="+99" swimtime="00:01:28.00" resultid="101994" heatid="105279" lane="3" entrytime="00:01:26.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.06" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99266" points="274" reactiontime="+105" swimtime="00:06:52.87" resultid="101995" heatid="106046" lane="2" entrytime="00:06:52.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.15" />
                    <SPLIT distance="100" swimtime="00:01:41.56" />
                    <SPLIT distance="150" swimtime="00:02:33.49" />
                    <SPLIT distance="200" swimtime="00:03:25.32" />
                    <SPLIT distance="250" swimtime="00:04:23.78" />
                    <SPLIT distance="300" swimtime="00:05:20.97" />
                    <SPLIT distance="350" swimtime="00:06:07.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="257" reactiontime="+93" swimtime="00:03:14.89" resultid="101996" heatid="105334" lane="9" entrytime="00:03:06.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.22" />
                    <SPLIT distance="100" swimtime="00:01:32.87" />
                    <SPLIT distance="150" swimtime="00:02:24.64" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99457" points="262" reactiontime="+104" swimtime="00:06:13.48" resultid="101997" heatid="106056" lane="3" entrytime="00:06:10.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.34" />
                    <SPLIT distance="100" swimtime="00:01:29.37" />
                    <SPLIT distance="150" swimtime="00:02:17.01" />
                    <SPLIT distance="200" swimtime="00:03:04.66" />
                    <SPLIT distance="250" swimtime="00:03:53.31" />
                    <SPLIT distance="300" swimtime="00:04:41.55" />
                    <SPLIT distance="350" swimtime="00:05:28.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-05-27" firstname="Krzysztof" gender="M" lastname="NOWAK" nation="POL" athleteid="101998">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="101999" heatid="105124" lane="8" entrytime="00:00:48.30" />
                <RESULT eventid="98924" status="DNS" swimtime="00:00:00.00" resultid="102000" heatid="105181" lane="2" entrytime="00:00:54.20" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="102001" heatid="105213" lane="5" entrytime="00:01:40.20" />
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="102002" heatid="105249" lane="5" entrytime="00:01:55.03" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="102004" heatid="105351" lane="3" entrytime="00:00:50.22" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-08-24" firstname="Adam" gender="M" lastname="WITKOWSKI" nation="POL" swrid="4992768" athleteid="102005">
              <RESULTS>
                <RESULT eventid="98891" status="WDR" swimtime="00:00:00.00" resultid="102006" entrytime="00:22:10.05" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="102007" heatid="105217" lane="5" entrytime="00:01:12.05" />
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="102008" heatid="105299" lane="6" entrytime="00:02:36.20" />
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="102009" entrytime="00:05:30.44" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-09-02" firstname="Stefan" gender="M" lastname="SKRZYPEK" nation="POL" swrid="4564008" athleteid="102010">
              <RESULTS>
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="102011" heatid="105152" lane="9" entrytime="00:03:10.00" />
                <RESULT eventid="98891" points="210" swimtime="00:24:23.95" resultid="102012" heatid="105423" lane="4" entrytime="00:23:30.00" />
                <RESULT eventid="98956" points="160" reactiontime="+97" swimtime="00:03:53.57" resultid="102013" heatid="105199" lane="8" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.45" />
                    <SPLIT distance="100" swimtime="00:01:51.00" />
                    <SPLIT distance="150" swimtime="00:02:51.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="139" reactiontime="+101" swimtime="00:03:35.04" resultid="102014" heatid="105234" lane="6" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.16" />
                    <SPLIT distance="100" swimtime="00:01:44.86" />
                    <SPLIT distance="150" swimtime="00:02:40.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="102015" heatid="105298" lane="0" entrytime="00:02:55.00" />
                <RESULT eventid="99282" points="166" reactiontime="+105" swimtime="00:07:23.10" resultid="102016" heatid="106050" lane="1" entrytime="00:06:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.26" />
                    <SPLIT distance="100" swimtime="00:01:44.59" />
                    <SPLIT distance="150" swimtime="00:02:44.08" />
                    <SPLIT distance="200" swimtime="00:03:44.45" />
                    <SPLIT distance="250" swimtime="00:04:46.85" />
                    <SPLIT distance="300" swimtime="00:05:51.07" />
                    <SPLIT distance="350" swimtime="00:06:37.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="138" reactiontime="+106" swimtime="00:01:36.25" resultid="102017" heatid="105328" lane="0" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="221" reactiontime="+99" swimtime="00:06:03.80" resultid="102018" heatid="106063" lane="9" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.82" />
                    <SPLIT distance="100" swimtime="00:01:25.88" />
                    <SPLIT distance="150" swimtime="00:02:13.40" />
                    <SPLIT distance="200" swimtime="00:03:00.41" />
                    <SPLIT distance="250" swimtime="00:03:47.77" />
                    <SPLIT distance="300" swimtime="00:04:33.67" />
                    <SPLIT distance="350" swimtime="00:05:19.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01910" nation="POL" region="POM" clubid="100469" name="KS Delfin Gdynia">
          <ATHLETES>
            <ATHLETE birthdate="1971-11-04" firstname="Jakub" gender="M" lastname="MAŃCZAK" nation="POL" license="101910200065" swrid="4186188" athleteid="100470">
              <RESULTS>
                <RESULT eventid="99020" points="292" reactiontime="+89" swimtime="00:02:48.06" resultid="100471" heatid="105235" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                    <SPLIT distance="100" swimtime="00:01:18.99" />
                    <SPLIT distance="150" swimtime="00:02:04.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="465" swimtime="00:00:28.94" resultid="100472" heatid="105274" lane="7" entrytime="00:00:29.50" />
                <RESULT eventid="99218" points="359" reactiontime="+73" swimtime="00:02:23.45" resultid="100473" heatid="105302" lane="8" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                    <SPLIT distance="100" swimtime="00:01:09.50" />
                    <SPLIT distance="150" swimtime="00:01:47.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="389" reactiontime="+74" swimtime="00:01:08.24" resultid="100474" heatid="105330" lane="7" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="DOL" clubid="100393" name="KS Masters Polkowice">
          <CONTACT city="Polkowice" email="bogdan.jawor@gmail.com" name="Jawor Bogdan" phone="519102742" state="DOL" street="ul.Kolejowa 6/5" zip="59-100" />
          <ATHLETES>
            <ATHLETE birthdate="1968-01-02" firstname="Pavlo" gender="M" lastname="VECHIRKO" nation="POL" athleteid="100394">
              <RESULTS>
                <RESULT eventid="98798" points="315" reactiontime="+90" swimtime="00:00:30.73" resultid="100395" heatid="105133" lane="5" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT eventid="98956" points="300" reactiontime="+98" swimtime="00:03:09.54" resultid="100396" heatid="105202" lane="2" entrytime="00:03:02.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.46" />
                    <SPLIT distance="100" swimtime="00:01:29.24" />
                    <SPLIT distance="150" swimtime="00:02:18.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="306" reactiontime="+103" swimtime="00:01:26.73" resultid="100397" heatid="105249" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="299" reactiontime="+89" swimtime="00:01:17.59" resultid="100398" heatid="105286" lane="6" entrytime="00:01:14.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="299" reactiontime="+84" swimtime="00:02:47.32" resultid="100399" heatid="105341" lane="7" entrytime="00:02:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.95" />
                    <SPLIT distance="100" swimtime="00:01:20.95" />
                    <SPLIT distance="150" swimtime="00:02:03.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WARTA" nation="POL" region="WIE" clubid="102347" name="KS Warta Poznań">
          <CONTACT city="Poznań" email="j.thiem@glos.com" name="Thiem Jacek" state="WIE" street="Os. Dębina 19 m 34" zip="61-450" />
          <ATHLETES>
            <ATHLETE birthdate="1994-07-23" firstname="Przemysław" gender="M" lastname="KUCA" nation="POL" license="100115200198" swrid="4213120" athleteid="100897">
              <RESULTS>
                <RESULT eventid="98798" points="574" reactiontime="+72" swimtime="00:00:25.16" resultid="100898" heatid="105143" lane="3" entrytime="00:00:24.55" />
                <RESULT eventid="98830" points="598" reactiontime="+70" swimtime="00:02:15.31" resultid="100899" heatid="105158" lane="5" entrytime="00:02:12.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.49" />
                    <SPLIT distance="100" swimtime="00:01:03.87" />
                    <SPLIT distance="150" swimtime="00:01:45.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="638" reactiontime="+67" swimtime="00:00:54.49" resultid="100900" heatid="105228" lane="6" entrytime="00:00:54.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="555" reactiontime="+71" swimtime="00:00:27.28" resultid="100901" heatid="105276" lane="2" entrytime="00:00:26.55" />
                <RESULT eventid="99361" points="615" reactiontime="+70" swimtime="00:00:58.58" resultid="100902" heatid="105331" lane="5" entrytime="00:00:57.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="581" reactiontime="+73" swimtime="00:04:23.66" resultid="100903" heatid="106059" lane="4" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                    <SPLIT distance="100" swimtime="00:01:02.89" />
                    <SPLIT distance="150" swimtime="00:01:37.04" />
                    <SPLIT distance="200" swimtime="00:02:11.63" />
                    <SPLIT distance="250" swimtime="00:02:44.85" />
                    <SPLIT distance="300" swimtime="00:03:19.06" />
                    <SPLIT distance="350" swimtime="00:03:51.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-02-17" firstname="Jacek" gender="M" lastname="THIEM" nation="POL" swrid="4754725" athleteid="102348">
              <RESULTS>
                <RESULT eventid="98891" points="167" swimtime="00:26:20.87" resultid="102349" heatid="105423" lane="8" entrytime="00:25:00.00" />
                <RESULT eventid="99020" points="188" reactiontime="+109" swimtime="00:03:14.44" resultid="102350" heatid="105234" lane="2" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.71" />
                    <SPLIT distance="100" swimtime="00:01:32.95" />
                    <SPLIT distance="150" swimtime="00:02:23.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="156" reactiontime="+110" swimtime="00:07:32.86" resultid="102351" heatid="106050" lane="9" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.84" />
                    <SPLIT distance="100" swimtime="00:01:41.26" />
                    <SPLIT distance="150" swimtime="00:02:44.09" />
                    <SPLIT distance="200" swimtime="00:03:45.85" />
                    <SPLIT distance="250" swimtime="00:04:52.27" />
                    <SPLIT distance="300" swimtime="00:05:55.64" />
                    <SPLIT distance="350" swimtime="00:06:46.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="192" reactiontime="+99" swimtime="00:01:26.28" resultid="102352" heatid="105327" lane="6" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="182" reactiontime="+107" swimtime="00:06:27.86" resultid="102353" heatid="106064" lane="2" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.26" />
                    <SPLIT distance="100" swimtime="00:01:32.17" />
                    <SPLIT distance="150" swimtime="00:02:22.45" />
                    <SPLIT distance="200" swimtime="00:03:12.64" />
                    <SPLIT distance="250" swimtime="00:04:02.27" />
                    <SPLIT distance="300" swimtime="00:04:51.64" />
                    <SPLIT distance="350" swimtime="00:05:40.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-27" firstname="Dariusz" gender="M" lastname="JANYGA" nation="POL" swrid="4992782" athleteid="102354">
              <RESULTS>
                <RESULT eventid="98891" points="293" swimtime="00:21:50.74" resultid="102355" heatid="105421" lane="0" entrytime="00:21:20.00" />
                <RESULT eventid="98924" points="347" reactiontime="+98" swimtime="00:00:34.21" resultid="102356" heatid="105187" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="98988" points="355" reactiontime="+80" swimtime="00:01:06.23" resultid="102357" heatid="105222" lane="5" entrytime="00:01:04.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="311" reactiontime="+87" swimtime="00:01:16.63" resultid="102358" heatid="105286" lane="7" entrytime="00:01:14.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="310" reactiontime="+96" swimtime="00:02:45.21" resultid="102359" heatid="105341" lane="6" entrytime="00:02:40.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.48" />
                    <SPLIT distance="100" swimtime="00:01:22.47" />
                    <SPLIT distance="150" swimtime="00:02:05.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-19" firstname="Przemysław" gender="M" lastname="WARACZEWSKI" nation="POL" swrid="4992781" athleteid="102360">
              <RESULTS>
                <RESULT eventid="98830" points="251" reactiontime="+85" swimtime="00:03:00.63" resultid="102361" heatid="105153" lane="3" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.51" />
                    <SPLIT distance="100" swimtime="00:01:28.77" />
                    <SPLIT distance="150" swimtime="00:02:19.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="303" swimtime="00:03:08.98" resultid="102362" heatid="105201" lane="7" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.27" />
                    <SPLIT distance="100" swimtime="00:01:30.28" />
                    <SPLIT distance="150" swimtime="00:02:19.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="288" reactiontime="+84" swimtime="00:01:28.43" resultid="102363" heatid="105253" lane="1" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="186" reactiontime="+73" swimtime="00:01:30.92" resultid="102364" heatid="105284" lane="9" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="322" reactiontime="+85" swimtime="00:00:38.89" resultid="102365" heatid="105355" lane="2" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-07-02" firstname="Tomasz" gender="M" lastname="TOMASZEWSKI" nation="POL" swrid="4992783" athleteid="102366">
              <RESULTS>
                <RESULT eventid="98798" points="432" reactiontime="+83" swimtime="00:00:27.64" resultid="102367" heatid="105140" lane="4" entrytime="00:00:27.00" />
                <RESULT eventid="98924" points="475" reactiontime="+76" swimtime="00:00:30.79" resultid="102368" heatid="105189" lane="5" entrytime="00:00:30.50" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="102369" heatid="105227" lane="8" entrytime="00:00:58.00" />
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="102370" heatid="105273" lane="1" entrytime="00:00:30.00" />
                <RESULT eventid="99186" points="451" reactiontime="+80" swimtime="00:01:07.69" resultid="102371" heatid="105287" lane="7" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="367" reactiontime="+88" swimtime="00:02:36.21" resultid="102372" heatid="105341" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="100" swimtime="00:01:14.92" />
                    <SPLIT distance="150" swimtime="00:01:56.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-05-14" firstname="Przemysław" gender="M" lastname="ISALSKI" nation="POL" swrid="4048170" athleteid="102373">
              <RESULTS>
                <RESULT eventid="98830" points="399" reactiontime="+84" swimtime="00:02:34.84" resultid="102374" heatid="105152" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                    <SPLIT distance="100" swimtime="00:01:12.82" />
                    <SPLIT distance="150" swimtime="00:01:58.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="418" swimtime="00:19:24.60" resultid="102375" heatid="105420" lane="7" entrytime="00:19:30.00" />
                <RESULT eventid="98956" points="387" reactiontime="+89" swimtime="00:02:54.23" resultid="102376" heatid="105201" lane="2" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.31" />
                    <SPLIT distance="100" swimtime="00:01:23.57" />
                    <SPLIT distance="150" swimtime="00:02:09.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="395" reactiontime="+87" swimtime="00:01:03.90" resultid="102377" heatid="105222" lane="1" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="422" reactiontime="+88" swimtime="00:02:15.94" resultid="102378" heatid="105303" lane="2" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                    <SPLIT distance="100" swimtime="00:01:05.60" />
                    <SPLIT distance="150" swimtime="00:01:40.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="391" reactiontime="+93" swimtime="00:05:33.39" resultid="102379" heatid="106053" lane="1" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                    <SPLIT distance="100" swimtime="00:01:16.24" />
                    <SPLIT distance="150" swimtime="00:02:01.80" />
                    <SPLIT distance="200" swimtime="00:02:45.29" />
                    <SPLIT distance="250" swimtime="00:03:32.25" />
                    <SPLIT distance="300" swimtime="00:04:19.45" />
                    <SPLIT distance="350" swimtime="00:04:57.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="417" reactiontime="+76" swimtime="00:00:35.68" resultid="102380" heatid="105360" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="99473" points="446" reactiontime="+82" swimtime="00:04:47.97" resultid="102381" heatid="106061" lane="8" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                    <SPLIT distance="100" swimtime="00:01:10.15" />
                    <SPLIT distance="150" swimtime="00:01:47.09" />
                    <SPLIT distance="200" swimtime="00:02:24.00" />
                    <SPLIT distance="250" swimtime="00:03:00.61" />
                    <SPLIT distance="300" swimtime="00:03:36.97" />
                    <SPLIT distance="350" swimtime="00:04:12.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-02" firstname="Paweł" gender="M" lastname="OLSZEWSKI" nation="POL" swrid="4877616" athleteid="102382">
              <RESULTS>
                <RESULT eventid="98798" points="415" reactiontime="+72" swimtime="00:00:28.03" resultid="102383" heatid="105137" lane="8" entrytime="00:00:28.50" />
                <RESULT eventid="98988" points="464" reactiontime="+75" swimtime="00:01:00.56" resultid="102384" heatid="105225" lane="8" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="422" reactiontime="+82" swimtime="00:02:15.92" resultid="102385" heatid="105303" lane="6" entrytime="00:02:14.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                    <SPLIT distance="100" swimtime="00:01:07.24" />
                    <SPLIT distance="150" swimtime="00:01:42.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="435" reactiontime="+82" swimtime="00:04:50.31" resultid="102386" heatid="106061" lane="5" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                    <SPLIT distance="100" swimtime="00:01:10.27" />
                    <SPLIT distance="150" swimtime="00:01:48.10" />
                    <SPLIT distance="200" swimtime="00:02:26.38" />
                    <SPLIT distance="250" swimtime="00:03:04.21" />
                    <SPLIT distance="300" swimtime="00:03:40.55" />
                    <SPLIT distance="350" swimtime="00:04:15.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-04-28" firstname="Kamila" gender="F" lastname="OLSZEWSKA" nation="POL" athleteid="102387">
              <RESULTS>
                <RESULT eventid="98777" points="193" reactiontime="+94" swimtime="00:00:41.06" resultid="102388" heatid="105116" lane="0" entrytime="00:00:36.50" />
                <RESULT eventid="98907" status="DNS" swimtime="00:00:00.00" resultid="102389" heatid="105174" lane="2" entrytime="00:00:45.00" />
                <RESULT eventid="98972" status="DNS" swimtime="00:00:00.00" resultid="102390" heatid="105208" lane="5" entrytime="00:01:18.00" />
                <RESULT eventid="99409" status="DNS" swimtime="00:00:00.00" resultid="102391" heatid="105346" lane="8" entrytime="00:00:49.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-22" firstname="Piotr" gender="M" lastname="BURZYŃSKI" nation="POL" athleteid="102392">
              <RESULTS>
                <RESULT eventid="98891" points="228" swimtime="00:23:45.23" resultid="102393" heatid="105422" lane="1" entrytime="00:22:35.00" />
                <RESULT eventid="98956" points="175" reactiontime="+129" swimtime="00:03:46.78" resultid="102394" heatid="105199" lane="1" entrytime="00:03:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.30" />
                    <SPLIT distance="100" swimtime="00:01:48.08" />
                    <SPLIT distance="150" swimtime="00:02:47.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="102" reactiontime="+130" swimtime="00:03:58.05" resultid="102395" heatid="105233" lane="5" entrytime="00:03:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.60" />
                    <SPLIT distance="100" swimtime="00:01:51.38" />
                    <SPLIT distance="150" swimtime="00:02:55.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="163" reactiontime="+120" swimtime="00:07:25.57" resultid="102396" heatid="106051" lane="1" entrytime="00:06:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.29" />
                    <SPLIT distance="100" swimtime="00:01:51.30" />
                    <SPLIT distance="150" swimtime="00:02:53.17" />
                    <SPLIT distance="200" swimtime="00:03:53.77" />
                    <SPLIT distance="250" swimtime="00:04:52.31" />
                    <SPLIT distance="300" swimtime="00:05:52.21" />
                    <SPLIT distance="350" swimtime="00:06:39.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="219" reactiontime="+115" swimtime="00:06:04.75" resultid="102397" heatid="106064" lane="6" entrytime="00:05:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.06" />
                    <SPLIT distance="100" swimtime="00:01:24.58" />
                    <SPLIT distance="150" swimtime="00:02:11.33" />
                    <SPLIT distance="200" swimtime="00:02:58.37" />
                    <SPLIT distance="250" swimtime="00:03:45.48" />
                    <SPLIT distance="300" swimtime="00:04:32.43" />
                    <SPLIT distance="350" swimtime="00:05:19.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99059" points="283" reactiontime="+89" swimtime="00:02:22.22" resultid="102398" heatid="105240" lane="4" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="100" swimtime="00:01:14.68" />
                    <SPLIT distance="150" swimtime="00:01:54.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102354" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="102360" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="102348" number="3" reactiontime="+82" />
                    <RELAYPOSITION athleteid="102382" number="4" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="99250" points="302" reactiontime="+89" swimtime="00:02:06.41" resultid="102399" heatid="105309" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.45" />
                    <SPLIT distance="100" swimtime="00:01:08.50" />
                    <SPLIT distance="150" swimtime="00:01:38.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102360" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="102392" number="2" reactiontime="+81" />
                    <RELAYPOSITION athleteid="102354" number="3" reactiontime="+74" />
                    <RELAYPOSITION athleteid="102382" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="NZWAW" nation="POL" clubid="101155" name="KS niezrzeszeni.pl">
          <CONTACT email="niezrzeszenipl@gmail.com" internet="niezrzeszeni.pl" name="Wawer Matylda Katarzyna" phone="505960036" />
          <ATHLETES>
            <ATHLETE birthdate="1959-12-27" firstname="Wojciech" gender="M" lastname="KORPETTA" nation="POL" swrid="4754654" athleteid="101156">
              <RESULTS>
                <RESULT eventid="98830" points="163" reactiontime="+133" swimtime="00:03:28.47" resultid="101157" heatid="105148" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.38" />
                    <SPLIT distance="100" swimtime="00:01:42.17" />
                    <SPLIT distance="150" swimtime="00:02:42.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="172" swimtime="00:26:03.92" resultid="101158" heatid="105424" lane="6" entrytime="00:27:00.00" />
                <RESULT eventid="98924" points="181" reactiontime="+76" swimtime="00:00:42.48" resultid="101159" heatid="105180" lane="7" />
                <RESULT eventid="98956" points="150" reactiontime="+133" swimtime="00:03:58.82" resultid="101160" heatid="105198" lane="9" entrytime="00:03:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.86" />
                    <SPLIT distance="100" swimtime="00:01:55.41" />
                    <SPLIT distance="150" swimtime="00:02:57.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="175" reactiontime="+91" swimtime="00:03:20.00" resultid="101161" heatid="105338" lane="1" entrytime="00:03:21.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.16" />
                    <SPLIT distance="100" swimtime="00:01:38.77" />
                    <SPLIT distance="150" swimtime="00:02:31.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="171" reactiontime="+134" swimtime="00:06:36.15" resultid="101162" heatid="106065" lane="7" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.52" />
                    <SPLIT distance="100" swimtime="00:01:32.95" />
                    <SPLIT distance="150" swimtime="00:02:23.11" />
                    <SPLIT distance="200" swimtime="00:03:15.61" />
                    <SPLIT distance="250" swimtime="00:04:08.12" />
                    <SPLIT distance="300" swimtime="00:05:00.22" />
                    <SPLIT distance="350" swimtime="00:05:52.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="100332" name="KSZO MOSiR Ostrowiec Św.">
          <CONTACT email="basen@mosir.ostrowiec.pl" name="Różalski" street="Józef" />
          <ATHLETES>
            <ATHLETE birthdate="1945-03-28" firstname="Józef" gender="M" lastname="RÓŻALSKI" nation="POL" swrid="4216999" athleteid="100348">
              <RESULTS>
                <RESULT eventid="98798" points="263" reactiontime="+90" swimtime="00:00:32.60" resultid="100349" heatid="105129" lane="5" entrytime="00:00:32.50" />
                <RESULT eventid="98830" points="172" reactiontime="+86" swimtime="00:03:24.80" resultid="100350" heatid="105151" lane="9" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.86" />
                    <SPLIT distance="100" swimtime="00:01:42.64" />
                    <SPLIT distance="150" swimtime="00:02:42.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="184" reactiontime="+101" swimtime="00:03:43.12" resultid="100351" heatid="105198" lane="2" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.93" />
                    <SPLIT distance="100" swimtime="00:01:49.35" />
                    <SPLIT distance="150" swimtime="00:02:48.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="98" reactiontime="+92" swimtime="00:04:01.51" resultid="100352" heatid="105233" lane="8" entrytime="00:03:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.56" />
                    <SPLIT distance="100" swimtime="00:01:55.63" />
                    <SPLIT distance="150" swimtime="00:03:02.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="244" swimtime="00:00:35.85" resultid="100353" heatid="105269" lane="7" entrytime="00:00:35.30" />
                <RESULT eventid="99282" points="145" reactiontime="+95" swimtime="00:07:43.78" resultid="100354" heatid="106049" lane="7" entrytime="00:07:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.83" />
                    <SPLIT distance="100" swimtime="00:01:47.61" />
                    <SPLIT distance="150" swimtime="00:02:50.90" />
                    <SPLIT distance="200" swimtime="00:03:55.57" />
                    <SPLIT distance="250" swimtime="00:04:59.40" />
                    <SPLIT distance="300" swimtime="00:06:03.55" />
                    <SPLIT distance="350" swimtime="00:06:55.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="136" reactiontime="+104" swimtime="00:01:36.83" resultid="100355" heatid="105326" lane="2" entrytime="00:01:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="247" reactiontime="+100" swimtime="00:00:42.46" resultid="100356" heatid="105354" lane="6" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="UAMPO" nation="POL" region="WIE" clubid="101115" name="KU AZS UAM Poznań">
          <CONTACT city="Poznań" email="bartekz009@wp.pl" name="Ziemniarski Bartosz" phone="691679381" state="WLKP" street="Bukowska 96/1" zip="60-396" />
          <ATHLETES>
            <ATHLETE birthdate="1977-03-14" firstname="Jarosław" gender="M" lastname="BYSTRY" nation="POL" swrid="4754758" athleteid="101131">
              <RESULTS>
                <RESULT eventid="98798" points="399" reactiontime="+86" swimtime="00:00:28.38" resultid="101132" heatid="105136" lane="5" entrytime="00:00:28.80" entrycourse="LCM" />
                <RESULT eventid="98988" points="402" reactiontime="+74" swimtime="00:01:03.56" resultid="101133" heatid="105223" lane="9" entrytime="00:01:03.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="305" reactiontime="+84" swimtime="00:02:31.49" resultid="101134" heatid="105301" lane="6" entrytime="00:02:24.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.69" />
                    <SPLIT distance="100" swimtime="00:01:12.78" />
                    <SPLIT distance="150" swimtime="00:01:52.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="289" reactiontime="+91" swimtime="00:05:32.66" resultid="101135" heatid="106062" lane="1" entrytime="00:05:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.92" />
                    <SPLIT distance="100" swimtime="00:01:15.36" />
                    <SPLIT distance="150" swimtime="00:01:57.38" />
                    <SPLIT distance="200" swimtime="00:02:40.92" />
                    <SPLIT distance="250" swimtime="00:03:24.94" />
                    <SPLIT distance="300" swimtime="00:04:09.22" />
                    <SPLIT distance="350" swimtime="00:04:52.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-04-18" firstname="Karolina" gender="F" lastname="STADNIK" nation="POL" license="103315100003" swrid="4060759" athleteid="101136">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski Masters" eventid="98777" points="610" reactiontime="+80" swimtime="00:00:27.98" resultid="101137" heatid="105121" lane="4" entrytime="00:00:27.48" entrycourse="LCM" />
                <RESULT eventid="98863" points="434" reactiontime="+89" swimtime="00:10:52.24" resultid="101138" heatid="105404" lane="6" entrytime="00:10:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                    <SPLIT distance="100" swimtime="00:01:11.23" />
                    <SPLIT distance="150" swimtime="00:01:50.00" />
                    <SPLIT distance="200" swimtime="00:02:29.75" />
                    <SPLIT distance="250" swimtime="00:03:09.78" />
                    <SPLIT distance="300" swimtime="00:03:50.37" />
                    <SPLIT distance="350" swimtime="00:04:31.68" />
                    <SPLIT distance="400" swimtime="00:05:13.19" />
                    <SPLIT distance="450" swimtime="00:05:54.77" />
                    <SPLIT distance="500" swimtime="00:06:36.54" />
                    <SPLIT distance="550" swimtime="00:07:18.84" />
                    <SPLIT distance="600" swimtime="00:08:01.68" />
                    <SPLIT distance="650" swimtime="00:08:44.64" />
                    <SPLIT distance="700" swimtime="00:09:27.33" />
                    <SPLIT distance="750" swimtime="00:10:10.53" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters, Rekord Polski Masters" eventid="98907" points="547" reactiontime="+83" swimtime="00:00:33.07" resultid="101139" heatid="105178" lane="2" entrytime="00:00:33.74" entrycourse="LCM" />
                <RESULT comment="Rekord Polski Masters" eventid="98972" points="594" reactiontime="+80" swimtime="00:01:01.93" resultid="101140" heatid="105212" lane="4" entrytime="00:01:00.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.62" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99202" points="531" reactiontime="+84" swimtime="00:02:19.45" resultid="101141" heatid="105294" lane="5" entrytime="00:02:14.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                    <SPLIT distance="100" swimtime="00:01:05.20" />
                    <SPLIT distance="150" swimtime="00:01:42.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="472" reactiontime="+88" swimtime="00:05:07.11" resultid="101142" heatid="106054" lane="3" entrytime="00:04:59.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                    <SPLIT distance="100" swimtime="00:01:10.36" />
                    <SPLIT distance="150" swimtime="00:01:49.39" />
                    <SPLIT distance="200" swimtime="00:02:29.26" />
                    <SPLIT distance="250" swimtime="00:03:08.90" />
                    <SPLIT distance="300" swimtime="00:03:49.31" />
                    <SPLIT distance="350" swimtime="00:04:29.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Jakub" gender="M" lastname="STERCZYŃSKI" nation="POL" license="103315200002" swrid="4061214" athleteid="101143">
              <RESULTS>
                <RESULT eventid="98830" points="529" reactiontime="+84" swimtime="00:02:20.95" resultid="101144" heatid="105158" lane="3" entrytime="00:02:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.63" />
                    <SPLIT distance="100" swimtime="00:01:04.61" />
                    <SPLIT distance="150" swimtime="00:01:45.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="504" reactiontime="+73" swimtime="00:00:30.20" resultid="101145" heatid="105190" lane="8" entrytime="00:00:29.90" entrycourse="LCM" />
                <RESULT eventid="99186" points="498" reactiontime="+80" swimtime="00:01:05.50" resultid="101146" heatid="105288" lane="2" entrytime="00:01:03.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="482" reactiontime="+77" swimtime="00:05:10.86" resultid="101147" heatid="106053" lane="4" entrytime="00:05:05.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.17" />
                    <SPLIT distance="100" swimtime="00:01:06.88" />
                    <SPLIT distance="150" swimtime="00:01:47.47" />
                    <SPLIT distance="200" swimtime="00:02:27.20" />
                    <SPLIT distance="250" swimtime="00:03:10.68" />
                    <SPLIT distance="300" swimtime="00:03:55.23" />
                    <SPLIT distance="350" swimtime="00:04:33.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="471" reactiontime="+76" swimtime="00:02:23.84" resultid="101148" heatid="105343" lane="5" entrytime="00:02:19.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                    <SPLIT distance="100" swimtime="00:01:08.96" />
                    <SPLIT distance="150" swimtime="00:01:46.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-09-22" firstname="Bartosz" gender="M" lastname="ZIEMNIARSKI" nation="POL" license="103315200001" swrid="4061212" athleteid="101149">
              <RESULTS>
                <RESULT eventid="98798" points="547" reactiontime="+81" swimtime="00:00:25.56" resultid="101150" heatid="105143" lane="2" entrytime="00:00:24.69" entrycourse="LCM" />
                <RESULT eventid="98988" points="605" reactiontime="+80" swimtime="00:00:55.46" resultid="101151" heatid="105228" lane="3" entrytime="00:00:54.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="526" reactiontime="+89" swimtime="00:00:27.77" resultid="101152" heatid="105275" lane="2" entrytime="00:00:27.69" entrycourse="LCM" />
                <RESULT eventid="99218" points="582" reactiontime="+77" swimtime="00:02:02.10" resultid="101153" heatid="105305" lane="5" entrytime="00:02:03.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.20" />
                    <SPLIT distance="100" swimtime="00:00:59.03" />
                    <SPLIT distance="150" swimtime="00:01:30.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="527" reactiontime="+79" swimtime="00:04:32.38" resultid="101154" heatid="106059" lane="6" entrytime="00:04:31.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.78" />
                    <SPLIT distance="100" swimtime="00:01:01.31" />
                    <SPLIT distance="150" swimtime="00:01:35.47" />
                    <SPLIT distance="200" swimtime="00:02:10.62" />
                    <SPLIT distance="250" swimtime="00:02:45.85" />
                    <SPLIT distance="300" swimtime="00:03:21.46" />
                    <SPLIT distance="350" swimtime="00:03:56.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="LTU" clubid="101376" name="Kaisiadoriu p.k.PLAUKIAM">
          <CONTACT email="alex@gedwood.eu" name="Raimondas Gincas" phone="+37065609220" street="Gedimino, 8-82" />
          <ATHLETES>
            <ATHLETE birthdate="1971-04-22" firstname="Aleksandras" gender="M" lastname="ZAMORSKIS" nation="LTU" swrid="4776503" athleteid="101400">
              <RESULTS>
                <RESULT eventid="98798" points="483" reactiontime="+68" swimtime="00:00:26.65" resultid="101401" heatid="105142" lane="8" entrytime="00:00:26.00" entrycourse="LCM" />
                <RESULT eventid="98830" points="497" reactiontime="+79" swimtime="00:02:23.90" resultid="101402" heatid="105158" lane="7" entrytime="00:02:21.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.15" />
                    <SPLIT distance="100" swimtime="00:01:07.42" />
                    <SPLIT distance="150" swimtime="00:01:50.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="542" reactiontime="+73" swimtime="00:00:57.50" resultid="101403" heatid="105227" lane="6" entrytime="00:00:57.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="524" reactiontime="+71" swimtime="00:01:12.48" resultid="101404" heatid="105257" lane="4" entrytime="00:01:13.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="461" reactiontime="+66" swimtime="00:01:07.20" resultid="101405" heatid="105288" lane="9" entrytime="00:01:08.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="454" reactiontime="+80" swimtime="00:01:04.79" resultid="101406" heatid="105330" lane="5" entrytime="00:01:04.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-07-20" firstname="Raimondas" gender="M" lastname="GINCAS" nation="LTU" swrid="4317387" athleteid="101407">
              <RESULTS>
                <RESULT eventid="98891" points="337" swimtime="00:20:51.51" resultid="101408" heatid="105420" lane="9" entrytime="00:20:00.00" />
                <RESULT eventid="98988" points="484" reactiontime="+69" swimtime="00:00:59.72" resultid="101409" heatid="105227" lane="9" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="431" reactiontime="+76" swimtime="00:02:15.00" resultid="101410" heatid="105304" lane="6" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                    <SPLIT distance="100" swimtime="00:01:06.32" />
                    <SPLIT distance="150" swimtime="00:01:40.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="409" reactiontime="+82" swimtime="00:04:56.26" resultid="101411" heatid="106060" lane="5" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.97" />
                    <SPLIT distance="100" swimtime="00:01:12.32" />
                    <SPLIT distance="150" swimtime="00:01:50.84" />
                    <SPLIT distance="200" swimtime="00:02:29.15" />
                    <SPLIT distance="250" swimtime="00:03:06.59" />
                    <SPLIT distance="300" swimtime="00:03:45.01" />
                    <SPLIT distance="350" swimtime="00:04:21.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-05-01" firstname="Mindaugas" gender="M" lastname="SAKYS" nation="LTU" swrid="4776502" athleteid="101412">
              <RESULTS>
                <RESULT eventid="98830" points="390" reactiontime="+90" swimtime="00:02:35.93" resultid="101413" heatid="105156" lane="5" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                    <SPLIT distance="100" swimtime="00:01:12.60" />
                    <SPLIT distance="150" swimtime="00:01:58.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="372" reactiontime="+79" swimtime="00:00:33.40" resultid="101414" heatid="105187" lane="7" entrytime="00:00:34.00" />
                <RESULT eventid="99186" points="377" reactiontime="+78" swimtime="00:01:11.88" resultid="101415" heatid="105287" lane="3" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="362" reactiontime="+77" swimtime="00:02:37.02" resultid="101416" heatid="105342" lane="0" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                    <SPLIT distance="100" swimtime="00:01:15.00" />
                    <SPLIT distance="150" swimtime="00:01:56.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-01-14" firstname="Eimantas" gender="M" lastname="FRANKONIS" nation="LTU" athleteid="101417">
              <RESULTS>
                <RESULT eventid="98798" points="374" reactiontime="+80" swimtime="00:00:29.01" resultid="101418" heatid="105136" lane="9" entrytime="00:00:29.00" />
                <RESULT eventid="98956" points="330" reactiontime="+68" swimtime="00:03:03.77" resultid="101419" heatid="105203" lane="8" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.19" />
                    <SPLIT distance="100" swimtime="00:01:27.06" />
                    <SPLIT distance="150" swimtime="00:02:15.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="379" reactiontime="+74" swimtime="00:01:20.75" resultid="101420" heatid="105256" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="364" reactiontime="+83" swimtime="00:00:37.32" resultid="101421" heatid="105360" lane="6" entrytime="00:00:34.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-08-22" firstname="Gintas" gender="M" lastname="KANAPICKAS" nation="LTU" swrid="4776500" athleteid="101422">
              <RESULTS>
                <RESULT comment="04" eventid="98798" reactiontime="+74" status="DSQ" swimtime="00:00:31.81" resultid="101423" heatid="105132" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="98988" points="281" reactiontime="+77" swimtime="00:01:11.54" resultid="101424" heatid="105219" lane="8" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="101425" heatid="105300" lane="7" entrytime="00:02:30.00" />
                <RESULT eventid="99393" points="217" reactiontime="+101" swimtime="00:03:05.98" resultid="101426" heatid="105339" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.86" />
                    <SPLIT distance="100" swimtime="00:01:29.67" />
                    <SPLIT distance="150" swimtime="00:02:18.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99250" points="463" reactiontime="+76" swimtime="00:01:49.66" resultid="101428" heatid="105311" lane="6" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.39" />
                    <SPLIT distance="100" swimtime="00:00:56.75" />
                    <SPLIT distance="150" swimtime="00:01:22.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101417" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="101412" number="2" reactiontime="+38" />
                    <RELAYPOSITION athleteid="101400" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="101407" number="4" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="99059" points="431" reactiontime="+70" swimtime="00:02:03.62" resultid="105085" heatid="105239" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                    <SPLIT distance="100" swimtime="00:01:09.00" />
                    <SPLIT distance="150" swimtime="00:01:36.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101412" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="101417" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="101400" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="101407" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="102075" name="Legia Warszawa">
          <CONTACT email="sekcja@plywanielegia.pl" name="Drzewiński" phone="600826305" />
          <ATHLETES>
            <ATHLETE birthdate="1990-06-24" firstname="Michał" gender="M" lastname="CHOIŃSKI" nation="POL" swrid="4071732" athleteid="102408">
              <RESULTS>
                <RESULT eventid="98798" points="492" reactiontime="+74" swimtime="00:00:26.48" resultid="102409" heatid="105142" lane="5" entrytime="00:00:25.50" />
                <RESULT eventid="98924" points="458" reactiontime="+63" swimtime="00:00:31.17" resultid="102410" heatid="105190" lane="3" entrytime="00:00:28.80" />
                <RESULT eventid="99170" points="570" reactiontime="+74" swimtime="00:00:27.04" resultid="102411" heatid="105276" lane="6" entrytime="00:00:26.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-09-01" firstname="Agata" gender="F" lastname="LESZCZYŃSKA" nation="POL" swrid="4806426" athleteid="102412">
              <RESULTS>
                <RESULT eventid="98777" points="504" reactiontime="+76" swimtime="00:00:29.80" resultid="102413" heatid="105120" lane="7" entrytime="00:00:30.25" entrycourse="LCM" />
                <RESULT eventid="98907" points="476" reactiontime="+74" swimtime="00:00:34.65" resultid="102414" heatid="105178" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="98972" status="DNS" swimtime="00:00:00.00" resultid="102415" heatid="105212" lane="6" entrytime="00:01:01.00" />
                <RESULT eventid="99154" points="456" swimtime="00:00:32.57" resultid="102416" heatid="105264" lane="7" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-03-18" firstname="Maciej" gender="M" lastname="PASIECZNY" nation="POL" swrid="4071778" athleteid="102417">
              <RESULTS>
                <RESULT eventid="98798" points="437" reactiontime="+70" swimtime="00:00:27.55" resultid="102418" heatid="105143" lane="9" entrytime="00:00:25.00" />
                <RESULT eventid="98988" points="474" reactiontime="+70" swimtime="00:01:00.14" resultid="102419" heatid="105228" lane="8" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="485" reactiontime="+77" swimtime="00:00:28.54" resultid="102420" heatid="105276" lane="1" entrytime="00:00:27.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-10-24" firstname="Marcin" gender="M" lastname="WILCZĘGA" nation="POL" swrid="4992879" athleteid="102812">
              <RESULTS>
                <RESULT eventid="98798" points="437" reactiontime="+78" swimtime="00:00:27.54" resultid="102813" heatid="105141" lane="0" entrytime="00:00:26.95" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-25" firstname="Marcin" gender="M" lastname="KACZMAREK" nation="POL" swrid="4043251" athleteid="102820">
              <RESULTS>
                <RESULT eventid="98924" points="579" reactiontime="+72" swimtime="00:00:28.84" resultid="102821" heatid="105190" lane="4" entrytime="00:00:27.10" />
                <RESULT eventid="99170" points="586" reactiontime="+86" swimtime="00:00:26.79" resultid="102822" heatid="105276" lane="3" entrytime="00:00:26.00" />
                <RESULT eventid="99186" points="560" reactiontime="+79" swimtime="00:01:03.01" resultid="102823" heatid="105288" lane="4" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99361" points="587" reactiontime="+95" swimtime="00:00:59.48" resultid="102824" heatid="105331" lane="3" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="539" reactiontime="+67" swimtime="00:02:17.52" resultid="102825" heatid="105343" lane="6" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                    <SPLIT distance="100" swimtime="00:01:07.26" />
                    <SPLIT distance="150" swimtime="00:01:43.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Krzysztof" gender="M" lastname="MICOREK" nation="POL" swrid="4086676" athleteid="102937">
              <RESULTS>
                <RESULT eventid="98798" points="551" reactiontime="+83" swimtime="00:00:25.50" resultid="103042" heatid="105143" lane="6" entrytime="00:00:24.60" />
                <RESULT eventid="98988" points="530" reactiontime="+88" swimtime="00:00:57.96" resultid="103043" heatid="105228" lane="2" entrytime="00:00:54.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="103044" heatid="105276" lane="0" entrytime="00:00:27.00" />
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="103045" heatid="105331" lane="1" entrytime="00:01:02.00" />
                <RESULT comment="            Z2" eventid="99425" reactiontime="+77" status="DSQ" swimtime="00:00:00.00" resultid="103046" heatid="105362" lane="5" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MKPIA" nation="POL" region="WAR" clubid="102523" name="MKS Piaseczno">
          <CONTACT city="PIASECZNO" name="ANDRZEJ RUBASZKIEWICZ" />
          <ATHLETES>
            <ATHLETE birthdate="1949-04-10" firstname="Andrzej" gender="M" lastname="RUBASZKIEWICZ" nation="POL" license="SO6414200002" swrid="4340487" athleteid="102524">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski Masters" eventid="98798" points="320" reactiontime="+74" swimtime="00:00:30.55" resultid="102525" heatid="105134" lane="8" entrytime="00:00:30.00" />
                <RESULT comment="Rekord Polski Masters, Rekord Polski Masters" eventid="98924" points="246" reactiontime="+89" swimtime="00:00:38.36" resultid="102526" heatid="105185" lane="3" entrytime="00:00:38.00" />
                <RESULT comment="Rekord Polski Masters" eventid="98988" points="315" reactiontime="+90" swimtime="00:01:08.88" resultid="102527" heatid="105221" lane="3" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="309" reactiontime="+86" swimtime="00:00:33.17" resultid="102528" heatid="105270" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="99218" points="233" reactiontime="+101" swimtime="00:02:45.63" resultid="102529" heatid="105300" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                    <SPLIT distance="100" swimtime="00:01:19.85" />
                    <SPLIT distance="150" swimtime="00:02:04.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="182" reactiontime="+89" swimtime="00:01:27.79" resultid="102530" heatid="105327" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOTYL" nation="POL" clubid="100737" name="MOTYL SENIOR MOSiR Stalowa Wola" shortname="MOTYL Stalowa W.">
          <CONTACT city="Stalowa Wola" email="lorkowska@wp.pl" name="Chmielewski Andrzej" street="Hutnicza 15" zip="37-450" />
          <ATHLETES>
            <ATHLETE birthdate="1975-03-19" firstname="Robert" gender="M" lastname="BARAN" nation="POL" swrid="4992836" athleteid="100750">
              <RESULTS>
                <RESULT eventid="98798" points="459" reactiontime="+83" swimtime="00:00:27.09" resultid="100751" heatid="105141" lane="8" entrytime="00:00:26.67" />
                <RESULT eventid="98830" points="418" reactiontime="+95" swimtime="00:02:32.38" resultid="100752" heatid="105155" lane="4" entrytime="00:02:39.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                    <SPLIT distance="100" swimtime="00:01:10.43" />
                    <SPLIT distance="150" swimtime="00:01:56.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="479" reactiontime="+75" swimtime="00:00:30.71" resultid="100753" heatid="105189" lane="7" entrytime="00:00:31.07" />
                <RESULT eventid="98988" points="467" reactiontime="+102" swimtime="00:01:00.46" resultid="100754" heatid="105225" lane="1" entrytime="00:01:00.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="451" reactiontime="+74" swimtime="00:01:07.71" resultid="100755" heatid="105287" lane="4" entrytime="00:01:08.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="335" reactiontime="+93" swimtime="00:02:26.76" resultid="100756" heatid="105302" lane="5" entrytime="00:02:19.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                    <SPLIT distance="100" swimtime="00:01:09.79" />
                    <SPLIT distance="150" swimtime="00:01:48.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="378" reactiontime="+86" swimtime="00:02:34.75" resultid="100757" heatid="105342" lane="2" entrytime="00:02:32.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                    <SPLIT distance="100" swimtime="00:01:15.83" />
                    <SPLIT distance="150" swimtime="00:01:56.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="321" reactiontime="+86" swimtime="00:00:38.94" resultid="100758" heatid="105358" lane="9" entrytime="00:00:37.93" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-14" firstname="Arkadiusz" gender="M" lastname="BERWECKI" nation="POL" swrid="4791744" athleteid="100759">
              <RESULTS>
                <RESULT eventid="98798" points="495" reactiontime="+71" swimtime="00:00:26.43" resultid="100760" heatid="105141" lane="7" entrytime="00:00:26.50" />
                <RESULT eventid="98830" points="532" reactiontime="+83" swimtime="00:02:20.66" resultid="100761" heatid="105158" lane="2" entrytime="00:02:21.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.34" />
                    <SPLIT distance="100" swimtime="00:01:05.02" />
                    <SPLIT distance="150" swimtime="00:01:46.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="406" reactiontime="+71" swimtime="00:00:32.45" resultid="100762" heatid="105189" lane="9" entrytime="00:00:32.50" />
                <RESULT eventid="99020" points="423" reactiontime="+94" swimtime="00:02:28.44" resultid="100763" heatid="105236" lane="4" entrytime="00:02:21.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                    <SPLIT distance="100" swimtime="00:01:09.29" />
                    <SPLIT distance="150" swimtime="00:01:48.02" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99091" points="520" reactiontime="+82" swimtime="00:01:12.68" resultid="100764" heatid="105257" lane="3" entrytime="00:01:14.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="458" reactiontime="+94" swimtime="00:05:16.16" resultid="100765" heatid="106053" lane="2" entrytime="00:05:18.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                    <SPLIT distance="100" swimtime="00:01:10.38" />
                    <SPLIT distance="150" swimtime="00:01:50.88" />
                    <SPLIT distance="200" swimtime="00:02:31.02" />
                    <SPLIT distance="250" swimtime="00:03:16.27" />
                    <SPLIT distance="300" swimtime="00:04:01.79" />
                    <SPLIT distance="350" swimtime="00:04:39.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="545" reactiontime="+85" swimtime="00:01:00.96" resultid="100766" heatid="105331" lane="2" entrytime="00:01:01.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="419" reactiontime="+74" swimtime="00:02:29.45" resultid="100767" heatid="105342" lane="5" entrytime="00:02:30.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.36" />
                    <SPLIT distance="100" swimtime="00:01:11.74" />
                    <SPLIT distance="150" swimtime="00:01:50.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-08-09" firstname="Włodzimierz" gender="M" lastname="JARZYNA" nation="POL" swrid="4992837" athleteid="100768">
              <RESULTS>
                <RESULT eventid="98798" points="258" reactiontime="+98" swimtime="00:00:32.84" resultid="100769" heatid="105127" lane="1" entrytime="00:00:35.61" />
                <RESULT eventid="98830" points="174" reactiontime="+102" swimtime="00:03:24.11" resultid="100770" heatid="105150" lane="5" entrytime="00:03:40.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.73" />
                    <SPLIT distance="100" swimtime="00:01:40.04" />
                    <SPLIT distance="150" swimtime="00:02:41.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="176" reactiontime="+84" swimtime="00:00:42.82" resultid="100771" heatid="105183" lane="9" entrytime="00:00:45.23" />
                <RESULT eventid="98956" points="184" reactiontime="+103" swimtime="00:03:43.16" resultid="100772" heatid="105198" lane="1" entrytime="00:03:46.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.11" />
                    <SPLIT distance="100" swimtime="00:01:51.09" />
                    <SPLIT distance="150" swimtime="00:02:50.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="173" reactiontime="+93" swimtime="00:01:33.05" resultid="100773" heatid="105283" lane="0" entrytime="00:01:36.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="170" reactiontime="+97" swimtime="00:07:19.54" resultid="100774" heatid="106049" lane="3" entrytime="00:07:21.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.11" />
                    <SPLIT distance="100" swimtime="00:01:52.79" />
                    <SPLIT distance="150" swimtime="00:02:51.18" />
                    <SPLIT distance="200" swimtime="00:03:44.94" />
                    <SPLIT distance="250" swimtime="00:04:46.77" />
                    <SPLIT distance="300" swimtime="00:05:47.28" />
                    <SPLIT distance="350" swimtime="00:06:35.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="155" reactiontime="+72" swimtime="00:03:28.04" resultid="100775" heatid="105338" lane="8" entrytime="00:03:33.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.58" />
                    <SPLIT distance="100" swimtime="00:01:43.60" />
                    <SPLIT distance="150" swimtime="00:02:39.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="196" reactiontime="+106" swimtime="00:06:18.45" resultid="100776" heatid="106065" lane="6" entrytime="00:06:28.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.13" />
                    <SPLIT distance="100" swimtime="00:01:30.02" />
                    <SPLIT distance="150" swimtime="00:02:20.04" />
                    <SPLIT distance="200" swimtime="00:03:09.67" />
                    <SPLIT distance="250" swimtime="00:04:00.28" />
                    <SPLIT distance="300" swimtime="00:04:49.17" />
                    <SPLIT distance="350" swimtime="00:05:36.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-18" firstname="Waldemar" gender="M" lastname="KALBARCZYK" nation="POL" athleteid="100777">
              <RESULTS>
                <RESULT eventid="98798" points="295" reactiontime="+92" swimtime="00:00:31.41" resultid="100778" heatid="105132" lane="5" entrytime="00:00:30.72" />
                <RESULT eventid="98830" points="237" reactiontime="+85" swimtime="00:03:04.12" resultid="100779" heatid="105153" lane="8" entrytime="00:02:57.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.02" />
                    <SPLIT distance="100" swimtime="00:01:26.52" />
                    <SPLIT distance="150" swimtime="00:02:21.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="242" reactiontime="+97" swimtime="00:03:23.67" resultid="100780" heatid="105200" lane="0" entrytime="00:03:25.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.46" />
                    <SPLIT distance="100" swimtime="00:01:37.18" />
                    <SPLIT distance="150" swimtime="00:02:30.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="272" reactiontime="+87" swimtime="00:01:12.35" resultid="100781" heatid="105219" lane="4" entrytime="00:01:09.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="256" reactiontime="+92" swimtime="00:00:35.30" resultid="100782" heatid="105270" lane="1" entrytime="00:00:34.51" />
                <RESULT eventid="99282" points="237" reactiontime="+108" swimtime="00:06:33.68" resultid="100783" heatid="106050" lane="2" entrytime="00:06:45.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.29" />
                    <SPLIT distance="100" swimtime="00:01:38.14" />
                    <SPLIT distance="150" swimtime="00:02:27.66" />
                    <SPLIT distance="200" swimtime="00:03:15.91" />
                    <SPLIT distance="250" swimtime="00:04:12.68" />
                    <SPLIT distance="300" swimtime="00:05:08.38" />
                    <SPLIT distance="350" swimtime="00:05:52.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="211" reactiontime="+88" swimtime="00:03:07.74" resultid="100784" heatid="105339" lane="3" entrytime="00:02:59.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.17" />
                    <SPLIT distance="100" swimtime="00:01:29.76" />
                    <SPLIT distance="150" swimtime="00:02:19.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="248" reactiontime="+87" swimtime="00:00:42.42" resultid="100785" heatid="105355" lane="4" entrytime="00:00:41.25" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-02-27" firstname="Robert" gender="M" lastname="LORKOWSKI" nation="POL" swrid="4992838" athleteid="100786">
              <RESULTS>
                <RESULT eventid="98830" points="288" reactiontime="+92" swimtime="00:02:52.43" resultid="100787" heatid="105154" lane="0" entrytime="00:02:53.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.39" />
                    <SPLIT distance="100" swimtime="00:00:40.50" />
                    <SPLIT distance="150" swimtime="00:02:13.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="235" swimtime="00:23:29.93" resultid="100788" heatid="105423" lane="6" entrytime="00:23:40.11" />
                <RESULT eventid="98988" points="319" reactiontime="+96" swimtime="00:01:08.62" resultid="100789" heatid="105218" lane="3" entrytime="00:01:10.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="193" reactiontime="+93" swimtime="00:03:12.76" resultid="100790" heatid="105234" lane="8" entrytime="00:03:25.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.37" />
                    <SPLIT distance="100" swimtime="00:01:29.20" />
                    <SPLIT distance="150" swimtime="00:02:22.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="249" reactiontime="+95" swimtime="00:01:22.51" resultid="100791" heatid="105284" lane="2" entrytime="00:01:21.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="253" reactiontime="+92" swimtime="00:06:25.40" resultid="100792" heatid="106051" lane="9" entrytime="00:06:32.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.16" />
                    <SPLIT distance="100" swimtime="00:01:28.81" />
                    <SPLIT distance="150" swimtime="00:02:18.09" />
                    <SPLIT distance="200" swimtime="00:03:07.27" />
                    <SPLIT distance="250" swimtime="00:04:05.18" />
                    <SPLIT distance="300" swimtime="00:05:01.29" />
                    <SPLIT distance="350" swimtime="00:05:44.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="239" reactiontime="+80" swimtime="00:03:00.27" resultid="100793" heatid="105339" lane="6" entrytime="00:02:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.84" />
                    <SPLIT distance="100" swimtime="00:01:26.17" />
                    <SPLIT distance="150" swimtime="00:02:13.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="100794" heatid="106064" lane="5" entrytime="00:05:55.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-07-07" firstname="Marcin" gender="M" lastname="MUSIALIK" nation="POL" swrid="4509577" athleteid="100795">
              <RESULTS>
                <RESULT eventid="98830" points="388" reactiontime="+92" swimtime="00:02:36.23" resultid="100796" heatid="105156" lane="6" entrytime="00:02:34.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                    <SPLIT distance="100" swimtime="00:01:14.15" />
                    <SPLIT distance="150" swimtime="00:02:00.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="382" swimtime="00:19:59.98" resultid="100797" heatid="105420" lane="8" entrytime="00:19:41.21" />
                <RESULT eventid="98924" points="309" reactiontime="+76" swimtime="00:00:35.53" resultid="100798" heatid="105187" lane="4" entrytime="00:00:33.28" />
                <RESULT eventid="99020" points="290" reactiontime="+98" swimtime="00:02:48.43" resultid="100799" heatid="105235" lane="5" entrytime="00:02:42.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                    <SPLIT distance="100" swimtime="00:01:20.11" />
                    <SPLIT distance="150" swimtime="00:02:04.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="361" reactiontime="+90" swimtime="00:02:23.23" resultid="100800" heatid="105303" lane="9" entrytime="00:02:16.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                    <SPLIT distance="100" swimtime="00:01:09.98" />
                    <SPLIT distance="150" swimtime="00:01:47.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="370" reactiontime="+103" swimtime="00:05:39.36" resultid="100801" heatid="106052" lane="4" entrytime="00:05:42.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                    <SPLIT distance="100" swimtime="00:01:16.52" />
                    <SPLIT distance="150" swimtime="00:02:00.43" />
                    <SPLIT distance="200" swimtime="00:02:44.02" />
                    <SPLIT distance="250" swimtime="00:03:33.34" />
                    <SPLIT distance="300" swimtime="00:04:23.57" />
                    <SPLIT distance="350" swimtime="00:05:02.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="314" reactiontime="+66" swimtime="00:02:44.49" resultid="100802" heatid="105342" lane="7" entrytime="00:02:32.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.99" />
                    <SPLIT distance="100" swimtime="00:01:18.45" />
                    <SPLIT distance="150" swimtime="00:02:00.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="405" reactiontime="+97" swimtime="00:04:57.25" resultid="100803" heatid="106060" lane="6" entrytime="00:04:45.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                    <SPLIT distance="100" swimtime="00:01:10.39" />
                    <SPLIT distance="150" swimtime="00:01:48.18" />
                    <SPLIT distance="200" swimtime="00:02:26.59" />
                    <SPLIT distance="250" swimtime="00:03:05.10" />
                    <SPLIT distance="300" swimtime="00:03:43.83" />
                    <SPLIT distance="350" swimtime="00:04:21.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-26" firstname="Krzysztof" gender="M" lastname="PAWŁOWSKI" nation="POL" swrid="4992839" athleteid="100804">
              <RESULTS>
                <RESULT eventid="98798" points="329" reactiontime="+85" swimtime="00:00:30.27" resultid="100805" heatid="105135" lane="1" entrytime="00:00:29.50" />
                <RESULT eventid="98891" points="238" swimtime="00:23:24.92" resultid="100806" heatid="105422" lane="6" entrytime="00:22:29.50" />
                <RESULT eventid="99020" points="155" reactiontime="+99" swimtime="00:03:27.30" resultid="100808" heatid="105233" lane="4" entrytime="00:03:30.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.52" />
                    <SPLIT distance="100" swimtime="00:01:37.31" />
                    <SPLIT distance="150" swimtime="00:02:33.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="300" reactiontime="+87" swimtime="00:01:27.24" resultid="100809" heatid="105253" lane="0" entrytime="00:01:28.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="241" reactiontime="+94" swimtime="00:06:31.52" resultid="100810" heatid="106050" lane="4" entrytime="00:06:34.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.33" />
                    <SPLIT distance="100" swimtime="00:01:37.10" />
                    <SPLIT distance="150" swimtime="00:02:27.46" />
                    <SPLIT distance="200" swimtime="00:03:17.35" />
                    <SPLIT distance="250" swimtime="00:04:11.07" />
                    <SPLIT distance="300" swimtime="00:05:05.41" />
                    <SPLIT distance="350" swimtime="00:05:48.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="241" reactiontime="+86" swimtime="00:02:59.83" resultid="100811" heatid="105339" lane="8" entrytime="00:03:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.61" />
                    <SPLIT distance="100" swimtime="00:01:25.74" />
                    <SPLIT distance="150" swimtime="00:02:12.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="100812" heatid="106064" lane="3" entrytime="00:05:55.20" />
                <RESULT eventid="98956" points="281" reactiontime="+98" swimtime="00:03:13.71" resultid="101987" heatid="105201" lane="1" entrytime="00:03:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.13" />
                    <SPLIT distance="100" swimtime="00:01:29.25" />
                    <SPLIT distance="150" swimtime="00:02:20.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-04-17" firstname="Maria" gender="F" lastname="PETECKA" nation="POL" swrid="4992840" athleteid="100813">
              <RESULTS>
                <RESULT eventid="98777" points="308" reactiontime="+94" swimtime="00:00:35.12" resultid="100814" heatid="105117" lane="3" entrytime="00:00:34.40" entrycourse="SCM" />
                <RESULT eventid="98814" points="304" reactiontime="+85" swimtime="00:03:07.53" resultid="100815" heatid="105145" lane="6" entrytime="00:03:18.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.28" />
                    <SPLIT distance="100" swimtime="00:01:32.87" />
                    <SPLIT distance="150" swimtime="00:02:25.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="281" reactiontime="+87" swimtime="00:03:32.33" resultid="100816" heatid="105193" lane="8" entrytime="00:03:35.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.92" />
                    <SPLIT distance="100" swimtime="00:01:44.40" />
                    <SPLIT distance="150" swimtime="00:02:40.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99004" points="176" reactiontime="+99" swimtime="00:03:36.95" resultid="100817" heatid="105230" lane="1" entrytime="00:03:30.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.54" />
                    <SPLIT distance="100" swimtime="00:01:40.64" />
                    <SPLIT distance="150" swimtime="00:02:39.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="234" reactiontime="+99" swimtime="00:01:44.28" resultid="100818" heatid="105245" lane="0" entrytime="00:01:50.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="227" reactiontime="+91" swimtime="00:00:41.08" resultid="100819" heatid="105261" lane="6" entrytime="00:00:39.00" />
                <RESULT eventid="99344" points="211" reactiontime="+95" swimtime="00:01:34.03" resultid="100820" heatid="105322" lane="7" entrytime="00:01:35.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="257" reactiontime="+92" swimtime="00:00:46.33" resultid="100821" heatid="105346" lane="3" entrytime="00:00:46.11" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-03-12" firstname="Adam" gender="M" lastname="PRZYBYLSKI" nation="POL" swrid="4992841" athleteid="100822">
              <RESULTS>
                <RESULT eventid="98798" points="399" reactiontime="+78" swimtime="00:00:28.39" resultid="100823" heatid="105136" lane="3" entrytime="00:00:28.89" />
                <RESULT eventid="98924" points="266" reactiontime="+67" swimtime="00:00:37.34" resultid="100824" heatid="105185" lane="7" entrytime="00:00:38.72" />
                <RESULT eventid="98988" points="366" reactiontime="+87" swimtime="00:01:05.55" resultid="100825" heatid="105222" lane="2" entrytime="00:01:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="356" reactiontime="+76" swimtime="00:00:31.62" resultid="100826" heatid="105268" lane="7" entrytime="00:00:36.57" />
                <RESULT eventid="99186" points="254" reactiontime="+72" swimtime="00:01:21.95" resultid="100827" heatid="105284" lane="3" entrytime="00:01:18.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="243" reactiontime="+87" swimtime="00:01:19.78" resultid="100828" heatid="105326" lane="5" entrytime="00:01:30.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="225" reactiontime="+83" swimtime="00:03:03.81" resultid="100829" heatid="105339" lane="1" entrytime="00:03:01.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.22" />
                    <SPLIT distance="100" swimtime="00:01:29.30" />
                    <SPLIT distance="150" swimtime="00:02:17.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-04-15" firstname="Michał" gender="M" lastname="SKROK" nation="POL" swrid="4992842" athleteid="100830">
              <RESULTS>
                <RESULT eventid="98798" points="422" reactiontime="+77" swimtime="00:00:27.86" resultid="100831" heatid="105134" lane="4" entrytime="00:00:29.90" />
                <RESULT eventid="98830" points="421" reactiontime="+85" swimtime="00:02:32.02" resultid="100832" heatid="105156" lane="3" entrytime="00:02:34.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.80" />
                    <SPLIT distance="100" swimtime="00:01:14.33" />
                    <SPLIT distance="150" swimtime="00:01:56.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="412" reactiontime="+73" swimtime="00:02:50.68" resultid="100833" heatid="105203" lane="6" entrytime="00:02:55.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.80" />
                    <SPLIT distance="100" swimtime="00:01:23.23" />
                    <SPLIT distance="150" swimtime="00:02:08.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="476" reactiontime="+79" swimtime="00:01:14.83" resultid="100834" heatid="105256" lane="4" entrytime="00:01:18.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="378" reactiontime="+90" swimtime="00:05:37.10" resultid="100835" heatid="106052" lane="1" entrytime="00:05:50.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.07" />
                    <SPLIT distance="100" swimtime="00:01:17.36" />
                    <SPLIT distance="150" swimtime="00:02:03.16" />
                    <SPLIT distance="200" swimtime="00:02:47.97" />
                    <SPLIT distance="250" swimtime="00:03:34.78" />
                    <SPLIT distance="300" swimtime="00:04:21.33" />
                    <SPLIT distance="350" swimtime="00:05:00.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="507" reactiontime="+80" swimtime="00:00:33.43" resultid="100836" heatid="105361" lane="0" entrytime="00:00:34.40" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="99059" points="489" reactiontime="+77" swimtime="00:01:58.53" resultid="100837" heatid="105242" lane="5" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                    <SPLIT distance="100" swimtime="00:01:03.18" />
                    <SPLIT distance="150" swimtime="00:01:30.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100750" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="100830" number="2" reactiontime="+29" />
                    <RELAYPOSITION athleteid="100759" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="100822" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="99250" points="371" reactiontime="+91" swimtime="00:01:57.98" resultid="100838" heatid="105310" lane="6" entrytime="00:02:00.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.06" />
                    <SPLIT distance="100" swimtime="00:00:59.76" />
                    <SPLIT distance="150" swimtime="00:01:30.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100750" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="100768" number="2" reactiontime="+12" />
                    <RELAYPOSITION athleteid="100786" number="3" reactiontime="+75" />
                    <RELAYPOSITION athleteid="100822" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="LU" clubid="102070" name="MTP Lublinianka">
          <CONTACT email="thomaswim@gazeta.pl" name="Tomasz Duszynski" phone="791846627" />
          <ATHLETES>
            <ATHLETE birthdate="1976-12-17" firstname="Tomasz" gender="M" lastname="DUSZYNSKI" nation="POL" swrid="4037875" athleteid="102071">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="98956" points="582" reactiontime="+88" swimtime="00:02:32.04" resultid="102072" heatid="105204" lane="4" entrytime="00:02:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="100" swimtime="00:01:14.22" />
                    <SPLIT distance="150" swimtime="00:01:52.36" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99091" points="579" reactiontime="+89" swimtime="00:01:10.10" resultid="102073" heatid="105258" lane="3" entrytime="00:01:09.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99425" points="599" reactiontime="+83" swimtime="00:00:31.63" resultid="102074" heatid="105362" lane="6" entrytime="00:00:31.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="DOL" clubid="102056" name="MUKP Just Swim Jelenia Góra">
          <CONTACT city="Jelenia Góra" email="marcin.binasiewicz@justswim.pl" name="Binasiewicz Marcin" phone="509071929" state="DOL" zip="58-506" />
          <ATHLETES>
            <ATHLETE birthdate="1986-05-26" firstname="Paweł" gender="M" lastname="Szkudlarek" nation="POL" athleteid="105104">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="105105" heatid="105143" lane="8" entrytime="00:00:25.00" />
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="105106" heatid="105275" lane="8" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-09-10" firstname="Mariusz" gender="M" lastname="Winogrodzki" nation="POL" license="50300120013" athleteid="105107">
              <RESULTS>
                <RESULT eventid="98798" points="574" reactiontime="+88" swimtime="00:00:25.15" resultid="105108" heatid="105143" lane="1" entrytime="00:00:25.00" />
                <RESULT comment="Rekord Polski Masters" eventid="99091" points="693" reactiontime="+82" swimtime="00:01:06.05" resultid="105109" heatid="105258" lane="5" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-05-01" firstname="Andrzej" gender="M" lastname="Waszkewicz" nation="POL" license="M0300120009" athleteid="105110">
              <RESULTS>
                <RESULT comment="04" eventid="98798" reactiontime="+80" status="DSQ" swimtime="00:00:00.00" resultid="105111" heatid="105143" lane="5" entrytime="00:00:23.82" />
                <RESULT eventid="99170" points="648" reactiontime="+95" swimtime="00:00:25.92" resultid="105112" heatid="105276" lane="5" entrytime="00:00:25.20" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="100913" name="Masters Bialystok">
          <CONTACT name="DOMINIKA MICHALIK" phone="608642788" />
          <ATHLETES>
            <ATHLETE birthdate="1965-01-01" firstname="Andrzej" gender="M" lastname="TWAROWSKI" nation="POL" athleteid="100914">
              <RESULTS>
                <RESULT eventid="98830" points="187" reactiontime="+91" swimtime="00:03:19.06" resultid="100915" heatid="105151" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.40" />
                    <SPLIT distance="100" swimtime="00:01:30.24" />
                    <SPLIT distance="150" swimtime="00:02:29.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="261" reactiontime="+111" swimtime="00:00:37.58" resultid="100916" heatid="105186" lane="9" entrytime="00:00:37.00" />
                <RESULT eventid="99020" points="126" reactiontime="+100" swimtime="00:03:42.24" resultid="100917" heatid="105233" lane="1" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.79" />
                    <SPLIT distance="100" swimtime="00:01:46.51" />
                    <SPLIT distance="150" swimtime="00:02:44.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="231" reactiontime="+70" swimtime="00:01:24.63" resultid="100918" heatid="105284" lane="0" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="177" reactiontime="+104" swimtime="00:07:14.05" resultid="100919" heatid="106049" lane="5" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.93" />
                    <SPLIT distance="100" swimtime="00:01:43.23" />
                    <SPLIT distance="150" swimtime="00:02:37.78" />
                    <SPLIT distance="200" swimtime="00:03:31.60" />
                    <SPLIT distance="250" swimtime="00:04:31.60" />
                    <SPLIT distance="300" swimtime="00:05:32.58" />
                    <SPLIT distance="350" swimtime="00:06:25.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="193" reactiontime="+80" swimtime="00:03:13.34" resultid="100920" heatid="105339" lane="9" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.93" />
                    <SPLIT distance="100" swimtime="00:01:31.39" />
                    <SPLIT distance="150" swimtime="00:02:23.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="248" reactiontime="+97" swimtime="00:00:42.41" resultid="100921" heatid="105356" lane="4" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-01" firstname="Dominika" gender="F" lastname="MICHALIK" nation="POL" swrid="4595750" athleteid="100922">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski Masters" eventid="98863" points="470" reactiontime="+103" swimtime="00:10:34.85" resultid="100923" heatid="105404" lane="3" entrytime="00:10:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.61" />
                    <SPLIT distance="100" swimtime="00:01:12.48" />
                    <SPLIT distance="150" swimtime="00:01:51.91" />
                    <SPLIT distance="200" swimtime="00:02:31.90" />
                    <SPLIT distance="250" swimtime="00:03:12.06" />
                    <SPLIT distance="300" swimtime="00:03:52.27" />
                    <SPLIT distance="350" swimtime="00:04:32.35" />
                    <SPLIT distance="400" swimtime="00:05:12.82" />
                    <SPLIT distance="450" swimtime="00:05:53.17" />
                    <SPLIT distance="500" swimtime="00:06:33.23" />
                    <SPLIT distance="550" swimtime="00:07:13.55" />
                    <SPLIT distance="600" swimtime="00:07:53.99" />
                    <SPLIT distance="650" swimtime="00:08:34.62" />
                    <SPLIT distance="700" swimtime="00:09:15.51" />
                    <SPLIT distance="750" swimtime="00:09:56.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="482" reactiontime="+85" swimtime="00:01:06.37" resultid="100924" heatid="105211" lane="3" entrytime="00:01:06.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99202" points="486" reactiontime="+77" swimtime="00:02:23.61" resultid="100925" heatid="105294" lane="1" entrytime="00:02:23.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                    <SPLIT distance="100" swimtime="00:01:08.06" />
                    <SPLIT distance="150" swimtime="00:01:45.69" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99457" points="474" reactiontime="+91" swimtime="00:05:06.55" resultid="100926" heatid="106054" lane="2" entrytime="00:05:04.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                    <SPLIT distance="100" swimtime="00:01:13.50" />
                    <SPLIT distance="150" swimtime="00:01:52.51" />
                    <SPLIT distance="200" swimtime="00:02:32.02" />
                    <SPLIT distance="250" swimtime="00:03:11.13" />
                    <SPLIT distance="300" swimtime="00:03:50.07" />
                    <SPLIT distance="350" swimtime="00:04:28.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Jaroslaw" gender="M" lastname="PAWLIK" nation="POL" swrid="4754662" athleteid="100927">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="100928" heatid="105127" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="100929" heatid="105215" lane="0" entrytime="00:01:25.00" />
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="100930" heatid="105267" lane="3" entrytime="00:00:39.00" />
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="100931" heatid="105326" lane="9" entrytime="00:01:50.00" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="100932" heatid="105352" lane="4" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Joanna" gender="F" lastname="WASILEWICZ" nation="POL" swrid="4876623" athleteid="100933">
              <RESULTS>
                <RESULT eventid="98777" points="247" reactiontime="+89" swimtime="00:00:37.80" resultid="100934" heatid="105115" lane="6" entrytime="00:00:38.17" entrycourse="LCM" />
                <RESULT eventid="98907" status="DNS" swimtime="00:00:00.00" resultid="100935" heatid="105172" lane="2" />
                <RESULT eventid="98972" points="204" swimtime="00:01:28.35" resultid="100936" heatid="105207" lane="0" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" status="DNS" swimtime="00:00:00.00" resultid="100937" heatid="105277" lane="4" entrytime="00:01:50.00" />
                <RESULT eventid="99202" points="188" reactiontime="+87" swimtime="00:03:17.00" resultid="100938" heatid="105290" lane="4" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.03" />
                    <SPLIT distance="100" swimtime="00:01:32.16" />
                    <SPLIT distance="150" swimtime="00:02:24.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" status="DNS" swimtime="00:00:00.00" resultid="100939" heatid="105344" lane="0" />
                <RESULT eventid="99457" points="181" reactiontime="+81" swimtime="00:07:02.16" resultid="100940" heatid="106056" lane="9" entrytime="00:06:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.46" />
                    <SPLIT distance="100" swimtime="00:01:32.10" />
                    <SPLIT distance="150" swimtime="00:02:26.53" />
                    <SPLIT distance="200" swimtime="00:03:22.23" />
                    <SPLIT distance="250" swimtime="00:04:18.42" />
                    <SPLIT distance="300" swimtime="00:05:15.67" />
                    <SPLIT distance="350" swimtime="00:06:11.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Miroslaw" gender="M" lastname="MATUSIK" nation="POL" swrid="4876624" athleteid="100941">
              <RESULTS>
                <RESULT eventid="98798" points="242" reactiontime="+97" swimtime="00:00:33.51" resultid="100942" heatid="105129" lane="7" entrytime="00:00:33.00" />
                <RESULT eventid="98891" points="199" swimtime="00:24:49.47" resultid="100943" heatid="105423" lane="2" entrytime="00:23:50.00" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="100944" heatid="105217" lane="6" entrytime="00:01:13.00" />
                <RESULT eventid="99020" status="DNS" swimtime="00:00:00.00" resultid="100945" heatid="105233" lane="3" entrytime="00:03:40.00" />
                <RESULT eventid="99170" points="257" reactiontime="+104" swimtime="00:00:35.24" resultid="100946" heatid="105270" lane="0" entrytime="00:00:35.00" />
                <RESULT eventid="99218" points="232" reactiontime="+104" swimtime="00:02:45.77" resultid="100947" heatid="105299" lane="0" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.24" />
                    <SPLIT distance="100" swimtime="00:01:18.87" />
                    <SPLIT distance="150" swimtime="00:02:02.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="100948" heatid="105326" lane="4" entrytime="00:01:30.00" />
                <RESULT eventid="99473" points="229" reactiontime="+113" swimtime="00:05:59.50" resultid="100949" heatid="106063" lane="0" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.96" />
                    <SPLIT distance="100" swimtime="00:01:23.35" />
                    <SPLIT distance="150" swimtime="00:02:09.26" />
                    <SPLIT distance="200" swimtime="00:02:55.49" />
                    <SPLIT distance="250" swimtime="00:03:41.86" />
                    <SPLIT distance="300" swimtime="00:04:29.30" />
                    <SPLIT distance="350" swimtime="00:05:16.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-01-01" firstname="Kazimiera" gender="F" lastname="RAINKO" nation="POL" athleteid="100950">
              <RESULTS>
                <RESULT eventid="98777" points="192" reactiontime="+102" swimtime="00:00:41.08" resultid="100951" heatid="105115" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="98907" points="91" reactiontime="+90" swimtime="00:01:00.14" resultid="100952" heatid="105173" lane="8" entrytime="00:00:55.00" />
                <RESULT eventid="98972" points="176" swimtime="00:01:32.80" resultid="100953" heatid="105206" lane="7" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="88" reactiontime="+132" swimtime="00:00:56.32" resultid="100954" heatid="105259" lane="1" entrytime="00:00:55.00" />
                <RESULT eventid="99202" points="140" reactiontime="+113" swimtime="00:03:37.20" resultid="100955" heatid="105289" lane="5" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.00" />
                    <SPLIT distance="100" swimtime="00:01:43.08" />
                    <SPLIT distance="150" swimtime="00:02:41.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="128" reactiontime="+103" swimtime="00:07:53.31" resultid="100956" heatid="106057" lane="5" entrytime="00:07:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.61" />
                    <SPLIT distance="100" swimtime="00:01:47.80" />
                    <SPLIT distance="150" swimtime="00:02:47.01" />
                    <SPLIT distance="200" swimtime="00:03:47.94" />
                    <SPLIT distance="250" swimtime="00:04:49.54" />
                    <SPLIT distance="300" swimtime="00:05:51.88" />
                    <SPLIT distance="350" swimtime="00:06:55.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-01" firstname="Maciej" gender="M" lastname="DASZUTA" nation="POL" athleteid="100957">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="100958" heatid="105138" lane="6" entrytime="00:00:28.00" />
                <RESULT eventid="98924" status="DNS" swimtime="00:00:00.00" resultid="100959" heatid="105188" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="100960" heatid="105256" lane="2" entrytime="00:01:20.00" />
                <RESULT eventid="99186" status="DNS" swimtime="00:00:00.00" resultid="100961" heatid="105285" lane="8" entrytime="00:01:18.00" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="100962" heatid="105361" lane="9" entrytime="00:00:34.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="100134" name="Masters Chełm">
          <CONTACT email="wepa56@interia.pl" name="Wiesław Wepa" />
          <ATHLETES>
            <ATHLETE birthdate="1941-10-11" firstname="Janusz" gender="M" lastname="GOLIK" nation="POL" swrid="4187077" athleteid="100135">
              <RESULTS>
                <RESULT eventid="98956" points="142" reactiontime="+114" swimtime="00:04:03.10" resultid="100136" heatid="105197" lane="8" entrytime="00:03:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.65" />
                    <SPLIT distance="100" swimtime="00:02:00.29" />
                    <SPLIT distance="150" swimtime="00:03:06.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="63" reactiontime="+119" swimtime="00:04:39.70" resultid="100137" heatid="105232" lane="2" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.14" />
                    <SPLIT distance="100" swimtime="00:02:13.19" />
                    <SPLIT distance="150" swimtime="00:03:26.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="161" reactiontime="+118" swimtime="00:01:47.25" resultid="100138" heatid="105250" lane="7" entrytime="00:01:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="92" reactiontime="+112" swimtime="00:00:49.58" resultid="100139" heatid="105265" lane="6" entrytime="00:00:58.00" />
                <RESULT eventid="99361" points="80" reactiontime="+125" swimtime="00:01:55.53" resultid="100140" heatid="105325" lane="5" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="190" reactiontime="+123" swimtime="00:00:46.38" resultid="100141" heatid="105353" lane="5" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="RUS" clubid="100118" name="Masters Club Sports Swimming YAMAL" shortname="Mrs CS Swimming YAMAL">
          <CONTACT email="www.swimmingyanao.ru" fax="3493633181" name="Lenchitskii Vladimir" phone="79224555665" street="glubokinsky 11 MKR. 94 house." />
          <ATHLETES>
            <ATHLETE birthdate="1962-10-07" firstname="Vladimir" gender="M" lastname="LENCHITSKII" nation="RUS" swrid="4595638" athleteid="100119">
              <RESULTS>
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="100120" heatid="105154" lane="9" entrytime="00:02:54.00" />
                <RESULT eventid="99020" status="DNS" swimtime="00:00:00.00" resultid="100121" heatid="105235" lane="7" entrytime="00:02:50.00" />
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="100122" heatid="105273" lane="9" entrytime="00:00:30.50" />
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="100123" heatid="105301" lane="0" entrytime="00:02:28.00" />
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="100124" heatid="105329" lane="0" entrytime="00:01:14.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="LBS" clubid="101883" name="Masters Gorzów">
          <CONTACT city="Kłodawa" email="mastersgorzow@onet.eu" name="Wojciechowicz Marek" phone="602891603" state="LUB" street="Skalna 2" zip="66-415" />
          <ATHLETES>
            <ATHLETE birthdate="1979-01-26" firstname="Stanisław" gender="M" lastname="KACZMAREK" nation="POL" athleteid="101918">
              <RESULTS>
                <RESULT eventid="98798" points="408" reactiontime="+79" swimtime="00:00:28.18" resultid="101919" heatid="105139" lane="6" entrytime="00:00:27.50" entrycourse="LCM" />
                <RESULT eventid="98830" points="431" reactiontime="+79" swimtime="00:02:30.81" resultid="101920" heatid="105157" lane="8" entrytime="00:02:31.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                    <SPLIT distance="100" swimtime="00:01:13.50" />
                    <SPLIT distance="150" swimtime="00:01:56.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="395" reactiontime="+80" swimtime="00:02:53.06" resultid="101921" heatid="105203" lane="9" entrytime="00:02:59.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                    <SPLIT distance="100" swimtime="00:01:23.00" />
                    <SPLIT distance="150" swimtime="00:02:09.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="361" reactiontime="+95" swimtime="00:02:36.58" resultid="101922" heatid="105236" lane="3" entrytime="00:02:28.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.86" />
                    <SPLIT distance="100" swimtime="00:01:14.39" />
                    <SPLIT distance="150" swimtime="00:01:55.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="415" reactiontime="+86" swimtime="00:02:16.66" resultid="101923" heatid="105299" lane="4" entrytime="00:02:35.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                    <SPLIT distance="100" swimtime="00:01:06.99" />
                    <SPLIT distance="150" swimtime="00:01:42.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="400" reactiontime="+88" swimtime="00:05:30.72" resultid="101924" heatid="106053" lane="7" entrytime="00:05:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                    <SPLIT distance="100" swimtime="00:01:10.42" />
                    <SPLIT distance="150" swimtime="00:01:57.49" />
                    <SPLIT distance="200" swimtime="00:02:42.86" />
                    <SPLIT distance="250" swimtime="00:03:30.25" />
                    <SPLIT distance="300" swimtime="00:04:17.48" />
                    <SPLIT distance="350" swimtime="00:04:55.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="372" reactiontime="+77" swimtime="00:01:09.23" resultid="101925" heatid="105331" lane="9" entrytime="00:01:04.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="423" reactiontime="+82" swimtime="00:04:53.06" resultid="101926" heatid="106059" lane="9" entrytime="00:04:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.98" />
                    <SPLIT distance="100" swimtime="00:01:10.39" />
                    <SPLIT distance="150" swimtime="00:01:47.35" />
                    <SPLIT distance="200" swimtime="00:02:24.93" />
                    <SPLIT distance="250" swimtime="00:03:02.64" />
                    <SPLIT distance="300" swimtime="00:03:40.08" />
                    <SPLIT distance="350" swimtime="00:04:17.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-05-08" firstname="Dawid" gender="M" lastname="BORUS" nation="POL" swrid="4992795" athleteid="101927">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="101928" heatid="105137" lane="0" entrytime="00:00:28.50" entrycourse="LCM" />
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="101929" heatid="105155" lane="5" entrytime="00:02:40.00" entrycourse="LCM" />
                <RESULT eventid="98924" status="DNS" swimtime="00:00:00.00" resultid="101930" heatid="105188" lane="3" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="101931" heatid="105254" lane="0" entrytime="00:01:25.00" entrycourse="LCM" />
                <RESULT eventid="99186" status="DNS" swimtime="00:00:00.00" resultid="101932" heatid="105286" lane="5" entrytime="00:01:11.50" entrycourse="LCM" />
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="101933" heatid="105341" lane="5" entrytime="00:02:38.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-02-20" firstname="Artur" gender="M" lastname="RUTKOWSKI" nation="POL" swrid="4992794" athleteid="101934">
              <RESULTS>
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="101935" heatid="105154" lane="6" entrytime="00:02:46.00" entrycourse="LCM" />
                <RESULT eventid="99020" status="DNS" swimtime="00:00:00.00" resultid="101936" heatid="105235" lane="8" entrytime="00:02:54.00" entrycourse="LCM" />
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="101937" heatid="105271" lane="5" entrytime="00:00:31.50" entrycourse="LCM" />
                <RESULT eventid="99282" status="DNS" swimtime="00:00:00.00" resultid="101938" heatid="106052" lane="9" entrytime="00:06:00.00" entrycourse="LCM" />
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="101939" heatid="105329" lane="7" entrytime="00:01:13.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-12-12" firstname="Marek" gender="M" lastname="WOJCIECHOWICZ" nation="POL" swrid="4967126" athleteid="101940">
              <RESULTS>
                <RESULT eventid="98798" status="WDR" swimtime="00:00:00.00" resultid="101941" heatid="105138" lane="4" entrytime="00:00:28.00" entrycourse="LCM" />
                <RESULT eventid="98891" status="WDR" swimtime="00:00:00.00" resultid="101942" entrytime="00:21:20.00" entrycourse="LCM" />
                <RESULT eventid="98988" status="WDR" swimtime="00:00:00.00" resultid="101943" heatid="105224" lane="1" entrytime="00:01:02.00" entrycourse="LCM" />
                <RESULT eventid="99170" status="WDR" swimtime="00:00:00.00" resultid="101944" heatid="105271" lane="7" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="99218" status="WDR" swimtime="00:00:00.00" resultid="101945" heatid="105302" lane="1" entrytime="00:02:20.00" entrycourse="LCM" />
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="101946" entrytime="00:05:10.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99059" status="DNS" swimtime="00:00:00.00" resultid="101947" heatid="105242" lane="8" entrytime="00:02:08.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101927" number="1" />
                    <RELAYPOSITION athleteid="101918" number="2" />
                    <RELAYPOSITION athleteid="101934" number="3" />
                    <RELAYPOSITION athleteid="101940" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" status="DNS" swimtime="00:00:00.00" resultid="101948" heatid="105311" lane="7" entrytime="00:01:52.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101934" number="1" />
                    <RELAYPOSITION athleteid="101927" number="2" />
                    <RELAYPOSITION athleteid="101940" number="3" />
                    <RELAYPOSITION athleteid="101918" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="KORONA KRA" nation="POL" region="MAL" clubid="103284" name="Masters Korona Kraków">
          <CONTACT city="Kraków" email="masterskorona@wp.pl" name="Mariola Kuliś" phone="500677133" state="MAŁ" street="Kalwaryjska" />
          <ATHLETES>
            <ATHLETE birthdate="1982-02-08" firstname="Tomasz" gender="M" lastname="CZERNIECKI" nation="POL" swrid="4992807" athleteid="103316">
              <RESULTS>
                <RESULT eventid="98798" points="507" reactiontime="+72" swimtime="00:00:26.22" resultid="103317" heatid="105142" lane="6" entrytime="00:00:26.00" />
                <RESULT eventid="98988" points="474" reactiontime="+77" swimtime="00:01:00.16" resultid="103318" heatid="105224" lane="8" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="396" reactiontime="+98" swimtime="00:00:30.54" resultid="103319" heatid="105272" lane="2" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-06-04" firstname="Andrzej" gender="M" lastname="DATA" nation="POL" swrid="4992806" athleteid="103320">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="103321" heatid="105128" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="98891" points="118" swimtime="00:29:31.00" resultid="103322" heatid="105425" lane="8" entrytime="00:24:00.00" />
                <RESULT eventid="98956" status="DNS" swimtime="00:00:00.00" resultid="103323" heatid="105199" lane="4" entrytime="00:03:27.00" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="103324" heatid="105216" lane="6" entrytime="00:01:16.00" />
                <RESULT eventid="99091" points="178" reactiontime="+134" swimtime="00:01:43.91" resultid="103325" heatid="105251" lane="3" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="136" reactiontime="+129" swimtime="00:03:17.91" resultid="103326" heatid="105297" lane="5" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.24" />
                    <SPLIT distance="100" swimtime="00:01:28.30" />
                    <SPLIT distance="150" swimtime="00:02:23.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="206" reactiontime="+116" swimtime="00:00:45.10" resultid="103327" heatid="105352" lane="5" entrytime="00:00:47.00" />
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="103328" entrytime="00:06:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-09-18" firstname="Izabela" gender="F" lastname="FRĄCZEK" nation="POL" swrid="4992822" athleteid="103329">
              <RESULTS>
                <RESULT eventid="98777" points="467" reactiontime="+80" swimtime="00:00:30.57" resultid="103330" heatid="105120" lane="2" entrytime="00:00:30.24" entrycourse="SCM" />
                <RESULT eventid="98907" points="345" reactiontime="+74" swimtime="00:00:38.57" resultid="103331" heatid="105177" lane="2" entrytime="00:00:37.50" />
                <RESULT eventid="98972" points="439" reactiontime="+87" swimtime="00:01:08.48" resultid="103332" heatid="105211" lane="2" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="390" reactiontime="+85" swimtime="00:00:34.31" resultid="103333" heatid="105262" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="99202" points="321" reactiontime="+85" swimtime="00:02:44.91" resultid="103334" heatid="105293" lane="8" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                    <SPLIT distance="100" swimtime="00:01:17.97" />
                    <SPLIT distance="150" swimtime="00:02:01.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="265" reactiontime="+86" swimtime="00:00:45.88" resultid="103335" heatid="105348" lane="8" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-08-18" firstname="Jadwiga" gender="F" lastname="GORECKA- BURKOT" nation="POL" swrid="4992800" athleteid="103336">
              <RESULTS>
                <RESULT eventid="98777" points="306" reactiontime="+79" swimtime="00:00:35.19" resultid="103337" heatid="105117" lane="2" entrytime="00:00:34.85" entrycourse="SCM" />
                <RESULT eventid="98972" points="254" reactiontime="+89" swimtime="00:01:22.20" resultid="103338" heatid="105207" lane="5" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="187" swimtime="00:00:43.78" resultid="103339" heatid="105260" lane="7" entrytime="00:00:43.00" />
                <RESULT eventid="99202" status="DNS" swimtime="00:00:00.00" resultid="103340" heatid="105289" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-12-23" firstname="Anna" gender="F" lastname="JANECZKO" nation="POL" swrid="4218717" athleteid="103341">
              <RESULTS>
                <RESULT eventid="98777" points="307" reactiontime="+104" swimtime="00:00:35.14" resultid="103342" heatid="105117" lane="5" entrytime="00:00:34.38" entrycourse="SCM" />
                <RESULT eventid="98814" points="199" reactiontime="+101" swimtime="00:03:36.07" resultid="103343" heatid="105144" lane="5" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.63" />
                    <SPLIT distance="100" swimtime="00:01:45.07" />
                    <SPLIT distance="150" swimtime="00:02:48.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" status="DNS" swimtime="00:00:00.00" resultid="103344" heatid="105175" lane="2" entrytime="00:00:41.98" />
                <RESULT eventid="99154" status="DNS" swimtime="00:00:00.00" resultid="103345" heatid="105261" lane="5" entrytime="00:00:37.68" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-07-27" firstname="Mariola" gender="F" lastname="KULIŚ" nation="POL" swrid="4992797" athleteid="103346">
              <RESULTS>
                <RESULT eventid="98777" points="411" reactiontime="+70" swimtime="00:00:31.91" resultid="103347" heatid="105120" lane="9" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="98907" points="394" reactiontime="+72" swimtime="00:00:36.91" resultid="103348" heatid="105173" lane="3" entrytime="00:00:50.00" />
                <RESULT eventid="98972" points="366" reactiontime="+74" swimtime="00:01:12.79" resultid="103349" heatid="105210" lane="8" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="349" reactiontime="+87" swimtime="00:01:31.38" resultid="103350" heatid="105243" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="381" reactiontime="+66" swimtime="00:00:34.58" resultid="103351" heatid="105263" lane="8" entrytime="00:00:34.50" />
                <RESULT eventid="99409" points="389" reactiontime="+79" swimtime="00:00:40.37" resultid="103352" heatid="105348" lane="4" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-09-12" firstname="Joanna" gender="F" lastname="KWATERA" nation="POL" swrid="4992811" athleteid="103353">
              <RESULTS>
                <RESULT eventid="98814" points="245" reactiontime="+67" swimtime="00:03:21.60" resultid="103354" heatid="105145" lane="8" entrytime="00:03:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.96" />
                    <SPLIT distance="100" swimtime="00:01:42.11" />
                    <SPLIT distance="150" swimtime="00:02:33.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="310" reactiontime="+86" swimtime="00:03:25.54" resultid="103355" heatid="105194" lane="9" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.36" />
                    <SPLIT distance="100" swimtime="00:01:38.03" />
                    <SPLIT distance="150" swimtime="00:02:32.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="269" reactiontime="+87" swimtime="00:01:39.63" resultid="103356" heatid="105246" lane="2" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" status="WDR" swimtime="00:00:00.00" resultid="103357" heatid="106045" lane="3" />
                <RESULT eventid="99409" points="295" reactiontime="+83" swimtime="00:00:44.26" resultid="103358" heatid="105347" lane="4" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-07-24" firstname="Bogusław" gender="M" lastname="KWIATKOWSKI" nation="POL" athleteid="103359">
              <RESULTS>
                <RESULT eventid="98798" points="35" reactiontime="+112" swimtime="00:01:03.61" resultid="103360" heatid="105123" lane="8" />
                <RESULT eventid="98924" points="26" reactiontime="+81" swimtime="00:01:20.58" resultid="103361" heatid="105180" lane="1" />
                <RESULT eventid="99091" points="31" reactiontime="+109" swimtime="00:03:05.46" resultid="103362" heatid="105248" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="20" reactiontime="+96" swimtime="00:03:10.79" resultid="103363" heatid="105281" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:30.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="44" reactiontime="+107" swimtime="00:01:15.42" resultid="103364" heatid="105350" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-16" firstname="Kamil" gender="M" lastname="LATUSZEK" nation="POL" swrid="4072741" athleteid="103365">
              <RESULTS>
                <RESULT eventid="98798" points="459" reactiontime="+82" swimtime="00:00:27.09" resultid="103366" heatid="105140" lane="3" entrytime="00:00:27.00" />
                <RESULT eventid="98988" points="491" reactiontime="+79" swimtime="00:00:59.44" resultid="103367" heatid="105225" lane="7" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="431" reactiontime="+83" swimtime="00:00:29.69" resultid="103368" heatid="105272" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="99218" points="370" reactiontime="+84" swimtime="00:02:22.03" resultid="103369" heatid="105302" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                    <SPLIT distance="100" swimtime="00:01:08.79" />
                    <SPLIT distance="150" swimtime="00:01:46.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="103370" entrytime="00:05:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-08-26" firstname="Andrzej" gender="M" lastname="MLECZKO" nation="POL" swrid="4992812" athleteid="103371">
              <RESULTS>
                <RESULT eventid="98798" points="220" reactiontime="+119" swimtime="00:00:34.62" resultid="103372" heatid="105127" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="98891" points="130" swimtime="00:28:37.04" resultid="103373" heatid="105424" lane="8" entrytime="00:28:08.00" />
                <RESULT eventid="98988" points="205" reactiontime="+122" swimtime="00:01:19.49" resultid="103374" heatid="105216" lane="3" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" status="DNS" swimtime="00:00:00.00" resultid="103375" heatid="105232" lane="6" entrytime="00:04:30.00" />
                <RESULT eventid="99218" points="164" reactiontime="+140" swimtime="00:03:06.10" resultid="103376" heatid="105297" lane="4" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.08" />
                    <SPLIT distance="100" swimtime="00:01:29.13" />
                    <SPLIT distance="150" swimtime="00:02:19.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="88" reactiontime="+143" swimtime="00:09:06.86" resultid="103377" heatid="106048" lane="1" entrytime="00:08:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.50" />
                    <SPLIT distance="100" swimtime="00:02:07.44" />
                    <SPLIT distance="150" swimtime="00:03:20.83" />
                    <SPLIT distance="200" swimtime="00:04:38.19" />
                    <SPLIT distance="250" swimtime="00:05:54.81" />
                    <SPLIT distance="300" swimtime="00:07:14.09" />
                    <SPLIT distance="350" swimtime="00:08:13.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="72" reactiontime="+119" swimtime="00:01:59.54" resultid="103378" heatid="105326" lane="8" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="146" reactiontime="+140" swimtime="00:06:57.29" resultid="103379" heatid="106065" lane="8" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.89" />
                    <SPLIT distance="100" swimtime="00:01:41.98" />
                    <SPLIT distance="150" swimtime="00:02:38.27" />
                    <SPLIT distance="200" swimtime="00:03:33.79" />
                    <SPLIT distance="250" swimtime="00:04:29.04" />
                    <SPLIT distance="300" swimtime="00:05:22.48" />
                    <SPLIT distance="350" swimtime="00:06:11.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-10-22" firstname="Maria" gender="F" lastname="MLECZKO" nation="POL" swrid="4992813" athleteid="103380">
              <RESULTS>
                <RESULT eventid="98777" points="48" reactiontime="+127" swimtime="00:01:05.04" resultid="103381" heatid="105113" lane="0" entrytime="00:00:59.29" entrycourse="SCM" />
                <RESULT eventid="98814" points="47" reactiontime="+120" swimtime="00:05:47.82" resultid="103382" heatid="105144" lane="9" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.59" />
                    <SPLIT distance="150" swimtime="00:04:35.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="67" reactiontime="+120" swimtime="00:05:42.02" resultid="103383" heatid="105191" lane="1" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.46" />
                    <SPLIT distance="100" swimtime="00:02:42.56" />
                    <SPLIT distance="150" swimtime="00:04:15.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="57" reactiontime="+106" swimtime="00:02:15.03" resultid="103384" heatid="105206" lane="9" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="34" reactiontime="+121" swimtime="00:01:16.95" resultid="103385" heatid="105259" lane="9" entrytime="00:01:17.00" />
                <RESULT eventid="99202" points="55" reactiontime="+117" swimtime="00:04:55.65" resultid="103386" heatid="105289" lane="7" entrytime="00:05:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.01" />
                    <SPLIT distance="100" swimtime="00:02:22.60" />
                    <SPLIT distance="150" swimtime="00:03:40.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="83" reactiontime="+124" swimtime="00:01:07.41" resultid="103387" heatid="105344" lane="2" entrytime="00:01:05.00" />
                <RESULT eventid="99457" points="51" reactiontime="+106" swimtime="00:10:44.56" resultid="103388" heatid="106057" lane="8" entrytime="00:10:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.49" />
                    <SPLIT distance="100" swimtime="00:02:19.52" />
                    <SPLIT distance="150" swimtime="00:03:37.70" />
                    <SPLIT distance="200" swimtime="00:04:57.92" />
                    <SPLIT distance="250" swimtime="00:06:17.14" />
                    <SPLIT distance="300" swimtime="00:07:40.09" />
                    <SPLIT distance="350" swimtime="00:09:15.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-08-01" firstname="Paulina" gender="F" lastname="PALMOWSKA" nation="POL" swrid="4992815" athleteid="103389">
              <RESULTS>
                <RESULT eventid="98814" points="434" reactiontime="+72" swimtime="00:02:46.60" resultid="103390" heatid="105146" lane="4" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.60" />
                    <SPLIT distance="100" swimtime="00:01:17.21" />
                    <SPLIT distance="150" swimtime="00:02:06.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="478" reactiontime="+75" swimtime="00:00:34.60" resultid="103391" heatid="105177" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="99314" points="464" reactiontime="+80" swimtime="00:01:15.05" resultid="103392" heatid="105280" lane="2" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.10" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99377" points="419" reactiontime="+78" swimtime="00:02:45.72" resultid="103393" heatid="105334" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.57" />
                    <SPLIT distance="100" swimtime="00:01:19.49" />
                    <SPLIT distance="150" swimtime="00:02:03.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="347" reactiontime="+86" swimtime="00:05:40.02" resultid="103394" heatid="106055" lane="5" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                    <SPLIT distance="100" swimtime="00:01:18.37" />
                    <SPLIT distance="150" swimtime="00:02:01.09" />
                    <SPLIT distance="200" swimtime="00:02:44.62" />
                    <SPLIT distance="250" swimtime="00:03:28.80" />
                    <SPLIT distance="300" swimtime="00:04:13.31" />
                    <SPLIT distance="350" swimtime="00:04:56.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-12-18" firstname="Szymon" gender="M" lastname="PYRĆ" nation="POL" swrid="4992817" athleteid="103395">
              <RESULTS>
                <RESULT eventid="98891" points="374" swimtime="00:20:07.93" resultid="103396" heatid="105421" lane="6" entrytime="00:20:35.00" />
                <RESULT eventid="99020" points="364" reactiontime="+77" swimtime="00:02:36.13" resultid="103397" heatid="105236" lane="9" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.48" />
                    <SPLIT distance="100" swimtime="00:01:13.55" />
                    <SPLIT distance="150" swimtime="00:01:54.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="337" reactiontime="+73" swimtime="00:00:32.21" resultid="103398" heatid="105272" lane="9" entrytime="00:00:31.30" />
                <RESULT eventid="99282" points="368" reactiontime="+67" swimtime="00:05:40.10" resultid="103399" heatid="106052" lane="8" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.52" />
                    <SPLIT distance="100" swimtime="00:01:12.03" />
                    <SPLIT distance="150" swimtime="00:01:59.28" />
                    <SPLIT distance="200" swimtime="00:02:44.79" />
                    <SPLIT distance="250" swimtime="00:03:34.40" />
                    <SPLIT distance="300" swimtime="00:04:23.87" />
                    <SPLIT distance="350" swimtime="00:05:03.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="375" reactiontime="+68" swimtime="00:01:09.03" resultid="103400" heatid="105330" lane="8" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-03-26" firstname="Józef" gender="M" lastname="ŚMIGIELSKI" nation="POL" athleteid="103401">
              <RESULTS>
                <RESULT eventid="98924" points="69" reactiontime="+109" swimtime="00:00:58.35" resultid="103402" heatid="105179" lane="4" />
                <RESULT eventid="99186" points="69" reactiontime="+131" swimtime="00:02:06.37" resultid="103403" heatid="105281" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="73" reactiontime="+112" swimtime="00:04:27.39" resultid="103404" heatid="105335" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.12" />
                    <SPLIT distance="100" swimtime="00:02:10.78" />
                    <SPLIT distance="150" swimtime="00:03:19.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="103405" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-07-04" firstname="Stanisław" gender="M" lastname="WAGA" nation="POL" swrid="4992823" athleteid="103406">
              <RESULTS>
                <RESULT eventid="98798" reactiontime="+82" status="DSQ" swimtime="00:00:00.00" resultid="103407" heatid="105124" lane="1" entrytime="00:00:45.00" />
                <RESULT eventid="98891" points="98" swimtime="00:31:23.00" resultid="103408" heatid="105425" lane="3" entrytime="00:30:30.00" />
                <RESULT eventid="98988" points="92" reactiontime="+119" swimtime="00:01:43.91" resultid="103409" heatid="105213" lane="3" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.36" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="07" eventid="99218" reactiontime="+127" status="DSQ" swimtime="00:00:00.00" resultid="103410" heatid="105295" lane="3" entrytime="00:03:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.02" />
                    <SPLIT distance="100" swimtime="00:01:50.67" />
                    <SPLIT distance="150" swimtime="00:02:51.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="85" reactiontime="+134" swimtime="00:08:18.81" resultid="103411" heatid="106066" lane="0" entrytime="00:07:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.85" />
                    <SPLIT distance="100" swimtime="00:02:02.38" />
                    <SPLIT distance="150" swimtime="00:03:06.84" />
                    <SPLIT distance="200" swimtime="00:04:11.06" />
                    <SPLIT distance="250" swimtime="00:05:14.31" />
                    <SPLIT distance="300" swimtime="00:06:16.87" />
                    <SPLIT distance="350" swimtime="00:07:19.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-26" firstname="Marta" gender="F" lastname="WYSOCKA" nation="POL" swrid="4992821" athleteid="103412">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski Masters" eventid="98940" points="346" reactiontime="+96" swimtime="00:03:18.14" resultid="103413" heatid="105193" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.07" />
                    <SPLIT distance="100" swimtime="00:01:35.61" />
                    <SPLIT distance="150" swimtime="00:02:26.99" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99089" points="340" reactiontime="+97" swimtime="00:01:32.11" resultid="103414" heatid="105246" lane="4" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.72" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99409" points="336" reactiontime="+89" swimtime="00:00:42.40" resultid="103415" heatid="105348" lane="7" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Masters Korona Kraków C" number="1">
              <RESULTS>
                <RESULT eventid="99250" points="366" reactiontime="+78" swimtime="00:01:58.52" resultid="103424" heatid="105310" lane="4" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.11" />
                    <SPLIT distance="100" swimtime="00:01:02.96" />
                    <SPLIT distance="150" swimtime="00:01:32.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103365" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="103320" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="103395" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="103316" number="4" reactiontime="+52" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Masters Korona Kraków C" number="1">
              <RESULTS>
                <RESULT eventid="99059" points="283" reactiontime="+100" swimtime="00:02:22.25" resultid="103425" heatid="105241" lane="0" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.95" />
                    <SPLIT distance="100" swimtime="00:01:24.00" />
                    <SPLIT distance="150" swimtime="00:01:56.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103371" number="1" reactiontime="+100" />
                    <RELAYPOSITION athleteid="103365" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="103395" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="103316" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="Masters Korona Kraków D" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="99036" points="360" reactiontime="+65" swimtime="00:02:29.07" resultid="103422" heatid="105238" lane="7" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.89" />
                    <SPLIT distance="100" swimtime="00:01:19.60" />
                    <SPLIT distance="150" swimtime="00:01:53.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103346" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="103412" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="103329" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="103336" number="4" reactiontime="+76" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99234" points="375" swimtime="00:02:14.18" resultid="103423" heatid="105307" lane="7" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                    <SPLIT distance="100" swimtime="00:01:07.41" />
                    <SPLIT distance="150" swimtime="00:01:38.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103336" number="1" />
                    <RELAYPOSITION athleteid="103329" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="103346" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="103412" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="Masters Korona Kraków B" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="286" reactiontime="+83" swimtime="00:02:08.69" resultid="103420" heatid="105160" lane="3" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                    <SPLIT distance="100" swimtime="00:01:07.54" />
                    <SPLIT distance="150" swimtime="00:01:42.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103389" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="103320" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="103341" number="3" reactiontime="+80" />
                    <RELAYPOSITION athleteid="103365" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" points="270" reactiontime="+76" swimtime="00:02:24.54" resultid="103421" heatid="105364" lane="3" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.14" />
                    <SPLIT distance="100" swimtime="00:01:19.32" />
                    <SPLIT distance="150" swimtime="00:01:48.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103389" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="103353" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="103365" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="103320" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Masters Korona Kraków C" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski Masters" eventid="98846" points="388" reactiontime="+83" swimtime="00:01:56.25" resultid="103418" heatid="105161" lane="1" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.20" />
                    <SPLIT distance="100" swimtime="00:01:00.54" />
                    <SPLIT distance="150" swimtime="00:01:30.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103346" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="103395" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="103329" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="103316" number="4" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" points="324" reactiontime="+81" swimtime="00:02:16.03" resultid="103419" heatid="105365" lane="1" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.99" />
                    <SPLIT distance="100" swimtime="00:01:18.75" />
                    <SPLIT distance="150" swimtime="00:01:50.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103329" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="103346" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="103395" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="103316" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" name="Masters Korona Kraków E" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="186" reactiontime="+94" swimtime="00:02:28.50" resultid="103416" heatid="105159" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                    <SPLIT distance="100" swimtime="00:01:19.37" />
                    <SPLIT distance="150" swimtime="00:01:54.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103336" number="1" reactiontime="+94" />
                    <RELAYPOSITION athleteid="103406" number="2" reactiontime="+7" />
                    <RELAYPOSITION athleteid="103412" number="3" reactiontime="+70" />
                    <RELAYPOSITION athleteid="103371" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" points="149" reactiontime="+70" swimtime="00:02:56.17" resultid="103417" heatid="105363" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.85" />
                    <SPLIT distance="100" swimtime="00:01:28.99" />
                    <SPLIT distance="150" swimtime="00:02:13.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103336" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="103412" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="103371" number="3" reactiontime="+64" />
                    <RELAYPOSITION athleteid="103406" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="LU" clubid="102019" name="Masters Kraśnik">
          <CONTACT city="Krasnik" email="jurek@krasnik.info" internet="www.masterskrasnik.za.pl" name="Michalczyk Jerzy" phone="601698977" state="LUB." street="Żwirki i Wigury 2" zip="23-210" />
          <ATHLETES>
            <ATHLETE birthdate="1953-09-27" firstname="Janusz" gender="M" lastname="WASIUK" nation="POL" swrid="4313185" athleteid="102020">
              <RESULTS>
                <RESULT eventid="98891" status="WDR" swimtime="00:00:00.00" resultid="102021" entrytime="00:33:13.21" />
                <RESULT eventid="98956" points="168" reactiontime="+127" swimtime="00:03:49.84" resultid="102022" heatid="105198" lane="0" entrytime="00:03:50.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.89" />
                    <SPLIT distance="100" swimtime="00:01:51.36" />
                    <SPLIT distance="150" swimtime="00:02:51.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="101" reactiontime="+129" swimtime="00:03:59.26" resultid="102023" heatid="105232" lane="0" entrytime="00:04:47.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.14" />
                    <SPLIT distance="100" swimtime="00:01:49.16" />
                    <SPLIT distance="150" swimtime="00:02:55.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="105" reactiontime="+137" swimtime="00:08:36.05" resultid="102024" heatid="106048" lane="8" entrytime="00:08:50.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.18" />
                    <SPLIT distance="100" swimtime="00:01:45.30" />
                    <SPLIT distance="150" swimtime="00:03:03.61" />
                    <SPLIT distance="200" swimtime="00:04:26.00" />
                    <SPLIT distance="250" swimtime="00:05:33.78" />
                    <SPLIT distance="300" swimtime="00:06:36.30" />
                    <SPLIT distance="350" swimtime="00:07:38.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="72" reactiontime="+110" swimtime="00:04:28.93" resultid="102025" heatid="105336" lane="2" entrytime="00:04:34.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.38" />
                    <SPLIT distance="100" swimtime="00:02:08.83" />
                    <SPLIT distance="150" swimtime="00:03:20.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-11-05" firstname="Krzysztof" gender="M" lastname="SAMONEK" nation="POL" swrid="4934017" athleteid="102026">
              <RESULTS>
                <RESULT eventid="98830" points="105" reactiontime="+107" swimtime="00:04:01.11" resultid="102027" heatid="105149" lane="3" entrytime="00:04:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.29" />
                    <SPLIT distance="100" swimtime="00:01:49.54" />
                    <SPLIT distance="150" swimtime="00:03:05.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="136" reactiontime="+74" swimtime="00:00:46.72" resultid="102028" heatid="105182" lane="1" entrytime="00:00:49.20" />
                <RESULT eventid="99020" points="62" reactiontime="+109" swimtime="00:04:40.64" resultid="102029" heatid="105232" lane="7" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.40" />
                    <SPLIT distance="100" swimtime="00:02:17.73" />
                    <SPLIT distance="150" swimtime="00:03:36.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="111" reactiontime="+84" swimtime="00:01:47.93" resultid="102030" heatid="105282" lane="6" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="94" reactiontime="+122" swimtime="00:08:54.55" resultid="102031" heatid="106048" lane="5" entrytime="00:08:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.65" />
                    <SPLIT distance="100" swimtime="00:02:09.82" />
                    <SPLIT distance="150" swimtime="00:03:19.16" />
                    <SPLIT distance="200" swimtime="00:04:23.64" />
                    <SPLIT distance="250" swimtime="00:05:42.76" />
                    <SPLIT distance="300" swimtime="00:06:58.38" />
                    <SPLIT distance="350" swimtime="00:07:58.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="102" reactiontime="+101" swimtime="00:03:58.81" resultid="105392" heatid="105337" lane="0" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.33" />
                    <SPLIT distance="100" swimtime="00:01:57.93" />
                    <SPLIT distance="150" swimtime="00:03:01.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-12-19" firstname="Waldemar" gender="M" lastname="RUSOWICZ" nation="POL" swrid="4934019" athleteid="102032">
              <RESULTS>
                <RESULT eventid="98830" points="105" reactiontime="+100" swimtime="00:04:01.60" resultid="102033" heatid="105149" lane="9" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.35" />
                    <SPLIT distance="100" swimtime="00:02:05.63" />
                    <SPLIT distance="150" swimtime="00:03:07.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="79" reactiontime="+91" swimtime="00:00:55.88" resultid="102034" heatid="105181" lane="7" entrytime="00:00:55.00" />
                <RESULT eventid="98956" points="168" reactiontime="+105" swimtime="00:03:49.93" resultid="102035" heatid="105197" lane="6" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.41" />
                    <SPLIT distance="100" swimtime="00:01:52.47" />
                    <SPLIT distance="150" swimtime="00:02:52.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="175" reactiontime="+96" swimtime="00:01:44.46" resultid="102036" heatid="105250" lane="8" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="121" reactiontime="+94" swimtime="00:01:44.97" resultid="102037" heatid="105282" lane="9" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="186" reactiontime="+110" swimtime="00:00:46.66" resultid="102038" heatid="105352" lane="2" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-03-04" firstname="Mirosław" gender="M" lastname="LESZCZYŃSKI" nation="POL" athleteid="102039">
              <RESULTS>
                <RESULT eventid="98956" points="299" reactiontime="+105" swimtime="00:03:09.93" resultid="102040" heatid="105200" lane="1" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.62" />
                    <SPLIT distance="100" swimtime="00:01:30.77" />
                    <SPLIT distance="150" swimtime="00:02:19.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="303" reactiontime="+99" swimtime="00:01:26.97" resultid="102041" heatid="105254" lane="8" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="102042" heatid="105336" lane="0" entrytime="00:05:00.00" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="102043" heatid="105356" lane="5" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-09" firstname="Jerzy" gender="M" lastname="MICHALCZYK" nation="POL" swrid="4934020" athleteid="102044">
              <RESULTS>
                <RESULT eventid="98830" points="105" reactiontime="+99" swimtime="00:04:01.36" resultid="102045" heatid="105149" lane="2" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.23" />
                    <SPLIT distance="100" swimtime="00:01:57.92" />
                    <SPLIT distance="150" swimtime="00:03:03.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="130" swimtime="00:04:10.20" resultid="102046" heatid="105197" lane="7" entrytime="00:03:55.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.21" />
                    <SPLIT distance="100" swimtime="00:02:00.03" />
                    <SPLIT distance="150" swimtime="00:03:08.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="142" reactiontime="+97" swimtime="00:01:51.96" resultid="102047" heatid="105249" lane="3" entrytime="00:01:55.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="108" reactiontime="+92" swimtime="00:00:46.99" resultid="102048" heatid="105265" lane="5" entrytime="00:00:55.00" />
                <RESULT eventid="99361" points="74" reactiontime="+98" swimtime="00:01:58.46" resultid="102049" heatid="105325" lane="3" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="152" reactiontime="+100" swimtime="00:00:49.97" resultid="102050" heatid="105352" lane="0" entrytime="00:00:48.35" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="101505" name="Masters MKP Szczecin">
          <CONTACT city="WOŁCZKOWO" email="mk@mastersswim.pl" internet="www.mastersswim.pl" name="KACZANOWSKI MIŁOSZ" phone="888181234" state="ZACHO" street="SŁONECZNA 5" zip="72-003" />
          <ATHLETES>
            <ATHLETE birthdate="1968-05-22" firstname="Miłosz" gender="M" lastname="KACZANOWSKI" nation="POL" swrid="4967269" athleteid="104998">
              <RESULTS>
                <RESULT eventid="98798" points="465" reactiontime="+72" swimtime="00:00:26.99" resultid="104999" heatid="105123" lane="7" />
                <RESULT eventid="98830" points="434" reactiontime="+68" swimtime="00:02:30.47" resultid="105000" heatid="105158" lane="9" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.80" />
                    <SPLIT distance="100" swimtime="00:01:09.75" />
                    <SPLIT distance="150" swimtime="00:01:53.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="413" swimtime="00:02:50.53" resultid="105001" heatid="105196" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                    <SPLIT distance="100" swimtime="00:01:20.45" />
                    <SPLIT distance="150" swimtime="00:02:05.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="473" reactiontime="+76" swimtime="00:01:00.18" resultid="105002" heatid="105226" lane="6" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="495" reactiontime="+82" swimtime="00:00:28.35" resultid="105003" heatid="105265" lane="1" />
                <RESULT eventid="99218" points="435" reactiontime="+83" swimtime="00:02:14.58" resultid="105004" heatid="105303" lane="5" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                    <SPLIT distance="100" swimtime="00:01:05.06" />
                    <SPLIT distance="150" swimtime="00:01:40.77" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99361" points="481" reactiontime="+78" swimtime="00:01:03.56" resultid="105005" heatid="105324" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="440" reactiontime="+79" swimtime="00:00:35.06" resultid="105006" heatid="105361" lane="1" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-09-25" firstname="Sławomir" gender="M" lastname="GRZESZEWSKI" nation="POL" athleteid="105007">
              <RESULTS>
                <RESULT eventid="98830" points="179" reactiontime="+97" swimtime="00:03:22.27" resultid="105008" heatid="105151" lane="0" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                    <SPLIT distance="100" swimtime="00:01:35.88" />
                    <SPLIT distance="150" swimtime="00:02:32.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="209" reactiontime="+93" swimtime="00:03:33.93" resultid="105009" heatid="105198" lane="4" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.29" />
                    <SPLIT distance="100" swimtime="00:01:42.99" />
                    <SPLIT distance="150" swimtime="00:02:38.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="233" reactiontime="+90" swimtime="00:01:34.94" resultid="105010" heatid="105251" lane="4" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="262" reactiontime="+91" swimtime="00:00:41.63" resultid="105011" heatid="105350" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-08-10" firstname="Małgorzata" gender="F" lastname="SERBIN" nation="POL" athleteid="105012">
              <RESULTS>
                <RESULT eventid="98777" points="399" reactiontime="+81" swimtime="00:00:32.21" resultid="105013" heatid="105120" lane="0" entrytime="00:00:30.69" />
                <RESULT eventid="98863" points="427" reactiontime="+77" swimtime="00:10:55.71" resultid="105014" heatid="105404" lane="7" entrytime="00:10:45.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                    <SPLIT distance="100" swimtime="00:01:14.49" />
                    <SPLIT distance="150" swimtime="00:01:55.04" />
                    <SPLIT distance="200" swimtime="00:02:35.65" />
                    <SPLIT distance="250" swimtime="00:03:16.81" />
                    <SPLIT distance="300" swimtime="00:03:58.45" />
                    <SPLIT distance="350" swimtime="00:04:39.98" />
                    <SPLIT distance="400" swimtime="00:05:21.51" />
                    <SPLIT distance="450" swimtime="00:06:03.40" />
                    <SPLIT distance="500" swimtime="00:06:45.07" />
                    <SPLIT distance="550" swimtime="00:07:27.20" />
                    <SPLIT distance="600" swimtime="00:08:09.05" />
                    <SPLIT distance="650" swimtime="00:08:51.19" />
                    <SPLIT distance="700" swimtime="00:09:33.11" />
                    <SPLIT distance="750" swimtime="00:10:15.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="405" swimtime="00:01:10.33" resultid="105015" heatid="105211" lane="7" entrytime="00:01:08.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="402" reactiontime="+73" swimtime="00:02:33.03" resultid="105016" heatid="105294" lane="7" entrytime="00:02:23.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                    <SPLIT distance="100" swimtime="00:01:13.79" />
                    <SPLIT distance="150" swimtime="00:01:53.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="357" reactiontime="+79" swimtime="00:02:54.79" resultid="105017" heatid="105334" lane="5" entrytime="00:02:49.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.98" />
                    <SPLIT distance="100" swimtime="00:01:26.59" />
                    <SPLIT distance="150" swimtime="00:02:11.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="378" reactiontime="+79" swimtime="00:05:30.50" resultid="105018" heatid="106054" lane="7" entrytime="00:05:07.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                    <SPLIT distance="100" swimtime="00:01:15.84" />
                    <SPLIT distance="150" swimtime="00:01:57.35" />
                    <SPLIT distance="200" swimtime="00:02:39.81" />
                    <SPLIT distance="250" swimtime="00:03:22.61" />
                    <SPLIT distance="300" swimtime="00:04:05.94" />
                    <SPLIT distance="350" swimtime="00:04:49.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-10-02" firstname="Jadwiga" gender="F" lastname="WEBER" nation="POL" athleteid="105019">
              <RESULTS>
                <RESULT eventid="98777" points="266" reactiontime="+92" swimtime="00:00:36.88" resultid="105020" heatid="105115" lane="0" entrytime="00:00:40.00" />
                <RESULT eventid="98907" points="272" reactiontime="+93" swimtime="00:00:41.72" resultid="105021" heatid="105174" lane="4" entrytime="00:00:43.00" />
                <RESULT eventid="98972" points="245" swimtime="00:01:23.13" resultid="105022" heatid="105207" lane="7" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.56" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99314" points="275" reactiontime="+91" swimtime="00:01:29.35" resultid="105023" heatid="105278" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.01" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99377" points="271" reactiontime="+90" swimtime="00:03:11.49" resultid="105024" heatid="105333" lane="7" entrytime="00:03:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.06" />
                    <SPLIT distance="100" swimtime="00:01:32.23" />
                    <SPLIT distance="150" swimtime="00:02:22.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1935-08-21" firstname="Stefania" gender="F" lastname="NOETZEL" nation="POL" athleteid="105025">
              <RESULTS>
                <RESULT eventid="98940" points="101" swimtime="00:04:58.32" resultid="105026" heatid="105191" lane="7" entrytime="00:04:55.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.01" />
                    <SPLIT distance="100" swimtime="00:02:26.80" />
                    <SPLIT distance="150" swimtime="00:03:43.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="93" swimtime="00:02:21.65" resultid="105027" heatid="105244" lane="8" entrytime="00:02:16.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="74" swimtime="00:01:10.07" resultid="105028" heatid="105344" lane="7" entrytime="00:01:05.72" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-11-14" firstname="Anna" gender="F" lastname="FRANKOWSKA" nation="POL" athleteid="105029">
              <RESULTS>
                <RESULT eventid="98777" points="248" reactiontime="+103" swimtime="00:00:37.77" resultid="105030" heatid="105115" lane="9" entrytime="00:00:40.00" />
                <RESULT eventid="98907" points="245" swimtime="00:00:43.21" resultid="105031" heatid="105173" lane="6" entrytime="00:00:50.00" />
                <RESULT eventid="99409" points="269" reactiontime="+101" swimtime="00:00:45.66" resultid="105032" heatid="105345" lane="4" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-02" firstname="Piotr" gender="M" lastname="KOWALCZYK" nation="POL" swrid="4992788" athleteid="105033">
              <RESULTS>
                <RESULT eventid="98891" points="374" swimtime="00:20:08.63" resultid="105034" heatid="105421" lane="4" entrytime="00:20:05.34" entrycourse="LCM" />
                <RESULT eventid="98988" points="416" reactiontime="+78" swimtime="00:01:02.82" resultid="105035" heatid="105223" lane="3" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="388" reactiontime="+84" swimtime="00:02:19.83" resultid="105036" heatid="105302" lane="4" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                    <SPLIT distance="100" swimtime="00:01:07.27" />
                    <SPLIT distance="150" swimtime="00:01:44.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="105037" heatid="105340" lane="6" entrytime="00:02:50.00" />
                <RESULT comment="04" eventid="99473" reactiontime="+83" status="DSQ" swimtime="00:00:00.00" resultid="105038" heatid="106061" lane="4" entrytime="00:04:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                    <SPLIT distance="100" swimtime="00:01:11.17" />
                    <SPLIT distance="150" swimtime="00:01:49.60" />
                    <SPLIT distance="200" swimtime="00:02:27.49" />
                    <SPLIT distance="250" swimtime="00:03:05.66" />
                    <SPLIT distance="300" swimtime="00:03:44.37" />
                    <SPLIT distance="350" swimtime="00:04:22.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT comment="Z 4 z 2/3 zmianę" eventid="98846" reactiontime="+89" status="DSQ" swimtime="00:02:18.31" resultid="105039" heatid="105160" lane="0" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.40" />
                    <SPLIT distance="100" swimtime="00:01:09.32" />
                    <SPLIT distance="150" swimtime="00:01:42.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="104998" number="1" reactiontime="+89" status="DSQ" />
                    <RELAYPOSITION athleteid="105019" number="2" reactiontime="+53" status="DSQ" />
                    <RELAYPOSITION athleteid="105029" number="3" reactiontime="-196" status="DSQ" />
                    <RELAYPOSITION athleteid="105007" number="4" reactiontime="+49" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="99441" points="156" reactiontime="+89" swimtime="00:02:53.31" resultid="105040" heatid="105363" lane="4" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:17.54" />
                    <SPLIT distance="100" swimtime="00:01:52.27" />
                    <SPLIT distance="150" swimtime="00:02:18.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="105019" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="105025" number="2" />
                    <RELAYPOSITION athleteid="104998" number="3" />
                    <RELAYPOSITION athleteid="105007" number="4" reactiontime="+69" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="UKR" clubid="101262" name="Masters Swimming Club EURO-LVIV" shortname="Mrs Swim. Club EURO-LV">
          <CONTACT city="Lviv" email="riff@mail.lviv.ua" fax="+380322430304" name="Ruslan Friauf" phone="+380676734796" street="Karpincya, 18A/3" zip="79012" />
          <ATHLETES>
            <ATHLETE birthdate="1976-02-23" firstname="Oleksandr" gender="M" lastname="SHAVROV" nation="UKR" swrid="4776479" athleteid="101263">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="101264" heatid="105135" lane="6" entrytime="00:00:29.40" />
                <RESULT eventid="98956" points="369" reactiontime="+92" swimtime="00:02:56.92" resultid="101265" heatid="105202" lane="3" entrytime="00:03:00.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.27" />
                    <SPLIT distance="100" swimtime="00:01:24.90" />
                    <SPLIT distance="150" swimtime="00:02:10.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="417" reactiontime="+77" swimtime="00:01:18.23" resultid="101266" heatid="105256" lane="8" entrytime="00:01:20.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="470" reactiontime="+76" swimtime="00:00:34.30" resultid="101267" heatid="105359" lane="4" entrytime="00:00:35.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-06-24" firstname="Inna" gender="F" lastname="HORDII" nation="UKR" swrid="4967000" athleteid="101268">
              <RESULTS>
                <RESULT eventid="98777" points="415" reactiontime="+89" swimtime="00:00:31.81" resultid="101269" heatid="105118" lane="4" entrytime="00:00:32.45" entrycourse="LCM" />
                <RESULT eventid="98907" points="312" reactiontime="+80" swimtime="00:00:39.88" resultid="101270" heatid="105176" lane="1" entrytime="00:00:39.20" />
                <RESULT eventid="98972" points="364" reactiontime="+87" swimtime="00:01:12.87" resultid="101271" heatid="105211" lane="8" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="325" reactiontime="+89" swimtime="00:00:36.46" resultid="101272" heatid="105262" lane="8" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-06-05" firstname="Mykhailo" gender="M" lastname="SHELEST" nation="UKR" swrid="4776480" athleteid="101273">
              <RESULTS>
                <RESULT eventid="98924" points="222" reactiontime="+80" swimtime="00:00:39.68" resultid="101274" heatid="105185" lane="4" entrytime="00:00:37.50" />
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="101275" heatid="105253" lane="3" entrytime="00:01:27.00" />
                <RESULT eventid="99425" points="300" reactiontime="+107" swimtime="00:00:39.83" resultid="101276" heatid="105358" lane="1" entrytime="00:00:37.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-07-31" firstname="Roman" gender="M" lastname="KORETSKYY" nation="UKR" swrid="4743142" athleteid="101277">
              <RESULTS>
                <RESULT eventid="98798" points="162" reactiontime="+118" swimtime="00:00:38.31" resultid="101278" heatid="105127" lane="0" entrytime="00:00:36.00" />
                <RESULT eventid="98924" points="123" reactiontime="+98" swimtime="00:00:48.29" resultid="101279" heatid="105183" lane="2" entrytime="00:00:43.00" />
                <RESULT eventid="98988" points="145" reactiontime="+108" swimtime="00:01:29.10" resultid="101280" heatid="105215" lane="8" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="101" reactiontime="+82" swimtime="00:01:51.50" resultid="101281" heatid="105282" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-05-09" firstname="Lidiya" gender="F" lastname="TYMOSHENKO" nation="UKR" swrid="4776490" athleteid="101282">
              <RESULTS>
                <RESULT eventid="98777" points="127" reactiontime="+129" swimtime="00:00:47.19" resultid="101283" heatid="105113" lane="3" entrytime="00:00:45.59" entrycourse="LCM" />
                <RESULT eventid="98907" points="72" reactiontime="+102" swimtime="00:01:04.83" resultid="101284" heatid="105173" lane="0" entrytime="00:00:55.66" />
                <RESULT eventid="99089" points="122" reactiontime="+115" swimtime="00:02:09.67" resultid="101285" heatid="105244" lane="1" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="118" reactiontime="+140" swimtime="00:01:00.09" resultid="101286" heatid="105345" lane="0" entrytime="00:00:53.15" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-03-31" firstname="Myron" gender="M" lastname="KOLODKO" nation="UKR" swrid="5023956" athleteid="101287">
              <RESULTS>
                <RESULT eventid="98830" points="139" reactiontime="+114" swimtime="00:03:39.83" resultid="101288" heatid="105151" lane="8" entrytime="00:03:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.14" />
                    <SPLIT distance="100" swimtime="00:01:40.15" />
                    <SPLIT distance="150" swimtime="00:02:47.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="77" reactiontime="+122" swimtime="00:04:21.76" resultid="101289" heatid="105233" lane="2" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.83" />
                    <SPLIT distance="100" swimtime="00:01:54.22" />
                    <SPLIT distance="150" swimtime="00:03:07.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="101290" heatid="105267" lane="9" entrytime="00:00:41.00" />
                <RESULT eventid="99282" points="119" reactiontime="+144" swimtime="00:08:15.43" resultid="101291" heatid="106049" lane="0" entrytime="00:07:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.98" />
                    <SPLIT distance="100" swimtime="00:02:01.89" />
                    <SPLIT distance="150" swimtime="00:03:05.42" />
                    <SPLIT distance="200" swimtime="00:04:07.10" />
                    <SPLIT distance="250" swimtime="00:05:17.04" />
                    <SPLIT distance="300" swimtime="00:06:26.87" />
                    <SPLIT distance="350" swimtime="00:07:21.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="86" reactiontime="+136" swimtime="00:01:52.48" resultid="101292" heatid="105326" lane="6" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-02-05" firstname="Lyudmyla" gender="F" lastname="KHIRESH" nation="UKR" swrid="4743144" athleteid="101293">
              <RESULTS>
                <RESULT eventid="98907" points="288" reactiontime="+79" swimtime="00:00:40.96" resultid="101294" heatid="105177" lane="9" entrytime="00:00:39.00" />
                <RESULT eventid="99314" status="DNS" swimtime="00:00:00.00" resultid="101295" heatid="105279" lane="2" entrytime="00:01:27.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-06-23" firstname="Nadiya" gender="F" lastname="SANNIKOVA" nation="UKR" swrid="4743147" athleteid="101296">
              <RESULTS>
                <RESULT eventid="99089" status="DNS" swimtime="00:00:00.00" resultid="101297" heatid="105245" lane="9" entrytime="00:01:52.00" />
                <RESULT eventid="99409" status="DNS" swimtime="00:00:00.00" resultid="101298" heatid="105346" lane="7" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-31" firstname="Dmytro" gender="M" lastname="ANTIPOV" nation="UKR" swrid="4967001" athleteid="101299">
              <RESULTS>
                <RESULT eventid="98798" points="305" reactiontime="+92" swimtime="00:00:31.03" resultid="101300" heatid="105138" lane="8" entrytime="00:00:28.00" />
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="101301" heatid="105257" lane="9" entrytime="00:01:18.00" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="101302" heatid="105359" lane="6" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-02-03" firstname="Romana" gender="F" lastname="SIRENKO" nation="UKR" swrid="4743148" athleteid="101303">
              <RESULTS>
                <RESULT eventid="98814" status="DNS" swimtime="00:00:00.00" resultid="101304" heatid="105146" lane="1" entrytime="00:03:05.00" />
                <RESULT eventid="98907" status="DNS" swimtime="00:00:00.00" resultid="101305" heatid="105177" lane="0" entrytime="00:00:38.00" />
                <RESULT eventid="99154" status="DNS" swimtime="00:00:00.00" resultid="101306" heatid="105262" lane="3" entrytime="00:00:35.50" />
                <RESULT eventid="99344" status="DNS" swimtime="00:00:00.00" resultid="101307" heatid="105322" lane="5" entrytime="00:01:27.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-05-11" firstname="Nataliya" gender="F" lastname="HERTSYK" nation="UKR" swrid="4743141" athleteid="101308">
              <RESULTS>
                <RESULT eventid="98777" status="DNS" swimtime="00:00:00.00" resultid="101309" heatid="105114" lane="3" entrytime="00:00:40.39" entrycourse="LCM" />
                <RESULT eventid="99154" status="DNS" swimtime="00:00:00.00" resultid="101310" heatid="105260" lane="6" entrytime="00:00:40.87" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-01-07" firstname="Ruslan" gender="M" lastname="FRIAUF" nation="UKR" swrid="4776473" athleteid="101311">
              <RESULTS>
                <RESULT eventid="98830" points="232" reactiontime="+73" swimtime="00:03:05.36" resultid="101312" heatid="105154" lane="8" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                    <SPLIT distance="100" swimtime="00:01:25.55" />
                    <SPLIT distance="150" swimtime="00:02:19.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="249" reactiontime="+81" swimtime="00:00:38.21" resultid="101313" heatid="105186" lane="0" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-03-11" firstname="Taras" gender="M" lastname="KUNETS" nation="UKR" swrid="4966999" athleteid="101314">
              <RESULTS>
                <RESULT eventid="98798" points="386" reactiontime="+75" swimtime="00:00:28.71" resultid="101315" heatid="105139" lane="8" entrytime="00:00:27.50" />
                <RESULT eventid="98891" points="226" swimtime="00:23:49.36" resultid="101316" heatid="105420" lane="0" entrytime="00:19:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-11" firstname="Anatoliy" gender="M" lastname="PETRINKO" nation="UKR" swrid="4967004" athleteid="101317">
              <RESULTS>
                <RESULT eventid="98798" points="258" reactiontime="+104" swimtime="00:00:32.83" resultid="101318" heatid="105138" lane="5" entrytime="00:00:28.00" />
                <RESULT eventid="98988" points="202" reactiontime="+111" swimtime="00:01:19.90" resultid="101319" heatid="105218" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="101320" heatid="105273" lane="5" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-10-27" firstname="Yuriy" gender="M" lastname="DENISOV" nation="UKR" swrid="4595558" athleteid="101321">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="101322" heatid="105129" lane="1" entrytime="00:00:33.00" />
                <RESULT eventid="98988" points="319" reactiontime="+90" swimtime="00:01:08.63" resultid="101323" heatid="105215" lane="5" entrytime="00:01:20.00" />
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="101324" heatid="105252" lane="3" entrytime="00:01:30.00" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="101325" heatid="105353" lane="3" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-03-11" firstname="Lyudmyla" gender="F" lastname="MAKSYMIV" nation="UKR" swrid="4876576" athleteid="101326">
              <RESULTS>
                <RESULT eventid="98940" status="DNS" swimtime="00:00:00.00" resultid="101327" heatid="105193" lane="0" entrytime="00:03:42.00" />
                <RESULT eventid="99089" status="DNS" swimtime="00:00:00.00" resultid="101328" heatid="105245" lane="2" entrytime="00:01:45.00" />
                <RESULT eventid="99314" status="DNS" swimtime="00:00:00.00" resultid="101329" heatid="105278" lane="7" entrytime="00:01:40.00" />
                <RESULT eventid="99377" status="DNS" swimtime="00:00:00.00" resultid="101330" heatid="105332" lane="5" entrytime="00:03:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-11-13" firstname="Ihor" gender="M" lastname="YASKEVYCH" nation="UKR" swrid="4595559" athleteid="101331">
              <RESULTS>
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="101332" heatid="105253" lane="6" entrytime="00:01:27.00" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="101333" heatid="105357" lane="2" entrytime="00:00:38.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-05-31" firstname="Zenoviy" gender="M" lastname="KUSHNIR" nation="UKR" swrid="4743143" athleteid="101334">
              <RESULTS>
                <RESULT eventid="98924" points="72" reactiontime="+91" swimtime="00:00:57.53" resultid="101335" heatid="105181" lane="6" entrytime="00:00:54.00" />
                <RESULT eventid="99186" points="68" reactiontime="+85" swimtime="00:02:06.79" resultid="101336" heatid="105281" lane="4" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="68" reactiontime="+85" swimtime="00:04:33.96" resultid="101337" heatid="105336" lane="4" entrytime="00:04:15.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.42" />
                    <SPLIT distance="100" swimtime="00:02:16.58" />
                    <SPLIT distance="150" swimtime="00:03:29.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-06-27" firstname="Iurii" gender="M" lastname="MARTYNIUK" nation="UKR" swrid="4743145" athleteid="101338">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="101339" heatid="105135" lane="9" entrytime="00:00:29.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-02-18" firstname="Vladyslav" gender="M" lastname="HOROVOY" nation="UKR" swrid="4967005" athleteid="101340">
              <RESULTS>
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="101341" heatid="105226" lane="5" entrytime="00:00:58.50" />
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="101342" heatid="105304" lane="5" entrytime="00:02:11.00" />
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="101343" entrytime="00:04:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-06-28" firstname="Valentyna" gender="F" lastname="KVITA" nation="UKR" athleteid="101344">
              <RESULTS>
                <RESULT eventid="98777" status="DNS" swimtime="00:00:00.00" resultid="101345" heatid="105121" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="98863" status="WDR" swimtime="00:00:00.00" resultid="101346" entrytime="00:10:00.00" />
                <RESULT eventid="98972" status="DNS" swimtime="00:00:00.00" resultid="101347" heatid="105212" lane="0" entrytime="00:01:04.00" />
                <RESULT eventid="99202" status="DNS" swimtime="00:00:00.00" resultid="101348" heatid="105294" lane="2" entrytime="00:02:20.00" />
                <RESULT eventid="99457" status="DNS" swimtime="00:00:00.00" resultid="101349" heatid="106054" lane="6" entrytime="00:05:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-07-18" firstname="Igor" gender="M" lastname="SHCHOTKIN" nation="UKR" swrid="4301793" athleteid="101350">
              <RESULTS>
                <RESULT eventid="98798" points="547" reactiontime="+81" swimtime="00:00:25.56" resultid="101351" heatid="105142" lane="4" entrytime="00:00:25.10" />
                <RESULT eventid="98988" points="524" reactiontime="+80" swimtime="00:00:58.15" resultid="101352" heatid="105227" lane="5" entrytime="00:00:57.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="511" reactiontime="+77" swimtime="00:00:28.05" resultid="101353" heatid="105275" lane="6" entrytime="00:00:27.60" />
                <RESULT eventid="99425" points="529" reactiontime="+78" swimtime="00:00:32.97" resultid="101354" heatid="105361" lane="4" entrytime="00:00:32.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-08-05" firstname="Iryna" gender="F" lastname="PONOMARENKO" nation="UKR" swrid="4301791" athleteid="101355">
              <RESULTS>
                <RESULT eventid="98777" points="396" reactiontime="+110" swimtime="00:00:32.30" resultid="101356" heatid="105118" lane="1" entrytime="00:00:33.47" entrycourse="LCM" />
                <RESULT eventid="98972" points="400" reactiontime="+83" swimtime="00:01:10.65" resultid="101357" heatid="105211" lane="9" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="382" reactiontime="+92" swimtime="00:02:35.65" resultid="101358" heatid="105292" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                    <SPLIT distance="100" swimtime="00:01:14.92" />
                    <SPLIT distance="150" swimtime="00:01:55.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="319" reactiontime="+90" swimtime="00:00:43.11" resultid="101359" heatid="105348" lane="1" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="8">
              <RESULTS>
                <RESULT eventid="99059" points="239" reactiontime="+89" swimtime="00:02:30.54" resultid="101367" heatid="105242" lane="1" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                    <SPLIT distance="100" swimtime="00:01:13.83" />
                    <SPLIT distance="150" swimtime="00:01:57.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101340" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="101263" number="2" reactiontime="+33" />
                    <RELAYPOSITION athleteid="101317" number="3" reactiontime="+91" />
                    <RELAYPOSITION athleteid="101338" number="4" reactiontime="+63" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="9">
              <RESULTS>
                <RESULT eventid="99250" status="DNS" swimtime="00:00:00.00" resultid="101368" heatid="105311" lane="1" entrytime="00:01:54.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101338" number="1" />
                    <RELAYPOSITION athleteid="101350" number="2" />
                    <RELAYPOSITION athleteid="101314" number="3" />
                    <RELAYPOSITION athleteid="101311" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="10">
              <RESULTS>
                <RESULT comment="1 zmiana S 4" eventid="99059" reactiontime="+80" status="DSQ" swimtime="00:00:00.00" resultid="101369" heatid="105241" lane="3" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.41" />
                    <SPLIT distance="100" swimtime="00:01:13.79" />
                    <SPLIT distance="150" swimtime="00:01:41.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101311" number="1" reactiontime="+80" status="DSQ" />
                    <RELAYPOSITION athleteid="101273" number="2" reactiontime="-9" status="DSQ" />
                    <RELAYPOSITION athleteid="101350" number="3" reactiontime="+50" status="DSQ" />
                    <RELAYPOSITION athleteid="101321" number="4" reactiontime="+38" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="11">
              <RESULTS>
                <RESULT eventid="99250" points="305" reactiontime="+77" swimtime="00:02:05.93" resultid="101370" heatid="105310" lane="8" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.75" />
                    <SPLIT distance="100" swimtime="00:01:04.22" />
                    <SPLIT distance="150" swimtime="00:01:40.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101340" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="101321" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="101277" number="3" />
                    <RELAYPOSITION athleteid="101263" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="12">
              <RESULTS>
                <RESULT eventid="99036" status="DNS" swimtime="00:00:00.00" resultid="101371" heatid="105238" lane="6" entrytime="00:02:26.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101293" number="1" />
                    <RELAYPOSITION athleteid="101355" number="2" />
                    <RELAYPOSITION athleteid="101303" number="3" />
                    <RELAYPOSITION athleteid="101344" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="13">
              <RESULTS>
                <RESULT eventid="99234" status="DNS" swimtime="00:00:00.00" resultid="101372" heatid="105307" lane="2" entrytime="00:02:09.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101344" number="1" />
                    <RELAYPOSITION athleteid="101303" number="2" />
                    <RELAYPOSITION athleteid="101355" number="3" />
                    <RELAYPOSITION athleteid="101293" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="14">
              <RESULTS>
                <RESULT eventid="99036" points="258" reactiontime="+80" swimtime="00:02:46.54" resultid="101373" heatid="105237" lane="5" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.97" />
                    <SPLIT distance="100" swimtime="00:01:35.99" />
                    <SPLIT distance="150" swimtime="00:02:14.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101326" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="101296" number="2" reactiontime="+22" />
                    <RELAYPOSITION athleteid="101268" number="3" reactiontime="+26" />
                    <RELAYPOSITION athleteid="101308" number="4" reactiontime="+75" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="15">
              <RESULTS>
                <RESULT eventid="99234" points="281" reactiontime="+92" swimtime="00:02:27.59" resultid="101374" heatid="105306" lane="4" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                    <SPLIT distance="100" swimtime="00:01:19.24" />
                    <SPLIT distance="150" swimtime="00:01:54.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101268" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="101308" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="101326" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="101282" number="4" reactiontime="+77" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" status="DNS" swimtime="00:00:00.00" resultid="101360" heatid="105161" lane="5" entrytime="00:01:55.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101350" number="1" />
                    <RELAYPOSITION athleteid="101303" number="2" />
                    <RELAYPOSITION athleteid="101344" number="3" />
                    <RELAYPOSITION athleteid="101314" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="98846" points="393" reactiontime="+77" swimtime="00:01:55.83" resultid="101361" heatid="105161" lane="6" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.59" />
                    <SPLIT distance="100" swimtime="00:00:56.44" />
                    <SPLIT distance="150" swimtime="00:01:24.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101299" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="101268" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="101355" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="101263" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="99441" status="DNS" swimtime="00:00:00.00" resultid="101362" heatid="105365" lane="0" entrytime="00:02:16.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101303" number="1" />
                    <RELAYPOSITION athleteid="101299" number="2" />
                    <RELAYPOSITION athleteid="101317" number="3" />
                    <RELAYPOSITION athleteid="101355" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="98846" status="DNS" swimtime="00:00:00.00" resultid="101363" heatid="105160" lane="2" entrytime="00:02:13.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101321" number="1" />
                    <RELAYPOSITION athleteid="101293" number="2" />
                    <RELAYPOSITION athleteid="101308" number="3" />
                    <RELAYPOSITION athleteid="101340" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="5">
              <RESULTS>
                <RESULT eventid="99441" status="DNS" swimtime="00:00:00.00" resultid="101364" heatid="105364" lane="6" entrytime="00:02:25.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101340" number="1" />
                    <RELAYPOSITION athleteid="101273" number="2" />
                    <RELAYPOSITION athleteid="101268" number="3" />
                    <RELAYPOSITION athleteid="101308" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="6">
              <RESULTS>
                <RESULT eventid="98846" points="170" reactiontime="+117" swimtime="00:02:33.01" resultid="101365" heatid="105159" lane="7" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.21" />
                    <SPLIT distance="100" swimtime="00:01:11.34" />
                    <SPLIT distance="150" swimtime="00:01:57.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101287" number="1" reactiontime="+117" />
                    <RELAYPOSITION athleteid="101326" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="101282" number="3" reactiontime="+29" />
                    <RELAYPOSITION athleteid="101277" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="7">
              <RESULTS>
                <RESULT eventid="99441" points="151" reactiontime="+77" swimtime="00:02:55.20" resultid="101366" heatid="105363" lane="3" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.59" />
                    <SPLIT distance="100" swimtime="00:01:41.13" />
                    <SPLIT distance="150" swimtime="00:02:23.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101277" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="101296" number="2" reactiontime="+17" />
                    <RELAYPOSITION athleteid="101287" number="3" reactiontime="+77" />
                    <RELAYPOSITION athleteid="101282" number="4" reactiontime="+64" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="16">
              <RESULTS>
                <RESULT eventid="99441" points="331" reactiontime="+71" swimtime="00:02:15.00" resultid="101375" heatid="105365" lane="5" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.86" />
                    <SPLIT distance="100" swimtime="00:01:14.82" />
                    <SPLIT distance="150" swimtime="00:01:42.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101293" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="101263" number="2" reactiontime="+6" />
                    <RELAYPOSITION athleteid="101350" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="101344" number="4" reactiontime="+73" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="102935" name="Namysłów">
          <ATHLETES>
            <ATHLETE birthdate="1969-01-24" firstname="Katarzyna" gender="F" lastname="DOLAN" nation="POL" athleteid="102936">
              <RESULTS>
                <RESULT eventid="98777" points="376" swimtime="00:00:32.86" resultid="103426" heatid="105117" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="98907" points="366" reactiontime="+91" swimtime="00:00:37.80" resultid="103427" heatid="105177" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="99314" points="354" reactiontime="+98" swimtime="00:01:22.10" resultid="103428" heatid="105280" lane="0" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="327" reactiontime="+79" swimtime="00:03:00.01" resultid="103429" heatid="105334" lane="8" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.69" />
                    <SPLIT distance="100" swimtime="00:01:27.73" />
                    <SPLIT distance="150" swimtime="00:02:14.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ORSOPOLE" nation="POL" clubid="104386" name="Odrzańskie Ratownictwo Specjalistyczne Opole" shortname="ORS Opole">
          <CONTACT email="wkania62@gmail.com" name="Kania Waldemar" />
          <ATHLETES>
            <ATHLETE birthdate="1962-01-01" firstname="Waldemar" gender="M" lastname="KANIA" nation="POL" swrid="4302335" athleteid="104387">
              <RESULTS>
                <RESULT eventid="98891" points="265" swimtime="00:22:34.53" resultid="104388" heatid="105421" lane="9" entrytime="00:21:59.00" />
                <RESULT eventid="99218" points="257" reactiontime="+102" swimtime="00:02:40.42" resultid="104389" heatid="105300" lane="0" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                    <SPLIT distance="100" swimtime="00:01:17.10" />
                    <SPLIT distance="150" swimtime="00:01:59.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="174" reactiontime="+88" swimtime="00:03:20.35" resultid="104390" heatid="105338" lane="7" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.83" />
                    <SPLIT distance="100" swimtime="00:01:38.51" />
                    <SPLIT distance="150" swimtime="00:02:31.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="104391" entrytime="00:05:29.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02705" nation="POL" region="LOD" clubid="102224" name="Pływak Tomaszów Mazowiecki">
          <CONTACT email="tsplywak@wp.pl" name="Bucholz" phone="606 135 860" />
          <ATHLETES>
            <ATHLETE birthdate="1975-05-02" firstname="Bernard" gender="M" lastname="WIERZBIK" nation="POL" swrid="4992867" athleteid="102246">
              <RESULTS>
                <RESULT eventid="98830" points="214" reactiontime="+110" swimtime="00:03:10.55" resultid="102247" heatid="105152" lane="2" entrytime="00:03:04.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                    <SPLIT distance="100" swimtime="00:01:30.83" />
                    <SPLIT distance="150" swimtime="00:02:24.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="219" reactiontime="+105" swimtime="00:01:17.79" resultid="102248" heatid="105221" lane="1" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="241" reactiontime="+95" swimtime="00:00:36.01" resultid="102249" heatid="105270" lane="5" entrytime="00:00:33.82" />
                <RESULT eventid="99361" points="199" reactiontime="+94" swimtime="00:01:25.28" resultid="102250" heatid="105328" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-23" firstname="Bartek" gender="M" lastname="MASLOCHA" nation="POL" athleteid="102251">
              <RESULTS>
                <RESULT eventid="98798" points="195" reactiontime="+107" swimtime="00:00:36.02" resultid="102252" heatid="105128" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="98924" points="159" reactiontime="+72" swimtime="00:00:44.34" resultid="102253" heatid="105183" lane="4" entrytime="00:00:42.40" />
                <RESULT eventid="98988" points="166" reactiontime="+110" swimtime="00:01:25.32" resultid="102254" heatid="105216" lane="7" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="104" reactiontime="+126" swimtime="00:00:47.60" resultid="102255" heatid="105266" lane="3" entrytime="00:00:42.00" />
                <RESULT eventid="99425" points="146" reactiontime="+117" swimtime="00:00:50.56" resultid="102256" heatid="105353" lane="0" entrytime="00:00:46.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="RAAS+" nation="POL" clubid="100357" name="Rydułtowska Akademia A Seniora 60+" shortname="Rydułtowska Akademia">
          <CONTACT email="zurekt@poczta.onet.pl" name="Żurczak Tomasz" phone="504152136" />
          <ATHLETES>
            <ATHLETE birthdate="1940-05-16" firstname="Rudolf" gender="M" lastname="BUGLA" nation="POL" swrid="4831499" athleteid="100366">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="100367" heatid="105124" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="98830" points="78" reactiontime="+118" swimtime="00:04:26.04" resultid="100368" heatid="105149" lane="5" entrytime="00:04:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.87" />
                    <SPLIT distance="100" swimtime="00:02:10.16" />
                    <SPLIT distance="150" swimtime="00:03:24.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="76" reactiontime="+82" swimtime="00:00:56.66" resultid="100369" heatid="105181" lane="4" entrytime="00:00:52.00" />
                <RESULT eventid="99020" points="52" reactiontime="+108" swimtime="00:04:56.93" resultid="100370" heatid="105232" lane="3" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.33" />
                    <SPLIT distance="100" swimtime="00:02:14.20" />
                    <SPLIT distance="150" swimtime="00:03:31.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="100371" heatid="105266" lane="9" entrytime="00:00:49.00" />
                <RESULT eventid="99282" points="69" reactiontime="+110" swimtime="00:09:53.90" resultid="100372" heatid="106048" lane="0" entrytime="00:09:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.04" />
                    <SPLIT distance="100" swimtime="00:02:26.87" />
                    <SPLIT distance="150" swimtime="00:03:44.90" />
                    <SPLIT distance="200" swimtime="00:05:01.77" />
                    <SPLIT distance="250" swimtime="00:06:18.61" />
                    <SPLIT distance="300" swimtime="00:07:35.66" />
                    <SPLIT distance="350" swimtime="00:08:45.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="49" reactiontime="+109" swimtime="00:02:15.59" resultid="100373" heatid="105325" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="71" reactiontime="+93" swimtime="00:04:30.23" resultid="100374" heatid="105336" lane="5" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.45" />
                    <SPLIT distance="100" swimtime="00:02:13.71" />
                    <SPLIT distance="150" swimtime="00:03:23.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-11-24" firstname="Jerzy" gender="M" lastname="CIECIOR" nation="POL" swrid="4934027" athleteid="100375">
              <RESULTS>
                <RESULT eventid="98830" points="184" reactiontime="+107" swimtime="00:03:20.31" resultid="100376" heatid="105151" lane="6" entrytime="00:03:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.95" />
                    <SPLIT distance="100" swimtime="00:01:32.01" />
                    <SPLIT distance="150" swimtime="00:02:34.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="195" swimtime="00:25:01.78" resultid="100377" heatid="105423" lane="1" entrytime="00:24:40.00" />
                <RESULT eventid="98924" points="189" reactiontime="+82" swimtime="00:00:41.87" resultid="100378" heatid="105184" lane="6" entrytime="00:00:41.00" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="100379" heatid="105217" lane="7" entrytime="00:01:14.00" />
                <RESULT eventid="99170" points="217" reactiontime="+86" swimtime="00:00:37.28" resultid="100380" heatid="105268" lane="0" entrytime="00:00:37.00" />
                <RESULT eventid="99186" points="148" reactiontime="+100" swimtime="00:01:38.09" resultid="100381" heatid="105283" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="168" reactiontime="+94" swimtime="00:01:30.26" resultid="100382" heatid="105327" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="161" reactiontime="+101" swimtime="00:03:25.66" resultid="100383" heatid="105338" lane="2" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.98" />
                    <SPLIT distance="100" swimtime="00:01:40.10" />
                    <SPLIT distance="150" swimtime="00:02:34.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-09-07" firstname="Leon" gender="M" lastname="IRCZYK" nation="POL" swrid="4934026" athleteid="100384">
              <RESULTS>
                <RESULT eventid="98830" points="91" reactiontime="+136" swimtime="00:04:12.88" resultid="100385" heatid="105149" lane="1" entrytime="00:04:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.00" />
                    <SPLIT distance="100" swimtime="00:02:15.01" />
                    <SPLIT distance="150" swimtime="00:03:16.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="100" swimtime="00:31:15.00" resultid="100386" heatid="105425" lane="6" entrytime="00:31:00.00" />
                <RESULT eventid="98956" points="162" reactiontime="+118" swimtime="00:03:52.82" resultid="100387" heatid="105197" lane="9" entrytime="00:04:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.88" />
                    <SPLIT distance="100" swimtime="00:01:54.76" />
                    <SPLIT distance="150" swimtime="00:02:55.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="52" reactiontime="+130" swimtime="00:04:57.93" resultid="100388" heatid="105232" lane="9" entrytime="00:05:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.80" />
                    <SPLIT distance="100" swimtime="00:02:19.74" />
                    <SPLIT distance="150" swimtime="00:03:37.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="160" reactiontime="+136" swimtime="00:01:47.67" resultid="100389" heatid="105250" lane="6" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="86" reactiontime="+133" swimtime="00:09:10.64" resultid="100390" heatid="106048" lane="7" entrytime="00:08:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.88" />
                    <SPLIT distance="100" swimtime="00:02:16.36" />
                    <SPLIT distance="150" swimtime="00:03:40.25" />
                    <SPLIT distance="200" swimtime="00:04:59.91" />
                    <SPLIT distance="250" swimtime="00:06:03.54" />
                    <SPLIT distance="300" swimtime="00:07:06.45" />
                    <SPLIT distance="350" swimtime="00:08:08.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="49" reactiontime="+120" swimtime="00:05:05.16" resultid="100391" heatid="105337" lane="1" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.75" />
                    <SPLIT distance="100" swimtime="00:02:32.41" />
                    <SPLIT distance="150" swimtime="00:03:49.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="97" reactiontime="+134" swimtime="00:07:58.60" resultid="100392" heatid="106066" lane="1" entrytime="00:07:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.45" />
                    <SPLIT distance="100" swimtime="00:01:53.19" />
                    <SPLIT distance="150" swimtime="00:02:54.40" />
                    <SPLIT distance="200" swimtime="00:03:56.76" />
                    <SPLIT distance="250" swimtime="00:04:58.22" />
                    <SPLIT distance="300" swimtime="00:05:58.78" />
                    <SPLIT distance="350" swimtime="00:06:59.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="SUI" clubid="100102" name="Schwimmverein beider Basel (SVB)">
          <CONTACT city="Basel" email="quiri.zumbach@yetnet.ch" name="Swen Schubert" street="Postfach 73" zip="4020" />
          <ATHLETES>
            <ATHLETE birthdate="1977-03-27" firstname="Swen" gender="M" lastname="SCHUBERT" nation="SUI" swrid="4870232" athleteid="100103">
              <RESULTS>
                <RESULT eventid="98798" points="288" reactiontime="+80" swimtime="00:00:31.64" resultid="100104" heatid="105130" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="98830" points="242" reactiontime="+77" swimtime="00:03:02.92" resultid="100105" heatid="105152" lane="7" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                    <SPLIT distance="100" swimtime="00:01:28.56" />
                    <SPLIT distance="150" swimtime="00:02:22.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="248" reactiontime="+78" swimtime="00:00:38.22" resultid="100106" heatid="105179" lane="3" />
                <RESULT eventid="98988" points="286" reactiontime="+75" swimtime="00:01:11.15" resultid="100107" heatid="105218" lane="6" entrytime="00:01:10.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="227" reactiontime="+88" swimtime="00:00:36.74" resultid="100108" heatid="105268" lane="2" entrytime="00:00:36.46" />
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="100109" heatid="105299" lane="7" entrytime="00:02:40.35" />
                <RESULT eventid="99361" points="158" reactiontime="+91" swimtime="00:01:32.12" resultid="100110" heatid="105326" lane="3" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="188" reactiontime="+72" swimtime="00:03:15.08" resultid="100111" heatid="105335" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.93" />
                    <SPLIT distance="100" swimtime="00:01:35.74" />
                    <SPLIT distance="150" swimtime="00:02:27.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-03-21" firstname="Quirina" gender="F" lastname="ZUMBACH" nation="SUI" swrid="4895263" athleteid="100112">
              <RESULTS>
                <RESULT eventid="98777" status="DNS" swimtime="00:00:00.00" resultid="100113" heatid="105118" lane="0" entrytime="00:00:34.00" />
                <RESULT eventid="98940" status="DNS" swimtime="00:00:00.00" resultid="100114" heatid="105192" lane="3" entrytime="00:03:47.26" />
                <RESULT eventid="98972" points="230" reactiontime="+76" swimtime="00:01:24.88" resultid="100115" heatid="105208" lane="9" entrytime="00:01:21.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="211" reactiontime="+89" swimtime="00:01:48.05" resultid="100116" heatid="105245" lane="5" entrytime="00:01:42.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="233" reactiontime="+81" swimtime="00:00:47.86" resultid="100117" heatid="105346" lane="6" entrytime="00:00:47.17" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="102767" name="Sikret Gliwice">
          <CONTACT city="GLIWICE" email="joannaeco@tlen.pl" internet="www.sikret-plywnie.pl" name="JOANNA ZAGAŁA" phone="601427257" street="JAGIELOŃSKA 21" zip="44-100" />
          <ATHLETES>
            <ATHLETE birthdate="1958-02-05" firstname="Zofia" gender="F" lastname="DĄBROWSKA" nation="POL" swrid="4934035" athleteid="102777">
              <RESULTS>
                <RESULT eventid="98777" points="183" reactiontime="+82" swimtime="00:00:41.73" resultid="102778" heatid="105114" lane="6" entrytime="00:00:41.81" entrycourse="SCM" />
                <RESULT eventid="98814" points="110" reactiontime="+97" swimtime="00:04:22.73" resultid="102779" heatid="105144" lane="1" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.38" />
                    <SPLIT distance="100" swimtime="00:02:20.22" />
                    <SPLIT distance="150" swimtime="00:03:23.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="162" reactiontime="+85" swimtime="00:04:15.05" resultid="102780" heatid="105192" lane="9" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.97" />
                    <SPLIT distance="100" swimtime="00:02:02.49" />
                    <SPLIT distance="150" swimtime="00:03:10.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99004" status="DNS" swimtime="00:00:00.00" resultid="102781" heatid="105229" lane="6" entrytime="00:05:00.00" />
                <RESULT eventid="99089" points="166" reactiontime="+90" swimtime="00:01:56.96" resultid="102782" heatid="105244" lane="6" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="109" reactiontime="+83" swimtime="00:00:52.47" resultid="102783" heatid="105259" lane="7" entrytime="00:00:52.10" />
                <RESULT eventid="99344" points="84" reactiontime="+90" swimtime="00:02:07.48" resultid="102784" heatid="105321" lane="2" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="183" reactiontime="+91" swimtime="00:00:51.86" resultid="102785" heatid="105345" lane="1" entrytime="00:00:53.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-06-24" firstname="Joanna" gender="F" lastname="ZAGAŁA" nation="POL" swrid="4934034" athleteid="102786">
              <RESULTS>
                <RESULT eventid="98777" points="221" reactiontime="+84" swimtime="00:00:39.24" resultid="102787" heatid="105115" lane="1" entrytime="00:00:39.23" entrycourse="LCM" />
                <RESULT eventid="98814" points="166" reactiontime="+77" swimtime="00:03:49.44" resultid="102788" heatid="105144" lane="7" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.66" />
                    <SPLIT distance="100" swimtime="00:01:54.49" />
                    <SPLIT distance="150" swimtime="00:02:56.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="150" reactiontime="+86" swimtime="00:00:50.82" resultid="102789" heatid="105173" lane="2" entrytime="00:00:52.00" />
                <RESULT eventid="98940" points="180" reactiontime="+114" swimtime="00:04:06.29" resultid="102790" heatid="105192" lane="0" entrytime="00:04:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.31" />
                    <SPLIT distance="100" swimtime="00:02:00.55" />
                    <SPLIT distance="150" swimtime="00:03:04.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="189" reactiontime="+76" swimtime="00:01:51.96" resultid="102791" heatid="105244" lane="7" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="163" reactiontime="+73" swimtime="00:03:26.67" resultid="102792" heatid="105290" lane="9" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.65" />
                    <SPLIT distance="100" swimtime="00:01:40.57" />
                    <SPLIT distance="150" swimtime="00:02:36.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="144" reactiontime="+78" swimtime="00:03:56.63" resultid="102793" heatid="105332" lane="6" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.76" />
                    <SPLIT distance="100" swimtime="00:01:57.83" />
                    <SPLIT distance="150" swimtime="00:02:58.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="203" reactiontime="+81" swimtime="00:00:50.16" resultid="102794" heatid="105345" lane="3" entrytime="00:00:51.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-08-11" firstname="Agnieszka" gender="F" lastname="DREJKA" nation="POL" athleteid="102795">
              <RESULTS>
                <RESULT eventid="98777" points="173" reactiontime="+107" swimtime="00:00:42.55" resultid="102796" heatid="105114" lane="9" entrytime="00:00:44.00" />
                <RESULT eventid="98940" points="187" reactiontime="+104" swimtime="00:04:02.96" resultid="102797" heatid="105191" lane="4" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.09" />
                    <SPLIT distance="100" swimtime="00:01:56.01" />
                    <SPLIT distance="150" swimtime="00:02:59.78" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="04" eventid="99089" reactiontime="+43" status="DSQ" swimtime="00:01:53.50" resultid="102798" heatid="105244" lane="5" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="175" reactiontime="+111" swimtime="00:00:52.64" resultid="102799" heatid="105344" lane="4" entrytime="00:00:54.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SOPMAST" nation="POL" region="POM" clubid="101949" name="Sopot Masters">
          <CONTACT city="SOPOT" email="sopotmasters@o2.pl" internet="strona www chwilowo nieczynna" name="Gorbaczow Mirosław" phone="696 258 185" state="POMOR" street="ul. Haffnera 57" zip="81-715" />
          <ATHLETES>
            <ATHLETE birthdate="1958-12-28" firstname="Dariusz" gender="M" lastname="GORBACZOW" nation="POL" swrid="4191113" athleteid="102826">
              <RESULTS>
                <RESULT eventid="98798" points="345" reactiontime="+77" swimtime="00:00:29.79" resultid="102827" heatid="105133" lane="9" entrytime="00:00:30.40" entrycourse="LCM" />
                <RESULT eventid="98924" points="329" reactiontime="+101" swimtime="00:00:34.80" resultid="102828" heatid="105187" lane="1" entrytime="00:00:34.60" entrycourse="LCM" />
                <RESULT eventid="98988" points="357" reactiontime="+85" swimtime="00:01:06.07" resultid="102829" heatid="105221" lane="8" entrytime="00:01:07.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="393" reactiontime="+77" swimtime="00:00:30.60" resultid="102830" heatid="105272" lane="8" entrytime="00:00:31.20" entrycourse="LCM" />
                <RESULT eventid="99186" points="293" reactiontime="+93" swimtime="00:01:18.18" resultid="102831" heatid="105285" lane="0" entrytime="00:01:18.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="102832" heatid="105340" lane="9" entrytime="00:02:58.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-02-08" firstname="Anna" gender="F" lastname="MACIEJOWSKA" nation="POL" swrid="4191115" athleteid="102833">
              <RESULTS>
                <RESULT eventid="98777" points="280" reactiontime="+91" swimtime="00:00:36.23" resultid="102834" heatid="105118" lane="6" entrytime="00:00:33.03" entrycourse="LCM" />
                <RESULT eventid="98863" points="207" swimtime="00:13:53.64" resultid="102835" heatid="105406" lane="4" entrytime="00:14:00.00" entrycourse="LCM" />
                <RESULT eventid="98972" status="DNS" swimtime="00:00:00.00" resultid="102836" heatid="105208" lane="0" entrytime="00:01:21.00" entrycourse="LCM" />
                <RESULT eventid="99202" status="DNS" swimtime="00:00:00.00" resultid="102837" heatid="105291" lane="0" entrytime="00:03:06.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SQUOST" nation="POL" region="WAR" clubid="101240" name="Squatina Ostrołęka">
          <CONTACT city="Ostrołęka" email="biezunskamaja@gmail.com" name="Bieżuńska Maja" phone="666-353-028" state="MAZ" street="Łęczysk 10/14/26" zip="07-410" />
          <ATHLETES>
            <ATHLETE birthdate="1979-06-26" firstname="Maja" gender="F" lastname="BIEŻUŃSKA" nation="POL" swrid="4992888" athleteid="101241">
              <RESULTS>
                <RESULT eventid="98940" points="330" reactiontime="+99" swimtime="00:03:21.11" resultid="101242" heatid="105194" lane="3" entrytime="00:03:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.52" />
                    <SPLIT distance="100" swimtime="00:01:35.13" />
                    <SPLIT distance="150" swimtime="00:02:27.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="366" reactiontime="+90" swimtime="00:01:29.93" resultid="101243" heatid="105247" lane="3" entrytime="00:01:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="398" reactiontime="+89" swimtime="00:00:40.05" resultid="101244" heatid="105348" lane="5" entrytime="00:00:40.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="WIE" clubid="104962" name="Start Poznań">
          <CONTACT city="Poznań" email="robert.beym@gmail.com" name="Beym Robert" phone="+48 512111513" street="os. Stefana Batorego 8,67" zip="60-687" />
          <ATHLETES>
            <ATHLETE birthdate="1969-02-26" firstname="Robert" gender="M" lastname="BEYM" nation="POL" swrid="4992890" athleteid="104963">
              <RESULTS>
                <RESULT eventid="98798" points="426" reactiontime="+93" swimtime="00:00:27.78" resultid="104964" heatid="105134" lane="0" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT eventid="98891" points="313" swimtime="00:21:21.57" resultid="104965" heatid="105422" lane="9" entrytime="00:23:00.00" entrycourse="LCM" />
                <RESULT eventid="98924" points="393" reactiontime="+86" swimtime="00:00:32.80" resultid="104966" heatid="105186" lane="1" entrytime="00:00:36.00" entrycourse="LCM" />
                <RESULT eventid="98988" points="435" reactiontime="+98" swimtime="00:01:01.90" resultid="104967" heatid="105224" lane="2" entrytime="00:01:02.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="395" reactiontime="+83" swimtime="00:01:10.78" resultid="104968" heatid="105287" lane="0" entrytime="00:01:11.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.51" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G6" eventid="99393" reactiontime="+82" status="DSQ" swimtime="00:00:00.00" resultid="104969" heatid="105339" lane="7" entrytime="00:03:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.92" />
                    <SPLIT distance="100" swimtime="00:01:14.71" />
                    <SPLIT distance="150" swimtime="00:01:55.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="104970" entrytime="00:05:30.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-02-26" firstname="Piotr" gender="M" lastname="MOŃCZAK" nation="POL" athleteid="104971">
              <RESULTS>
                <RESULT eventid="98798" points="445" reactiontime="+72" swimtime="00:00:27.37" resultid="104972" heatid="105141" lane="9" entrytime="00:00:27.00" entrycourse="LCM" />
                <RESULT eventid="98830" points="406" reactiontime="+72" swimtime="00:02:33.88" resultid="104973" heatid="105157" lane="9" entrytime="00:02:32.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                    <SPLIT distance="100" swimtime="00:01:13.53" />
                    <SPLIT distance="150" swimtime="00:01:58.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="506" reactiontime="+88" swimtime="00:00:58.84" resultid="104974" heatid="105226" lane="0" entrytime="00:00:59.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="445" reactiontime="+88" swimtime="00:02:13.54" resultid="104975" heatid="105304" lane="2" entrytime="00:02:12.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                    <SPLIT distance="100" swimtime="00:01:05.33" />
                    <SPLIT distance="150" swimtime="00:01:41.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="425" reactiontime="+95" swimtime="00:04:52.48" resultid="104976" heatid="106060" lane="0" entrytime="00:04:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                    <SPLIT distance="100" swimtime="00:01:10.63" />
                    <SPLIT distance="150" swimtime="00:01:47.38" />
                    <SPLIT distance="200" swimtime="00:02:25.16" />
                    <SPLIT distance="250" swimtime="00:03:02.63" />
                    <SPLIT distance="300" swimtime="00:03:41.29" />
                    <SPLIT distance="350" swimtime="00:04:17.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-02-26" firstname="Krzysztof" gender="M" lastname="KAPAŁCZYŃSKI" nation="POL" athleteid="104977">
              <RESULTS>
                <RESULT eventid="98830" points="308" reactiontime="+82" swimtime="00:02:48.67" resultid="104978" heatid="105153" lane="9" entrytime="00:02:58.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                    <SPLIT distance="100" swimtime="00:01:19.33" />
                    <SPLIT distance="150" swimtime="00:02:08.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="209" reactiontime="+96" swimtime="00:03:07.85" resultid="104979" heatid="105234" lane="5" entrytime="00:03:08.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.38" />
                    <SPLIT distance="100" swimtime="00:01:30.03" />
                    <SPLIT distance="150" swimtime="00:02:20.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="288" reactiontime="+87" swimtime="00:06:08.90" resultid="104980" heatid="106051" lane="7" entrytime="00:06:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                    <SPLIT distance="100" swimtime="00:01:21.95" />
                    <SPLIT distance="150" swimtime="00:02:10.17" />
                    <SPLIT distance="200" swimtime="00:02:56.76" />
                    <SPLIT distance="250" swimtime="00:03:50.85" />
                    <SPLIT distance="300" swimtime="00:04:43.98" />
                    <SPLIT distance="350" swimtime="00:05:27.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="263" reactiontime="+97" swimtime="00:01:17.75" resultid="104981" heatid="105328" lane="1" entrytime="00:01:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="304" reactiontime="+87" swimtime="00:00:39.63" resultid="104982" heatid="105353" lane="7" entrytime="00:00:45.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="MAZ" clubid="102871" name="Swimmers SP Warszawa">
          <CONTACT city="WARSZAWA" email="info@swimmersteam.pl" internet="www.swimmersteam.pl" name="GOŁĘBIOWSKI REMIGIUSZ" phone="601333782" state="MAZ" street="GŁADKA 18" zip="02-172" />
          <ATHLETES>
            <ATHLETE birthdate="1976-07-07" firstname="Remigiusz" gender="M" lastname="GOŁĘBIOWSKI" nation="POL" swrid="4743284" athleteid="102879">
              <RESULTS>
                <RESULT eventid="98798" points="450" reactiontime="+87" swimtime="00:00:27.28" resultid="102880" heatid="105140" lane="7" entrytime="00:00:27.00" entrycourse="LCM" />
                <RESULT eventid="98891" points="426" swimtime="00:19:16.70" resultid="102881" heatid="105420" lane="2" entrytime="00:19:30.00" entrycourse="LCM" />
                <RESULT eventid="99170" points="432" reactiontime="+91" swimtime="00:00:29.66" resultid="102882" heatid="105275" lane="0" entrytime="00:00:28.00" entrycourse="LCM" />
                <RESULT eventid="99218" points="430" reactiontime="+96" swimtime="00:02:15.04" resultid="102883" heatid="105305" lane="0" entrytime="00:02:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                    <SPLIT distance="100" swimtime="00:01:02.99" />
                    <SPLIT distance="150" swimtime="00:01:38.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="441" reactiontime="+95" swimtime="00:04:49.09" resultid="102884" heatid="106059" lane="0" entrytime="00:04:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.85" />
                    <SPLIT distance="100" swimtime="00:01:08.82" />
                    <SPLIT distance="150" swimtime="00:01:46.22" />
                    <SPLIT distance="200" swimtime="00:02:23.35" />
                    <SPLIT distance="250" swimtime="00:03:00.55" />
                    <SPLIT distance="300" swimtime="00:03:37.68" />
                    <SPLIT distance="350" swimtime="00:04:14.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-08-29" firstname="Marek" gender="M" lastname="BROŻYNA" nation="POL" athleteid="102885">
              <RESULTS>
                <RESULT eventid="98798" points="314" reactiontime="+104" swimtime="00:00:30.74" resultid="102886" heatid="105135" lane="7" entrytime="00:00:29.50" entrycourse="LCM" />
                <RESULT eventid="98924" points="334" reactiontime="+63" swimtime="00:00:34.63" resultid="102887" heatid="105187" lane="6" entrytime="00:00:34.00" entrycourse="LCM" />
                <RESULT eventid="99186" points="294" reactiontime="+77" swimtime="00:01:18.11" resultid="102888" heatid="105286" lane="9" entrytime="00:01:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="288" reactiontime="+85" swimtime="00:02:49.31" resultid="102889" heatid="105341" lane="1" entrytime="00:02:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.94" />
                    <SPLIT distance="100" swimtime="00:01:21.78" />
                    <SPLIT distance="150" swimtime="00:02:06.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-12-11" firstname="Mikołaj" gender="M" lastname="TUSIŃSKI" nation="POL" athleteid="102890">
              <RESULTS>
                <RESULT eventid="98798" points="385" reactiontime="+88" swimtime="00:00:28.72" resultid="102891" heatid="105137" lane="7" entrytime="00:00:28.50" entrycourse="LCM" />
                <RESULT eventid="98988" points="427" reactiontime="+94" swimtime="00:01:02.27" resultid="102892" heatid="105224" lane="0" entrytime="00:01:02.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="408" reactiontime="+89" swimtime="00:00:30.24" resultid="102893" heatid="105274" lane="1" entrytime="00:00:29.80" entrycourse="LCM" />
                <RESULT eventid="99218" points="353" reactiontime="+85" swimtime="00:02:24.22" resultid="102894" heatid="105304" lane="4" entrytime="00:02:10.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.60" />
                    <SPLIT distance="100" swimtime="00:01:04.97" />
                    <SPLIT distance="150" swimtime="00:01:43.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-07-29" firstname="Urszula" gender="F" lastname="JAKUBOWSKA CŁAPIŃSKA" nation="POL" athleteid="102895">
              <RESULTS>
                <RESULT eventid="98814" points="213" reactiontime="+102" swimtime="00:03:31.08" resultid="102896" heatid="105146" lane="3" entrytime="00:02:59.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.03" />
                    <SPLIT distance="100" swimtime="00:01:37.91" />
                    <SPLIT distance="150" swimtime="00:02:41.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="249" reactiontime="+86" swimtime="00:00:42.96" resultid="102897" heatid="105175" lane="1" entrytime="00:00:42.00" entrycourse="LCM" />
                <RESULT eventid="98972" points="246" reactiontime="+102" swimtime="00:01:23.01" resultid="102898" heatid="105210" lane="1" entrytime="00:01:12.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="216" reactiontime="+103" swimtime="00:03:08.19" resultid="102899" heatid="105293" lane="2" entrytime="00:02:35.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.03" />
                    <SPLIT distance="100" swimtime="00:01:27.13" />
                    <SPLIT distance="150" swimtime="00:02:17.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-12-20" firstname="Arkadiusz" gender="M" lastname="APTEWICZ" nation="POL" swrid="4806379" athleteid="102900">
              <RESULTS>
                <RESULT eventid="98830" points="562" reactiontime="+68" swimtime="00:02:18.08" resultid="102901" heatid="105158" lane="8" entrytime="00:02:23.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.44" />
                    <SPLIT distance="100" swimtime="00:01:06.18" />
                    <SPLIT distance="150" swimtime="00:01:44.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="578" reactiontime="+78" swimtime="00:02:32.39" resultid="102902" heatid="105204" lane="2" entrytime="00:02:37.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.14" />
                    <SPLIT distance="100" swimtime="00:01:15.04" />
                    <SPLIT distance="150" swimtime="00:01:53.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="505" reactiontime="+72" swimtime="00:00:58.89" resultid="102903" heatid="105227" lane="4" entrytime="00:00:57.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="595" reactiontime="+79" swimtime="00:01:09.48" resultid="102904" heatid="105258" lane="1" entrytime="00:01:10.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="504" reactiontime="+81" swimtime="00:02:08.13" resultid="102905" heatid="105305" lane="2" entrytime="00:02:08.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.47" />
                    <SPLIT distance="100" swimtime="00:01:02.47" />
                    <SPLIT distance="150" swimtime="00:01:35.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="608" reactiontime="+65" swimtime="00:00:31.47" resultid="102906" heatid="105362" lane="9" entrytime="00:00:32.30" entrycourse="LCM" />
                <RESULT eventid="99473" points="493" reactiontime="+89" swimtime="00:04:38.51" resultid="102907" heatid="106059" lane="2" entrytime="00:04:32.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                    <SPLIT distance="100" swimtime="00:01:07.18" />
                    <SPLIT distance="150" swimtime="00:01:42.82" />
                    <SPLIT distance="200" swimtime="00:02:19.30" />
                    <SPLIT distance="250" swimtime="00:02:54.75" />
                    <SPLIT distance="300" swimtime="00:03:29.84" />
                    <SPLIT distance="350" swimtime="00:04:04.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-11-10" firstname="Anna" gender="F" lastname="TURCZYN" nation="POL" athleteid="102908">
              <RESULTS>
                <RESULT eventid="98777" status="DNS" swimtime="00:00:00.00" resultid="102909" heatid="105113" lane="5" entrytime="00:00:45.00" />
                <RESULT eventid="99409" status="DNS" swimtime="00:00:00.00" resultid="102910" heatid="105344" lane="5" entrytime="00:00:55.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="99441" points="233" reactiontime="+66" swimtime="00:02:31.69" resultid="106117" heatid="105363" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.62" />
                    <SPLIT distance="100" swimtime="00:01:24.41" />
                    <SPLIT distance="150" swimtime="00:01:26.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102885" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="102908" number="2" reactiontime="+78" />
                    <RELAYPOSITION athleteid="102895" number="3" />
                    <RELAYPOSITION athleteid="102890" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="100275" name="Swimming Masters Team Szczecin" shortname="Swim.Mrs Team Szczecin">
          <CONTACT name="Brodacki Maciej" />
          <ATHLETES>
            <ATHLETE birthdate="1983-02-24" firstname="Maciej" gender="M" lastname="BRODACKI" nation="POL" swrid="4751547" athleteid="100276">
              <RESULTS>
                <RESULT eventid="98798" points="480" reactiontime="+88" swimtime="00:00:26.69" resultid="100277" heatid="105141" lane="1" entrytime="00:00:26.50" />
                <RESULT eventid="98830" points="426" reactiontime="+82" swimtime="00:02:31.49" resultid="100278" heatid="105157" lane="7" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                    <SPLIT distance="100" swimtime="00:01:09.28" />
                    <SPLIT distance="150" swimtime="00:01:56.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="525" reactiontime="+80" swimtime="00:00:58.14" resultid="100279" heatid="105227" lane="7" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="403" reactiontime="+79" swimtime="00:02:17.98" resultid="100280" heatid="105302" lane="9" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.37" />
                    <SPLIT distance="100" swimtime="00:01:05.08" />
                    <SPLIT distance="150" swimtime="00:01:41.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="365" reactiontime="+90" swimtime="00:05:41.18" resultid="100281" heatid="106052" lane="5" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                    <SPLIT distance="100" swimtime="00:01:12.89" />
                    <SPLIT distance="150" swimtime="00:01:57.67" />
                    <SPLIT distance="200" swimtime="00:02:42.80" />
                    <SPLIT distance="250" swimtime="00:03:33.43" />
                    <SPLIT distance="300" swimtime="00:04:24.39" />
                    <SPLIT distance="350" swimtime="00:05:04.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="382" reactiontime="+94" swimtime="00:05:03.17" resultid="100282" heatid="106061" lane="0" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.97" />
                    <SPLIT distance="100" swimtime="00:01:10.82" />
                    <SPLIT distance="150" swimtime="00:01:48.96" />
                    <SPLIT distance="200" swimtime="00:02:27.40" />
                    <SPLIT distance="250" swimtime="00:03:06.41" />
                    <SPLIT distance="300" swimtime="00:03:46.41" />
                    <SPLIT distance="350" swimtime="00:04:26.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-02-27" firstname="Szymon" gender="M" lastname="KLUCZYK" nation="POL" swrid="4967270" athleteid="100283">
              <RESULTS>
                <RESULT eventid="98830" points="418" reactiontime="+94" swimtime="00:02:32.43" resultid="100284" heatid="105156" lane="1" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.89" />
                    <SPLIT distance="100" swimtime="00:01:11.23" />
                    <SPLIT distance="150" swimtime="00:01:56.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="423" swimtime="00:19:20.26" resultid="100285" heatid="105420" lane="4" entrytime="00:18:30.00" />
                <RESULT eventid="98956" status="DNS" swimtime="00:00:00.00" resultid="100286" heatid="105202" lane="8" entrytime="00:03:05.00" />
                <RESULT eventid="99020" points="354" reactiontime="+108" swimtime="00:02:37.49" resultid="100287" heatid="105236" lane="1" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="100" swimtime="00:01:14.98" />
                    <SPLIT distance="150" swimtime="00:01:58.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="410" reactiontime="+103" swimtime="00:05:28.04" resultid="100288" heatid="106053" lane="3" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                    <SPLIT distance="100" swimtime="00:01:10.71" />
                    <SPLIT distance="150" swimtime="00:01:54.41" />
                    <SPLIT distance="200" swimtime="00:02:37.13" />
                    <SPLIT distance="250" swimtime="00:03:26.01" />
                    <SPLIT distance="300" swimtime="00:04:15.13" />
                    <SPLIT distance="350" swimtime="00:04:51.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="449" reactiontime="+101" swimtime="00:04:47.38" resultid="100289" heatid="106059" lane="1" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.55" />
                    <SPLIT distance="100" swimtime="00:01:05.82" />
                    <SPLIT distance="150" swimtime="00:01:42.37" />
                    <SPLIT distance="200" swimtime="00:02:19.36" />
                    <SPLIT distance="250" swimtime="00:02:56.60" />
                    <SPLIT distance="300" swimtime="00:03:34.34" />
                    <SPLIT distance="350" swimtime="00:04:11.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-07-13" firstname="Piotr" gender="M" lastname="KOZŁOWSKI" nation="POL" athleteid="100290">
              <RESULTS>
                <RESULT eventid="98798" points="367" reactiontime="+80" swimtime="00:00:29.20" resultid="100291" heatid="105136" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="98988" points="370" reactiontime="+95" swimtime="00:01:05.32" resultid="100292" heatid="105222" lane="4" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="267" reactiontime="+96" swimtime="00:01:17.32" resultid="100293" heatid="105330" lane="1" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-25" firstname="Rafał" gender="M" lastname="LISIECKI" nation="POL" swrid="4992891" athleteid="100294">
              <RESULTS>
                <RESULT eventid="98798" points="435" reactiontime="+90" swimtime="00:00:27.59" resultid="100295" heatid="105139" lane="4" entrytime="00:00:27.30" />
                <RESULT eventid="98924" points="441" reactiontime="+84" swimtime="00:00:31.58" resultid="100296" heatid="105189" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="98988" points="470" reactiontime="+84" swimtime="00:01:00.32" resultid="100297" heatid="105224" lane="7" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="413" swimtime="00:01:09.74" resultid="100298" heatid="105287" lane="6" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-18" firstname="Jan" gender="M" lastname="ROENIG" nation="POL" swrid="4967271" athleteid="100299">
              <RESULTS>
                <RESULT eventid="98956" status="DNS" swimtime="00:00:00.00" resultid="100300" heatid="105203" lane="0" entrytime="00:02:59.00" />
                <RESULT eventid="99091" points="356" reactiontime="+98" swimtime="00:01:22.42" resultid="100301" heatid="105257" lane="1" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="403" reactiontime="+87" swimtime="00:00:36.09" resultid="100302" heatid="105361" lane="7" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-03-05" firstname="Rafał" gender="M" lastname="DOBROWOLSKI" nation="POL" athleteid="100303">
              <RESULTS>
                <RESULT eventid="98798" points="275" reactiontime="+80" swimtime="00:00:32.15" resultid="100304" heatid="105129" lane="3" entrytime="00:00:32.89" />
                <RESULT eventid="98924" status="DNS" swimtime="00:00:00.00" resultid="100305" heatid="105188" lane="0" entrytime="00:00:33.00" />
                <RESULT eventid="98988" points="203" reactiontime="+85" swimtime="00:01:19.71" resultid="100306" heatid="105228" lane="5" entrytime="00:00:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="100307" heatid="105258" lane="7" entrytime="00:01:10.00" />
                <RESULT eventid="99425" points="251" reactiontime="+99" swimtime="00:00:42.24" resultid="100308" heatid="105360" lane="1" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-20" firstname="Agnieszka" gender="F" lastname="KRZYŻOSTANIAK" nation="POL" swrid="4087097" athleteid="100309">
              <RESULTS>
                <RESULT eventid="98777" points="425" reactiontime="+91" swimtime="00:00:31.56" resultid="100310" heatid="105121" lane="2" entrytime="00:00:28.95" entrycourse="LCM" />
                <RESULT eventid="98863" points="506" reactiontime="+88" swimtime="00:10:19.51" resultid="100311" heatid="105404" lane="5" entrytime="00:10:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                    <SPLIT distance="100" swimtime="00:01:09.65" />
                    <SPLIT distance="150" swimtime="00:01:47.51" />
                    <SPLIT distance="200" swimtime="00:02:26.04" />
                    <SPLIT distance="250" swimtime="00:03:04.23" />
                    <SPLIT distance="300" swimtime="00:03:43.27" />
                    <SPLIT distance="350" swimtime="00:04:22.96" />
                    <SPLIT distance="400" swimtime="00:05:02.87" />
                    <SPLIT distance="450" swimtime="00:05:42.45" />
                    <SPLIT distance="500" swimtime="00:06:21.99" />
                    <SPLIT distance="550" swimtime="00:07:02.06" />
                    <SPLIT distance="600" swimtime="00:07:41.91" />
                    <SPLIT distance="650" swimtime="00:08:21.45" />
                    <SPLIT distance="700" swimtime="00:09:02.33" />
                    <SPLIT distance="750" swimtime="00:09:41.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="587" reactiontime="+76" swimtime="00:00:32.31" resultid="100312" heatid="105178" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="99154" points="439" reactiontime="+85" swimtime="00:00:32.98" resultid="100313" heatid="105263" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="99314" points="517" swimtime="00:01:12.39" resultid="100314" heatid="105280" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="530" reactiontime="+82" swimtime="00:04:55.48" resultid="100315" heatid="106054" lane="8" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                    <SPLIT distance="100" swimtime="00:01:09.06" />
                    <SPLIT distance="150" swimtime="00:01:46.11" />
                    <SPLIT distance="200" swimtime="00:02:24.07" />
                    <SPLIT distance="250" swimtime="00:03:01.85" />
                    <SPLIT distance="300" swimtime="00:03:40.28" />
                    <SPLIT distance="350" swimtime="00:04:18.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-04-21" firstname="Michał" gender="M" lastname="KRYSIAK" nation="POL" athleteid="100316">
              <RESULTS>
                <RESULT eventid="98798" points="437" reactiontime="+93" swimtime="00:00:27.54" resultid="100317" heatid="105141" lane="2" entrytime="00:00:26.50" />
                <RESULT eventid="98988" points="425" reactiontime="+89" swimtime="00:01:02.36" resultid="100318" heatid="105226" lane="2" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" status="DNS" swimtime="00:00:00.00" resultid="100319" heatid="105235" lane="4" entrytime="00:02:40.00" />
                <RESULT eventid="99170" points="428" reactiontime="+89" swimtime="00:00:29.76" resultid="100320" heatid="105274" lane="3" entrytime="00:00:29.00" />
                <RESULT eventid="99361" points="384" reactiontime="+88" swimtime="00:01:08.51" resultid="100321" heatid="105330" lane="3" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="335" reactiontime="+93" swimtime="00:05:16.66" resultid="100322" heatid="106061" lane="1" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                    <SPLIT distance="100" swimtime="00:01:12.46" />
                    <SPLIT distance="150" swimtime="00:01:53.50" />
                    <SPLIT distance="200" swimtime="00:02:34.61" />
                    <SPLIT distance="250" swimtime="00:03:17.43" />
                    <SPLIT distance="300" swimtime="00:04:00.81" />
                    <SPLIT distance="350" swimtime="00:04:39.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-03-20" firstname="Marcin" gender="M" lastname="ŁOGIN" nation="POL" swrid="4609021" athleteid="100323">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="100324" heatid="105133" lane="1" entrytime="00:00:30.23" />
                <RESULT eventid="98956" points="310" reactiontime="+126" swimtime="00:03:07.55" resultid="100325" heatid="105200" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.13" />
                    <SPLIT distance="100" swimtime="00:01:29.15" />
                    <SPLIT distance="150" swimtime="00:02:18.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="344" reactiontime="+110" swimtime="00:01:23.39" resultid="100326" heatid="105252" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="346" reactiontime="+92" swimtime="00:00:37.96" resultid="100327" heatid="105356" lane="9" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99250" points="410" reactiontime="+98" swimtime="00:01:54.16" resultid="100328" heatid="105311" lane="9" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.88" />
                    <SPLIT distance="100" swimtime="00:00:58.95" />
                    <SPLIT distance="150" swimtime="00:01:26.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100323" number="1" reactiontime="+98" />
                    <RELAYPOSITION athleteid="100283" number="2" />
                    <RELAYPOSITION athleteid="100294" number="3" reactiontime="+71" />
                    <RELAYPOSITION athleteid="100299" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99059" points="443" reactiontime="+82" swimtime="00:02:02.54" resultid="100329" heatid="105242" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                    <SPLIT distance="100" swimtime="00:01:07.55" />
                    <SPLIT distance="150" swimtime="00:01:36.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100294" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="100299" number="2" reactiontime="+70" />
                    <RELAYPOSITION athleteid="100316" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="100276" number="4" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="99250" points="414" reactiontime="+83" swimtime="00:01:53.84" resultid="100330" heatid="105311" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.45" />
                    <SPLIT distance="100" swimtime="00:00:59.12" />
                    <SPLIT distance="150" swimtime="00:01:27.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100316" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="100303" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="100290" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="100276" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99059" points="325" reactiontime="+91" swimtime="00:02:15.83" resultid="100331" heatid="105242" lane="0" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                    <SPLIT distance="100" swimtime="00:01:11.72" />
                    <SPLIT distance="150" swimtime="00:01:44.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100283" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="100323" number="2" reactiontime="+78" />
                    <RELAYPOSITION athleteid="100290" number="3" reactiontime="+67" />
                    <RELAYPOSITION athleteid="100303" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="105388" name="Szczecineckie Towarzystwo Pływackie Masters" shortname="Szczecineckie TP Mrs ">
          <ATHLETES>
            <ATHLETE birthdate="1933-02-19" firstname="Zbigniew" gender="M" lastname="LUDWICZAK" nation="POL" swrid="4992882" athleteid="100993">
              <RESULTS>
                <RESULT eventid="98798" points="69" swimtime="00:00:50.82" resultid="100994" heatid="105124" lane="0" entrytime="00:00:51.00" />
                <RESULT eventid="98924" points="59" reactiontime="+115" swimtime="00:01:01.53" resultid="100995" heatid="105181" lane="9" entrytime="00:00:57.00" />
                <RESULT eventid="98988" points="67" swimtime="00:01:55.03" resultid="100996" heatid="105213" lane="6" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="54" reactiontime="+137" swimtime="00:02:17.05" resultid="100997" heatid="105281" lane="2" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="65" swimtime="00:04:13.25" resultid="100998" heatid="105295" lane="2" entrytime="00:04:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.97" />
                    <SPLIT distance="100" swimtime="00:02:05.00" />
                    <SPLIT distance="150" swimtime="00:03:10.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="61" reactiontime="+114" swimtime="00:04:43.72" resultid="100999" heatid="105336" lane="1" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.58" />
                    <SPLIT distance="100" swimtime="00:02:19.27" />
                    <SPLIT distance="150" swimtime="00:03:33.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="73" swimtime="00:08:45.08" resultid="101000" heatid="106067" lane="4" entrytime="00:08:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.11" />
                    <SPLIT distance="100" swimtime="00:02:03.30" />
                    <SPLIT distance="150" swimtime="00:03:09.27" />
                    <SPLIT distance="200" swimtime="00:04:17.00" />
                    <SPLIT distance="250" swimtime="00:05:24.71" />
                    <SPLIT distance="300" swimtime="00:06:33.21" />
                    <SPLIT distance="350" swimtime="00:07:40.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="LTU" clubid="101429" name="TAKAS">
          <CONTACT city="Vilnius" email="abicka@takas.lt" internet="www.klubastakas.lt" name="Arlandas Antanas Juodeska" phone="+37068619471" street="Uzupio g. 3-4" zip="01200" />
          <ATHLETES>
            <ATHLETE birthdate="1951-06-04" firstname="Virginija" gender="F" lastname="VAISVILIENE" nation="LTU" swrid="4199518" athleteid="101432">
              <RESULTS>
                <RESULT eventid="98777" points="109" reactiontime="+115" swimtime="00:00:49.53" resultid="101433" heatid="105113" lane="4" entrytime="00:00:45.00" entrycourse="SCM" />
                <RESULT eventid="98814" points="114" reactiontime="+102" swimtime="00:04:20.10" resultid="101434" heatid="105144" lane="8" entrytime="00:04:18.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.04" />
                    <SPLIT distance="100" swimtime="00:02:08.97" />
                    <SPLIT distance="150" swimtime="00:03:22.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="120" reactiontime="+115" swimtime="00:04:41.49" resultid="101435" heatid="105191" lane="5" entrytime="00:04:18.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.74" />
                    <SPLIT distance="100" swimtime="00:02:18.58" />
                    <SPLIT distance="150" swimtime="00:03:29.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99004" points="88" reactiontime="+105" swimtime="00:04:33.78" resultid="101436" heatid="105229" lane="3" entrytime="00:04:21.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.01" />
                    <SPLIT distance="100" swimtime="00:02:07.89" />
                    <SPLIT distance="150" swimtime="00:03:22.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="85" swimtime="00:00:56.93" resultid="101437" heatid="105259" lane="8" entrytime="00:00:55.55" />
                <RESULT eventid="99202" points="97" reactiontime="+113" swimtime="00:04:05.19" resultid="101438" heatid="105289" lane="6" entrytime="00:04:09.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.77" />
                    <SPLIT distance="100" swimtime="00:02:00.07" />
                    <SPLIT distance="150" swimtime="00:03:04.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="85" reactiontime="+104" swimtime="00:02:07.04" resultid="101439" heatid="105321" lane="6" entrytime="00:01:59.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="102" reactiontime="+115" swimtime="00:01:02.97" resultid="101440" heatid="105344" lane="3" entrytime="00:00:56.25" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-09-25" firstname="Arturas" gender="M" lastname="TUOMAS" nation="LTU" swrid="4199517" athleteid="101441">
              <RESULTS>
                <RESULT eventid="98830" points="294" reactiontime="+78" swimtime="00:02:51.36" resultid="101442" heatid="105155" lane="9" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                    <SPLIT distance="100" swimtime="00:01:19.72" />
                    <SPLIT distance="150" swimtime="00:02:11.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="260" reactiontime="+85" swimtime="00:02:54.56" resultid="101443" heatid="105235" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.66" />
                    <SPLIT distance="100" swimtime="00:01:24.33" />
                    <SPLIT distance="150" swimtime="00:02:11.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" status="DNS" swimtime="00:00:00.00" resultid="101444" heatid="106052" lane="7" entrytime="00:05:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-02-06" firstname="Linas" gender="M" lastname="JOCIUS" nation="LTU" swrid="4267658" athleteid="101445">
              <RESULTS>
                <RESULT eventid="98798" points="241" reactiontime="+119" swimtime="00:00:33.56" resultid="101446" heatid="105128" lane="5" entrytime="00:00:33.50" />
                <RESULT eventid="98988" points="214" reactiontime="+90" swimtime="00:01:18.35" resultid="101447" heatid="105217" lane="8" entrytime="00:01:14.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-03-24" firstname="Ruta" gender="F" lastname="RIMKEVICIENE" nation="LTU" swrid="4595564" athleteid="101448">
              <RESULTS>
                <RESULT eventid="99202" points="293" reactiontime="+87" swimtime="00:02:50.03" resultid="101449" heatid="105292" lane="9" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.52" />
                    <SPLIT distance="100" swimtime="00:01:21.96" />
                    <SPLIT distance="150" swimtime="00:02:06.66" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="04" eventid="99344" reactiontime="+78" status="DSQ" swimtime="00:00:00.00" resultid="101450" heatid="105322" lane="6" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-02-12" firstname="Irena" gender="F" lastname="JOKUBAITIENE" nation="LTU" swrid="4270248" athleteid="101451">
              <RESULTS>
                <RESULT eventid="98777" points="111" reactiontime="+112" swimtime="00:00:49.36" resultid="101452" heatid="105113" lane="7" entrytime="00:00:50.00" />
                <RESULT eventid="98940" points="157" reactiontime="+106" swimtime="00:04:17.76" resultid="101453" heatid="105191" lane="6" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.21" />
                    <SPLIT distance="100" swimtime="00:02:03.46" />
                    <SPLIT distance="150" swimtime="00:03:10.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="144" reactiontime="+111" swimtime="00:02:02.76" resultid="101454" heatid="105244" lane="2" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="142" reactiontime="+100" swimtime="00:00:56.50" resultid="101455" heatid="105345" lane="9" entrytime="00:00:54.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-10-18" firstname="Ramune" gender="F" lastname="IVANAUSKAITE" nation="LTU" swrid="4750033" athleteid="101456">
              <RESULTS>
                <RESULT eventid="98814" points="272" reactiontime="+67" swimtime="00:03:14.61" resultid="101457" heatid="105146" lane="8" entrytime="00:03:06.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.96" />
                    <SPLIT distance="100" swimtime="00:01:32.45" />
                    <SPLIT distance="150" swimtime="00:02:29.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="268" reactiontime="+110" swimtime="00:00:41.95" resultid="101458" heatid="105176" lane="0" entrytime="00:00:39.70" />
                <RESULT eventid="98940" points="273" reactiontime="+80" swimtime="00:03:34.40" resultid="101459" heatid="105193" lane="6" entrytime="00:03:27.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.17" />
                    <SPLIT distance="100" swimtime="00:01:45.13" />
                    <SPLIT distance="150" swimtime="00:02:40.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="266" reactiontime="+92" swimtime="00:01:39.95" resultid="101460" heatid="105246" lane="3" entrytime="00:01:33.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="254" reactiontime="+91" swimtime="00:01:31.77" resultid="101461" heatid="105279" lane="7" entrytime="00:01:27.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="277" reactiontime="+100" swimtime="00:02:53.12" resultid="101462" heatid="105292" lane="2" entrytime="00:02:45.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.00" />
                    <SPLIT distance="100" swimtime="00:01:23.90" />
                    <SPLIT distance="150" swimtime="00:02:09.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="262" reactiontime="+92" swimtime="00:03:13.70" resultid="101463" heatid="105334" lane="0" entrytime="00:03:06.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.05" />
                    <SPLIT distance="100" swimtime="00:01:34.12" />
                    <SPLIT distance="150" swimtime="00:02:23.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="272" swimtime="00:06:08.67" resultid="101464" heatid="106055" lane="7" entrytime="00:05:51.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.35" />
                    <SPLIT distance="100" swimtime="00:01:25.12" />
                    <SPLIT distance="150" swimtime="00:02:11.41" />
                    <SPLIT distance="200" swimtime="00:02:58.94" />
                    <SPLIT distance="250" swimtime="00:03:46.86" />
                    <SPLIT distance="300" swimtime="00:04:35.13" />
                    <SPLIT distance="350" swimtime="00:05:23.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-08-22" firstname="Arvydas" gender="M" lastname="BURINSKAS" nation="LTU" swrid="4199513" athleteid="101465">
              <RESULTS>
                <RESULT eventid="99020" points="268" reactiontime="+77" swimtime="00:02:52.84" resultid="101466" heatid="105235" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.51" />
                    <SPLIT distance="100" swimtime="00:01:22.70" />
                    <SPLIT distance="150" swimtime="00:02:07.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="390" reactiontime="+80" swimtime="00:00:30.69" resultid="101467" heatid="105273" lane="0" entrytime="00:00:30.50" />
                <RESULT eventid="99361" points="300" reactiontime="+77" swimtime="00:01:14.38" resultid="101468" heatid="105329" lane="6" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1938-08-27" firstname="Aldona" gender="F" lastname="VILKIENE" nation="LTU" swrid="4477505" athleteid="101469">
              <RESULTS>
                <RESULT eventid="99202" points="128" reactiontime="+109" swimtime="00:03:44.08" resultid="101470" heatid="105289" lane="3" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.59" />
                    <SPLIT distance="100" swimtime="00:01:46.63" />
                    <SPLIT distance="150" swimtime="00:02:46.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="137" reactiontime="+101" swimtime="00:07:42.83" resultid="101471" heatid="106057" lane="3" entrytime="00:07:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.61" />
                    <SPLIT distance="100" swimtime="00:01:50.12" />
                    <SPLIT distance="150" swimtime="00:02:49.15" />
                    <SPLIT distance="200" swimtime="00:03:48.29" />
                    <SPLIT distance="250" swimtime="00:04:46.71" />
                    <SPLIT distance="300" swimtime="00:05:45.30" />
                    <SPLIT distance="350" swimtime="00:06:43.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-06-18" firstname="Linas" gender="M" lastname="KERSEVICIUS" nation="LTU" swrid="4199514" athleteid="101472">
              <RESULTS>
                <RESULT eventid="98830" points="368" reactiontime="+94" swimtime="00:02:39.03" resultid="101473" heatid="105155" lane="1" entrytime="00:02:40.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                    <SPLIT distance="100" swimtime="00:01:13.70" />
                    <SPLIT distance="150" swimtime="00:02:00.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="420" reactiontime="+81" swimtime="00:00:32.08" resultid="101474" heatid="105188" lane="4" entrytime="00:00:32.59" />
                <RESULT eventid="99186" points="427" reactiontime="+70" swimtime="00:01:08.94" resultid="101475" heatid="105287" lane="8" entrytime="00:01:10.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="412" reactiontime="+81" swimtime="00:02:30.31" resultid="101476" heatid="105342" lane="8" entrytime="00:02:33.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                    <SPLIT distance="100" swimtime="00:01:12.03" />
                    <SPLIT distance="150" swimtime="00:01:51.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-12-26" firstname="Arlandas Antanas" gender="M" lastname="JUODESKA" nation="LTU" athleteid="101477">
              <RESULTS>
                <RESULT eventid="98798" points="346" reactiontime="+84" swimtime="00:00:29.78" resultid="101478" heatid="105136" lane="4" entrytime="00:00:28.70" />
                <RESULT eventid="98924" points="358" reactiontime="+70" swimtime="00:00:33.83" resultid="101479" heatid="105187" lane="5" entrytime="00:00:33.40" />
                <RESULT eventid="99091" points="311" reactiontime="+77" swimtime="00:01:26.22" resultid="101480" heatid="105255" lane="9" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="289" reactiontime="+78" swimtime="00:01:18.54" resultid="101481" heatid="105285" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="359" reactiontime="+87" swimtime="00:00:37.52" resultid="101482" heatid="105358" lane="2" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-06-08" firstname="Viktoras" gender="M" lastname="SNIESKA" nation="LTU" swrid="4845234" athleteid="101483">
              <RESULTS>
                <RESULT eventid="98798" points="244" reactiontime="+97" swimtime="00:00:33.43" resultid="101484" heatid="105129" lane="0" entrytime="00:00:33.03" />
                <RESULT eventid="98891" points="171" swimtime="00:26:08.93" resultid="101485" heatid="105424" lane="5" entrytime="00:26:40.10" />
                <RESULT eventid="98924" points="189" reactiontime="+88" swimtime="00:00:41.89" resultid="101486" heatid="105184" lane="3" entrytime="00:00:40.23" />
                <RESULT eventid="98988" points="217" reactiontime="+112" swimtime="00:01:18.05" resultid="101487" heatid="105217" lane="1" entrytime="00:01:14.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="172" reactiontime="+91" swimtime="00:01:33.32" resultid="101488" heatid="105283" lane="2" entrytime="00:01:31.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="152" swimtime="00:07:36.61" resultid="101489" heatid="106049" lane="8" entrytime="00:07:41.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.23" />
                    <SPLIT distance="100" swimtime="00:01:59.34" />
                    <SPLIT distance="150" swimtime="00:02:54.38" />
                    <SPLIT distance="200" swimtime="00:03:50.53" />
                    <SPLIT distance="250" swimtime="00:04:54.58" />
                    <SPLIT distance="300" swimtime="00:05:58.00" />
                    <SPLIT distance="350" swimtime="00:06:47.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="155" reactiontime="+104" swimtime="00:03:27.93" resultid="101490" heatid="105343" lane="2" entrytime="00:02:21.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.08" />
                    <SPLIT distance="100" swimtime="00:01:38.75" />
                    <SPLIT distance="150" swimtime="00:02:33.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="167" reactiontime="+97" swimtime="00:06:39.01" resultid="101491" heatid="106064" lane="9" entrytime="00:06:21.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.83" />
                    <SPLIT distance="100" swimtime="00:01:32.18" />
                    <SPLIT distance="150" swimtime="00:02:22.08" />
                    <SPLIT distance="200" swimtime="00:03:13.09" />
                    <SPLIT distance="250" swimtime="00:04:04.43" />
                    <SPLIT distance="300" swimtime="00:04:56.96" />
                    <SPLIT distance="350" swimtime="00:05:49.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-04-12" firstname="Aleksandra" gender="F" lastname="YLIENE" nation="LTU" swrid="4182530" athleteid="101492">
              <RESULTS>
                <RESULT eventid="98777" points="151" reactiontime="+102" swimtime="00:00:44.49" resultid="101493" heatid="105114" lane="8" entrytime="00:00:43.16" entrycourse="LCM" />
                <RESULT eventid="98907" points="151" reactiontime="+89" swimtime="00:00:50.74" resultid="101494" heatid="105173" lane="4" entrytime="00:00:49.85" />
                <RESULT eventid="98972" points="137" reactiontime="+119" swimtime="00:01:40.82" resultid="101495" heatid="105206" lane="1" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="110" reactiontime="+97" swimtime="00:02:01.23" resultid="101496" heatid="105277" lane="3" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="101" reactiontime="+100" swimtime="00:04:25.54" resultid="101497" heatid="105332" lane="2" entrytime="00:04:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.76" />
                    <SPLIT distance="100" swimtime="00:02:11.88" />
                    <SPLIT distance="150" swimtime="00:03:22.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-21" firstname="Rimvydas" gender="M" lastname="ANIULIS" nation="LTU" athleteid="101498">
              <RESULTS>
                <RESULT eventid="98798" points="377" reactiontime="+87" swimtime="00:00:28.94" resultid="101499" heatid="105126" lane="8" entrytime="00:00:37.00" />
                <RESULT eventid="99170" points="387" reactiontime="+97" swimtime="00:00:30.77" resultid="101500" heatid="105267" lane="0" entrytime="00:00:41.00" />
                <RESULT eventid="99425" points="385" reactiontime="+100" swimtime="00:00:36.66" resultid="101501" heatid="105353" lane="1" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="102632" name="TKKF Koszalin Masters">
          <CONTACT city="Koszalin" email="jakubkielar3@gmail.com" name="Kielar" phone="693193137" street="ul Holenderska 6" zip="75-430" />
          <ATHLETES>
            <ATHLETE birthdate="1951-02-03" firstname="Andrzej" gender="M" lastname="MICHAŁKOWSKI" nation="POL" swrid="4754754" athleteid="102633">
              <RESULTS>
                <RESULT eventid="98798" points="152" reactiontime="+113" swimtime="00:00:39.13" resultid="102634" heatid="105125" lane="5" entrytime="00:00:38.50" />
                <RESULT eventid="98830" points="116" reactiontime="+131" swimtime="00:03:53.43" resultid="102635" heatid="105149" lane="4" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.54" />
                    <SPLIT distance="100" swimtime="00:01:57.31" />
                    <SPLIT distance="150" swimtime="00:02:58.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="161" swimtime="00:03:53.30" resultid="102636" heatid="105198" lane="7" entrytime="00:03:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.26" />
                    <SPLIT distance="100" swimtime="00:01:49.80" />
                    <SPLIT distance="150" swimtime="00:02:52.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="108" reactiontime="+115" swimtime="00:01:38.48" resultid="102637" heatid="105214" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="195" reactiontime="+118" swimtime="00:01:40.76" resultid="102638" heatid="105250" lane="4" entrytime="00:01:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="90" reactiontime="+123" swimtime="00:03:47.17" resultid="102639" heatid="105295" lane="5" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.40" />
                    <SPLIT distance="100" swimtime="00:01:45.59" />
                    <SPLIT distance="150" swimtime="00:02:48.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="258" reactiontime="+109" swimtime="00:00:41.86" resultid="102640" heatid="105355" lane="5" entrytime="00:00:41.30" />
                <RESULT eventid="99473" points="86" reactiontime="+97" swimtime="00:08:17.86" resultid="102641" heatid="106066" lane="8" entrytime="00:07:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.70" />
                    <SPLIT distance="100" swimtime="00:01:48.84" />
                    <SPLIT distance="150" swimtime="00:02:53.40" />
                    <SPLIT distance="200" swimtime="00:03:56.84" />
                    <SPLIT distance="250" swimtime="00:05:01.90" />
                    <SPLIT distance="300" swimtime="00:06:07.80" />
                    <SPLIT distance="350" swimtime="00:07:14.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="100400" name="TP Masters Opole">
          <CONTACT city="OPOLE" name="KRASNODĘBSKI" />
          <ATHLETES>
            <ATHLETE birthdate="1937-01-01" firstname="Tadeusz" gender="M" lastname="WITKOWSKI" nation="POL" swrid="4187082" athleteid="100401">
              <RESULTS>
                <RESULT eventid="98798" points="190" reactiontime="+121" swimtime="00:00:36.34" resultid="100402" heatid="105126" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="98830" points="61" reactiontime="+113" swimtime="00:04:48.20" resultid="100403" heatid="105149" lane="8" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.89" />
                    <SPLIT distance="100" swimtime="00:02:26.47" />
                    <SPLIT distance="150" swimtime="00:03:55.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="105" reactiontime="+99" swimtime="00:00:50.88" resultid="100404" heatid="105182" lane="2" entrytime="00:00:48.50" />
                <RESULT eventid="98988" points="140" reactiontime="+117" swimtime="00:01:30.20" resultid="100405" heatid="105214" lane="6" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="92" reactiontime="+96" swimtime="00:01:54.99" resultid="100406" heatid="105281" lane="5" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="97" reactiontime="+127" swimtime="00:03:41.42" resultid="100407" heatid="105296" lane="2" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.47" />
                    <SPLIT distance="100" swimtime="00:01:46.43" />
                    <SPLIT distance="150" swimtime="00:02:45.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="90" reactiontime="+85" swimtime="00:04:09.35" resultid="100408" heatid="105336" lane="6" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.43" />
                    <SPLIT distance="100" swimtime="00:02:03.48" />
                    <SPLIT distance="150" swimtime="00:03:08.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="110" reactiontime="+110" swimtime="00:00:55.53" resultid="100409" heatid="105351" lane="6" entrytime="00:00:51.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-02-23" firstname="Grzegorz" gender="M" lastname="RADOMSKI" nation="POL" swrid="4061108" athleteid="101007">
              <RESULTS>
                <RESULT eventid="98830" points="572" reactiontime="+80" swimtime="00:02:17.33" resultid="101008" heatid="105158" lane="6" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.28" />
                    <SPLIT distance="100" swimtime="00:01:04.73" />
                    <SPLIT distance="150" swimtime="00:01:43.51" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters, Rekord Polski Masters" eventid="98891" points="466" swimtime="00:18:42.89" resultid="101009" heatid="105420" lane="6" entrytime="00:19:30.00" />
                <RESULT comment="Rekord Polski Masters" eventid="99218" points="521" reactiontime="+83" swimtime="00:02:06.69" resultid="101010" heatid="105304" lane="3" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.27" />
                    <SPLIT distance="100" swimtime="00:00:59.77" />
                    <SPLIT distance="150" swimtime="00:01:32.82" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99282" points="532" reactiontime="+83" swimtime="00:05:00.77" resultid="101011" heatid="106053" lane="6" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                    <SPLIT distance="100" swimtime="00:01:09.66" />
                    <SPLIT distance="150" swimtime="00:01:47.88" />
                    <SPLIT distance="200" swimtime="00:02:26.39" />
                    <SPLIT distance="250" swimtime="00:03:07.18" />
                    <SPLIT distance="300" swimtime="00:03:49.50" />
                    <SPLIT distance="350" swimtime="00:04:25.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="493" reactiontime="+69" swimtime="00:02:21.63" resultid="101012" heatid="105343" lane="8" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                    <SPLIT distance="100" swimtime="00:01:08.08" />
                    <SPLIT distance="150" swimtime="00:01:45.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="527" reactiontime="+89" swimtime="00:04:32.29" resultid="101013" heatid="106060" lane="1" entrytime="00:04:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.67" />
                    <SPLIT distance="100" swimtime="00:01:02.74" />
                    <SPLIT distance="150" swimtime="00:01:36.82" />
                    <SPLIT distance="200" swimtime="00:02:11.97" />
                    <SPLIT distance="250" swimtime="00:02:47.11" />
                    <SPLIT distance="300" swimtime="00:03:22.37" />
                    <SPLIT distance="350" swimtime="00:03:57.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="MAŁ" clubid="100839" name="TS Masters Wisła Kraków">
          <CONTACT email="wislaplywanie@gmail.com" internet="http://www.wislaplywanie.pl/sekcja-masters/" name="Wolski Wojciech" phone="791126323" />
          <ATHLETES>
            <ATHLETE birthdate="1966-03-28" firstname="Wojciech" gender="M" lastname="WOLSKI" nation="POL" swrid="4754645" athleteid="100856">
              <RESULTS>
                <RESULT eventid="98798" points="247" reactiontime="+99" swimtime="00:00:33.29" resultid="100857" heatid="105130" lane="0" entrytime="00:00:32.25" />
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="100858" heatid="105152" lane="1" entrytime="00:03:05.69" />
                <RESULT eventid="98956" points="243" reactiontime="+95" swimtime="00:03:23.32" resultid="100859" heatid="105200" lane="6" entrytime="00:03:15.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.96" />
                    <SPLIT distance="100" swimtime="00:01:33.39" />
                    <SPLIT distance="150" swimtime="00:02:28.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="256" reactiontime="+88" swimtime="00:01:32.05" resultid="100860" heatid="105253" lane="9" entrytime="00:01:29.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="100861" heatid="105268" lane="1" entrytime="00:00:36.67" />
                <RESULT eventid="99282" points="186" reactiontime="+111" swimtime="00:07:07.12" resultid="100862" heatid="106050" lane="7" entrytime="00:06:52.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                    <SPLIT distance="100" swimtime="00:01:33.49" />
                    <SPLIT distance="150" swimtime="00:02:35.54" />
                    <SPLIT distance="200" swimtime="00:03:37.36" />
                    <SPLIT distance="250" swimtime="00:04:35.57" />
                    <SPLIT distance="300" swimtime="00:05:31.34" />
                    <SPLIT distance="350" swimtime="00:06:17.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="171" reactiontime="+100" swimtime="00:01:29.59" resultid="100863" heatid="105327" lane="7" entrytime="00:01:29.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="290" reactiontime="+94" swimtime="00:00:40.28" resultid="100864" heatid="105357" lane="8" entrytime="00:00:39.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-09-22" firstname="Mateusz" gender="M" lastname="DYBEK" nation="POL" swrid="4992906" athleteid="100865">
              <RESULTS>
                <RESULT eventid="98891" points="329" swimtime="00:21:00.45" resultid="100866" heatid="105422" lane="5" entrytime="00:22:20.50" entrycourse="LCM" />
                <RESULT eventid="98988" points="490" reactiontime="+88" swimtime="00:00:59.47" resultid="100867" heatid="105226" lane="3" entrytime="00:00:58.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="403" reactiontime="+84" swimtime="00:02:17.98" resultid="100868" heatid="105303" lane="3" entrytime="00:02:14.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.52" />
                    <SPLIT distance="100" swimtime="00:01:04.82" />
                    <SPLIT distance="150" swimtime="00:01:41.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="339" reactiontime="+89" swimtime="00:05:15.54" resultid="100869" heatid="106062" lane="3" entrytime="00:05:08.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                    <SPLIT distance="100" swimtime="00:01:13.81" />
                    <SPLIT distance="150" swimtime="00:01:53.31" />
                    <SPLIT distance="200" swimtime="00:02:33.05" />
                    <SPLIT distance="250" swimtime="00:03:13.06" />
                    <SPLIT distance="300" swimtime="00:03:54.22" />
                    <SPLIT distance="350" swimtime="00:04:35.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-05-28" firstname="Marta" gender="F" lastname="WOLSKA" nation="POL" swrid="4754644" athleteid="100870">
              <RESULTS>
                <RESULT eventid="98777" points="109" reactiontime="+168" swimtime="00:00:49.58" resultid="100871" heatid="105113" lane="1" entrytime="00:00:50.62" entrycourse="SCM" />
                <RESULT eventid="98907" points="112" reactiontime="+77" swimtime="00:00:56.09" resultid="100872" heatid="105173" lane="9" entrytime="00:00:56.94" />
                <RESULT eventid="98940" points="118" reactiontime="+155" swimtime="00:04:43.35" resultid="100873" heatid="105191" lane="2" entrytime="00:04:52.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.31" />
                    <SPLIT distance="100" swimtime="00:02:16.15" />
                    <SPLIT distance="150" swimtime="00:03:30.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="112" reactiontime="+143" swimtime="00:02:13.44" resultid="100874" heatid="105244" lane="0" entrytime="00:02:16.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="118" swimtime="00:01:58.36" resultid="100875" heatid="105277" lane="6" entrytime="00:02:09.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="110" reactiontime="+80" swimtime="00:04:18.83" resultid="100876" heatid="105332" lane="7" entrytime="00:04:38.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.15" />
                    <SPLIT distance="100" swimtime="00:02:06.81" />
                    <SPLIT distance="150" swimtime="00:03:14.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="124" reactiontime="+141" swimtime="00:00:58.97" resultid="100877" heatid="105344" lane="6" entrytime="00:00:58.58" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-04" firstname="Małgorzata" gender="F" lastname="SKALSKA" nation="POL" swrid="5023973" athleteid="100878">
              <RESULTS>
                <RESULT eventid="98777" points="194" reactiontime="+104" swimtime="00:00:40.94" resultid="100879" heatid="105114" lane="4" entrytime="00:00:40.03" />
                <RESULT eventid="98940" points="232" reactiontime="+110" swimtime="00:03:46.16" resultid="100880" heatid="105192" lane="6" entrytime="00:03:50.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.10" />
                    <SPLIT distance="100" swimtime="00:01:52.76" />
                    <SPLIT distance="150" swimtime="00:02:51.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" status="DNS" swimtime="00:00:00.00" resultid="100881" heatid="105206" lane="4" entrytime="00:01:30.74" />
                <RESULT eventid="99089" points="242" reactiontime="+98" swimtime="00:01:43.13" resultid="100882" heatid="105245" lane="6" entrytime="00:01:43.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="184" reactiontime="+103" swimtime="00:03:18.62" resultid="100883" heatid="105290" lane="5" entrytime="00:03:17.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.06" />
                    <SPLIT distance="100" swimtime="00:01:36.72" />
                    <SPLIT distance="150" swimtime="00:02:29.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="259" reactiontime="+99" swimtime="00:00:46.24" resultid="100884" heatid="105346" lane="1" entrytime="00:00:48.05" />
                <RESULT eventid="99457" points="175" reactiontime="+112" swimtime="00:07:07.30" resultid="100885" heatid="106057" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.32" />
                    <SPLIT distance="100" swimtime="00:01:40.85" />
                    <SPLIT distance="150" swimtime="00:02:35.77" />
                    <SPLIT distance="200" swimtime="00:03:30.82" />
                    <SPLIT distance="250" swimtime="00:04:26.28" />
                    <SPLIT distance="300" swimtime="00:05:21.86" />
                    <SPLIT distance="350" swimtime="00:06:16.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-03-19" firstname="Paulina" gender="F" lastname="PALKA" nation="POL" swrid="4072437" athleteid="100886">
              <RESULTS>
                <RESULT eventid="98814" points="353" reactiontime="+62" swimtime="00:02:58.48" resultid="100887" heatid="105147" lane="8" entrytime="00:02:52.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.16" />
                    <SPLIT distance="100" swimtime="00:01:23.04" />
                    <SPLIT distance="150" swimtime="00:02:16.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="433" reactiontime="+70" swimtime="00:00:35.76" resultid="100888" heatid="105178" lane="0" entrytime="00:00:35.20" entrycourse="LCM" />
                <RESULT eventid="99314" points="436" reactiontime="+60" swimtime="00:01:16.59" resultid="100889" heatid="105280" lane="6" entrytime="00:01:14.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="388" reactiontime="+70" swimtime="00:02:50.03" resultid="100890" heatid="105334" lane="4" entrytime="00:02:44.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                    <SPLIT distance="100" swimtime="00:01:22.50" />
                    <SPLIT distance="150" swimtime="00:02:06.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-09-10" firstname="Janusz" gender="M" lastname="MROZIK" nation="POL" athleteid="100891">
              <RESULTS>
                <RESULT eventid="98956" points="56" swimtime="00:05:31.40" resultid="100892" heatid="105196" lane="2" />
                <RESULT eventid="99091" points="55" reactiontime="+122" swimtime="00:02:33.16" resultid="100893" heatid="105248" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="48" swimtime="00:02:22.03" resultid="100894" heatid="105283" lane="7" />
                <RESULT eventid="99393" points="48" reactiontime="+129" swimtime="00:05:06.23" resultid="100895" heatid="105335" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:31.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="OLPOZ" nation="POL" region="WIE" clubid="102531" name="TS Olimpia Poznań">
          <CONTACT name="Pietraszewski" phone="501 648 415" />
          <ATHLETES>
            <ATHLETE birthdate="1950-01-01" firstname="Maria" gender="F" lastname="ŁUTOWICZ" nation="POL" swrid="4188428" athleteid="102532">
              <RESULTS>
                <RESULT eventid="98777" points="236" reactiontime="+93" swimtime="00:00:38.37" resultid="102533" heatid="105115" lane="3" entrytime="00:00:38.00" entrycourse="LCM" />
                <RESULT eventid="98907" points="164" swimtime="00:00:49.34" resultid="102534" heatid="105173" lane="1" entrytime="00:00:52.00" />
                <RESULT eventid="98972" points="204" reactiontime="+103" swimtime="00:01:28.31" resultid="102535" heatid="105206" lane="2" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="138" reactiontime="+92" swimtime="00:00:48.43" resultid="102536" heatid="105259" lane="3" entrytime="00:00:49.00" />
                <RESULT eventid="99202" points="173" reactiontime="+100" swimtime="00:03:22.41" resultid="102537" heatid="105290" lane="1" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.15" />
                    <SPLIT distance="100" swimtime="00:01:40.94" />
                    <SPLIT distance="150" swimtime="00:02:33.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="178" reactiontime="+103" swimtime="00:00:52.35" resultid="102538" heatid="105345" lane="5" entrytime="00:00:51.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Grażyna" gender="F" lastname="CABAJ- DRELA" nation="POL" swrid="4754706" athleteid="102539">
              <RESULTS>
                <RESULT eventid="98777" points="328" reactiontime="+80" swimtime="00:00:34.38" resultid="102540" heatid="105117" lane="7" entrytime="00:00:35.00" />
                <RESULT comment="Rekord Polski Masters, Rekord Polski " eventid="98814" points="299" reactiontime="+93" swimtime="00:03:08.60" resultid="102541" heatid="105145" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.08" />
                    <SPLIT distance="100" swimtime="00:01:29.61" />
                    <SPLIT distance="150" swimtime="00:02:23.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="279" reactiontime="+86" swimtime="00:00:41.38" resultid="102542" heatid="105175" lane="5" entrytime="00:00:41.00" />
                <RESULT eventid="98940" points="306" reactiontime="+92" swimtime="00:03:26.42" resultid="102543" heatid="105193" lane="3" entrytime="00:03:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.60" />
                    <SPLIT distance="100" swimtime="00:01:39.57" />
                    <SPLIT distance="150" swimtime="00:02:33.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="321" reactiontime="+81" swimtime="00:01:33.91" resultid="102544" heatid="105246" lane="7" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="230" reactiontime="+88" swimtime="00:00:40.87" resultid="102545" heatid="105259" lane="5" entrytime="00:00:45.00" />
                <RESULT comment="Rekord Polski Masters" eventid="99409" points="322" reactiontime="+85" swimtime="00:00:42.99" resultid="102546" heatid="105347" lane="8" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-01-01" firstname="Joanna" gender="F" lastname="PUCHALSKA" nation="POL" swrid="4435044" athleteid="102547">
              <RESULTS>
                <RESULT eventid="98814" status="DNS" swimtime="00:00:00.00" resultid="102548" heatid="105147" lane="1" entrytime="00:02:52.00" />
                <RESULT eventid="98940" status="DNS" swimtime="00:00:00.00" resultid="102549" heatid="105194" lane="2" entrytime="00:03:12.00" />
                <RESULT eventid="99089" status="DNS" swimtime="00:00:00.00" resultid="102550" heatid="105247" lane="0" entrytime="00:01:29.00" />
                <RESULT eventid="99154" status="DNS" swimtime="00:00:00.00" resultid="102551" heatid="105262" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="99344" status="DNS" swimtime="00:00:00.00" resultid="102552" heatid="105323" lane="1" entrytime="00:01:17.00" />
                <RESULT eventid="99457" status="WDR" swimtime="00:00:00.00" resultid="102553" entrytime="00:05:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-01-01" firstname="Jacek" gender="M" lastname="LESIŃSKI" nation="POL" swrid="4188190" athleteid="102554">
              <RESULTS>
                <RESULT eventid="98798" points="169" reactiontime="+106" swimtime="00:00:37.78" resultid="102555" heatid="105123" lane="2" />
                <RESULT eventid="98830" points="130" reactiontime="+112" swimtime="00:03:44.59" resultid="102556" heatid="105150" lane="1" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.97" />
                    <SPLIT distance="100" swimtime="00:01:49.68" />
                    <SPLIT distance="150" swimtime="00:02:54.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="159" reactiontime="+84" swimtime="00:00:44.37" resultid="102557" heatid="105183" lane="8" entrytime="00:00:45.00" />
                <RESULT eventid="98988" points="150" reactiontime="+114" swimtime="00:01:28.14" resultid="102558" heatid="105214" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="127" reactiontime="+81" swimtime="00:01:43.31" resultid="102559" heatid="105282" lane="5" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="113" reactiontime="+92" swimtime="00:03:51.34" resultid="102560" heatid="105337" lane="4" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.59" />
                    <SPLIT distance="100" swimtime="00:01:50.47" />
                    <SPLIT distance="150" swimtime="00:02:51.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Jerzy" gender="M" lastname="BORYSKI" nation="POL" swrid="4754708" athleteid="102561">
              <RESULTS>
                <RESULT eventid="98798" points="161" reactiontime="+115" swimtime="00:00:38.41" resultid="102562" heatid="105126" lane="2" entrytime="00:00:36.50" />
                <RESULT eventid="98924" points="158" reactiontime="+97" swimtime="00:00:44.41" resultid="102563" heatid="105183" lane="1" entrytime="00:00:43.50" />
                <RESULT eventid="99186" points="139" reactiontime="+85" swimtime="00:01:40.17" resultid="102564" heatid="105283" lane="8" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="115" reactiontime="+86" swimtime="00:03:49.93" resultid="102565" heatid="105338" lane="9" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.63" />
                    <SPLIT distance="100" swimtime="00:01:54.47" />
                    <SPLIT distance="150" swimtime="00:02:55.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="102566" entrytime="00:07:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Zbigniew" gender="M" lastname="PIETRASZEWSKI" nation="POL" swrid="4187282" athleteid="102567">
              <RESULTS>
                <RESULT eventid="98830" points="206" reactiontime="+91" swimtime="00:03:12.98" resultid="102568" heatid="105152" lane="8" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.22" />
                    <SPLIT distance="100" swimtime="00:01:36.03" />
                    <SPLIT distance="150" swimtime="00:02:29.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="177" reactiontime="+93" swimtime="00:00:42.81" resultid="102569" heatid="105184" lane="2" entrytime="00:00:41.00" />
                <RESULT eventid="99186" points="181" reactiontime="+86" swimtime="00:01:31.68" resultid="102570" heatid="105283" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="202" reactiontime="+105" swimtime="00:06:55.17" resultid="102571" heatid="106050" lane="5" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.00" />
                    <SPLIT distance="100" swimtime="00:01:47.19" />
                    <SPLIT distance="150" swimtime="00:02:39.43" />
                    <SPLIT distance="200" swimtime="00:03:30.87" />
                    <SPLIT distance="250" swimtime="00:04:26.37" />
                    <SPLIT distance="300" swimtime="00:05:22.31" />
                    <SPLIT distance="350" swimtime="00:06:09.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="191" reactiontime="+94" swimtime="00:03:14.17" resultid="102572" heatid="105339" lane="0" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.31" />
                    <SPLIT distance="100" swimtime="00:01:35.60" />
                    <SPLIT distance="150" swimtime="00:02:25.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Sławomir" gender="M" lastname="CYBERTOWICZ" nation="POL" swrid="4269915" athleteid="102573">
              <RESULTS>
                <RESULT eventid="98956" status="DNS" swimtime="00:00:00.00" resultid="102574" heatid="105202" lane="1" entrytime="00:03:05.00" />
                <RESULT eventid="99091" points="351" reactiontime="+82" swimtime="00:01:22.87" resultid="102575" heatid="105254" lane="3" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="291" reactiontime="+82" swimtime="00:02:33.76" resultid="102576" heatid="105300" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.87" />
                    <SPLIT distance="100" swimtime="00:01:13.77" />
                    <SPLIT distance="150" swimtime="00:01:54.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="102577" heatid="105357" lane="4" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-01" firstname="Bartłomiej" gender="M" lastname="ZADOROŻNY" nation="POL" swrid="4920304" athleteid="102578">
              <RESULTS>
                <RESULT eventid="98798" points="381" reactiontime="+70" swimtime="00:00:28.82" resultid="102579" heatid="105139" lane="9" entrytime="00:00:27.66" />
                <RESULT eventid="98924" points="270" reactiontime="+81" swimtime="00:00:37.16" resultid="102580" heatid="105186" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="98988" points="390" reactiontime="+79" swimtime="00:01:04.17" resultid="102581" heatid="105224" lane="5" entrytime="00:01:01.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="371" reactiontime="+81" swimtime="00:01:21.31" resultid="102582" heatid="105256" lane="5" entrytime="00:01:18.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="328" reactiontime="+82" swimtime="00:00:32.51" resultid="102583" heatid="105269" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="99425" points="416" reactiontime="+89" swimtime="00:00:35.71" resultid="102584" heatid="105360" lane="2" entrytime="00:00:34.95" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" status="DNS" swimtime="00:00:00.00" resultid="102585" heatid="105160" lane="4" entrytime="00:02:06.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102573" number="1" />
                    <RELAYPOSITION athleteid="102539" number="2" />
                    <RELAYPOSITION athleteid="102547" number="3" />
                    <RELAYPOSITION athleteid="102578" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="99441" points="220" reactiontime="+90" swimtime="00:02:34.61" resultid="102586" heatid="105364" lane="8" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.38" />
                    <SPLIT distance="100" swimtime="00:01:23.24" />
                    <SPLIT distance="150" swimtime="00:01:55.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102539" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="102567" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="102578" number="3" reactiontime="+72" />
                    <RELAYPOSITION athleteid="102532" number="4" reactiontime="+89" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="LTU" clubid="105041" name="Torpedos">
          <CONTACT city="Marijampole" email="vilmantasenator@gmail.com" name="Aldona Mazetiene" phone="+37068746068" street="Jukneviciaus 78-10" zip="68198" />
          <ATHLETES>
            <ATHLETE birthdate="1964-07-31" firstname="Vilmantas" gender="M" lastname="KRASAUSKAS" nation="LTU" athleteid="105042">
              <RESULTS>
                <RESULT eventid="98798" points="350" reactiontime="+83" swimtime="00:00:29.67" resultid="105043" heatid="105134" lane="5" entrytime="00:00:29.94" entrycourse="LCM" />
                <RESULT eventid="98891" points="334" swimtime="00:20:55.25" resultid="105044" heatid="105421" lane="5" entrytime="00:20:15.08" entrycourse="LCM" />
                <RESULT eventid="98988" points="357" reactiontime="+92" swimtime="00:01:06.08" resultid="105045" heatid="105222" lane="3" entrytime="00:01:04.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="373" reactiontime="+87" swimtime="00:02:21.67" resultid="105046" heatid="105301" lane="4" entrytime="00:02:20.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                    <SPLIT distance="100" swimtime="00:01:08.13" />
                    <SPLIT distance="150" swimtime="00:01:44.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="383" reactiontime="+85" swimtime="00:05:03.01" resultid="105047" heatid="106061" lane="7" entrytime="00:04:58.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                    <SPLIT distance="100" swimtime="00:01:12.29" />
                    <SPLIT distance="150" swimtime="00:01:50.06" />
                    <SPLIT distance="200" swimtime="00:02:28.88" />
                    <SPLIT distance="250" swimtime="00:03:07.11" />
                    <SPLIT distance="300" swimtime="00:03:46.25" />
                    <SPLIT distance="350" swimtime="00:04:24.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-05-04" firstname="Jurate" gender="F" lastname="PRANCKEVICIENE" nation="LTU" athleteid="105048">
              <RESULTS>
                <RESULT eventid="98777" points="363" reactiontime="+79" swimtime="00:00:33.26" resultid="105049" heatid="105118" lane="7" entrytime="00:00:33.33" entrycourse="LCM" />
                <RESULT eventid="98972" points="331" reactiontime="+77" swimtime="00:01:15.21" resultid="105050" heatid="105209" lane="8" entrytime="00:01:15.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="241" swimtime="00:00:40.28" resultid="105051" heatid="105261" lane="7" entrytime="00:00:39.32" entrycourse="SCM" />
                <RESULT eventid="99266" points="233" reactiontime="+81" swimtime="00:07:15.76" resultid="105052" heatid="106046" lane="8" entrytime="00:07:12.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.30" />
                    <SPLIT distance="100" swimtime="00:01:40.06" />
                    <SPLIT distance="150" swimtime="00:02:38.83" />
                    <SPLIT distance="200" swimtime="00:03:35.54" />
                    <SPLIT distance="250" swimtime="00:04:37.13" />
                    <SPLIT distance="300" swimtime="00:05:40.15" />
                    <SPLIT distance="350" swimtime="00:06:29.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-07-09" firstname="Antanas" gender="M" lastname="GUOGA" nation="LTU" swrid="4270245" athleteid="105053">
              <RESULTS>
                <RESULT eventid="98830" points="109" reactiontime="+103" swimtime="00:03:58.24" resultid="105054" heatid="105149" lane="7" entrytime="00:04:10.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.42" />
                    <SPLIT distance="100" swimtime="00:02:02.32" />
                    <SPLIT distance="150" swimtime="00:03:08.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="141" swimtime="00:27:49.91" resultid="105055" heatid="105424" lane="4" entrytime="00:26:35.99" entrycourse="SCM" />
                <RESULT eventid="99020" points="68" reactiontime="+116" swimtime="00:04:32.86" resultid="105056" heatid="105232" lane="1" entrytime="00:04:38.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.81" />
                    <SPLIT distance="100" swimtime="00:02:06.55" />
                    <SPLIT distance="150" swimtime="00:03:21.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="123" reactiontime="+114" swimtime="00:03:24.79" resultid="105057" heatid="105296" lane="1" entrytime="00:03:25.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.03" />
                    <SPLIT distance="100" swimtime="00:01:36.65" />
                    <SPLIT distance="150" swimtime="00:02:30.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="103" reactiontime="+114" swimtime="00:08:38.78" resultid="105058" heatid="106048" lane="3" entrytime="00:08:25.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.20" />
                    <SPLIT distance="100" swimtime="00:02:11.75" />
                    <SPLIT distance="150" swimtime="00:03:17.72" />
                    <SPLIT distance="200" swimtime="00:04:24.85" />
                    <SPLIT distance="250" swimtime="00:05:37.84" />
                    <SPLIT distance="300" swimtime="00:06:51.05" />
                    <SPLIT distance="350" swimtime="00:07:45.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="54" reactiontime="+92" swimtime="00:02:11.44" resultid="105059" heatid="105325" lane="8" entrytime="00:02:09.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="135" reactiontime="+106" swimtime="00:07:08.46" resultid="105060" heatid="106066" lane="6" entrytime="00:07:25.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.81" />
                    <SPLIT distance="100" swimtime="00:01:37.96" />
                    <SPLIT distance="150" swimtime="00:02:32.56" />
                    <SPLIT distance="200" swimtime="00:03:28.36" />
                    <SPLIT distance="250" swimtime="00:04:23.92" />
                    <SPLIT distance="300" swimtime="00:05:19.31" />
                    <SPLIT distance="350" swimtime="00:06:15.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-02-07" firstname="Margarita" gender="F" lastname="CINELIENE" nation="LTU" athleteid="105061">
              <RESULTS>
                <RESULT eventid="98940" points="209" reactiontime="+101" swimtime="00:03:54.22" resultid="105062" heatid="105193" lane="9" entrytime="00:03:42.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.84" />
                    <SPLIT distance="100" swimtime="00:01:50.19" />
                    <SPLIT distance="150" swimtime="00:02:52.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="230" reactiontime="+113" swimtime="00:01:44.96" resultid="105063" heatid="105245" lane="3" entrytime="00:01:43.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="253" reactiontime="+107" swimtime="00:00:46.58" resultid="105064" heatid="105347" lane="2" entrytime="00:00:44.23" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="196" reactiontime="+83" swimtime="00:02:26.01" resultid="105065" heatid="105159" lane="4" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.85" />
                    <SPLIT distance="100" swimtime="00:01:11.41" />
                    <SPLIT distance="150" swimtime="00:01:52.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="105042" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="105061" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="105053" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="105048" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" points="175" reactiontime="+89" swimtime="00:02:46.82" resultid="105066" heatid="105364" lane="9" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.47" />
                    <SPLIT distance="100" swimtime="00:01:26.55" />
                    <SPLIT distance="150" swimtime="00:02:05.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="105042" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="105061" number="2" />
                    <RELAYPOSITION athleteid="105048" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="105053" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="102089" name="Toruńczyk Masters Toruń">
          <CONTACT city="Toruń" email="szufar@o2.pl" name="Szufarski Andrzej" phone="600898866" state="KUJ-P" street="Matejki 60/7" zip="87-100" />
          <ATHLETES>
            <ATHLETE birthdate="1977-02-27" firstname="Magdalena" gender="F" lastname="ROGOZIŃSKA" nation="POL" swrid="4754678" athleteid="102090">
              <RESULTS>
                <RESULT eventid="98814" points="285" reactiontime="+108" swimtime="00:03:11.56" resultid="102091" heatid="105145" lane="0" entrytime="00:03:35.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.01" />
                    <SPLIT distance="100" swimtime="00:01:29.88" />
                    <SPLIT distance="150" swimtime="00:02:25.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="279" reactiontime="+83" swimtime="00:00:41.37" resultid="102092" heatid="105174" lane="1" entrytime="00:00:45.70" />
                <RESULT eventid="98940" points="273" reactiontime="+110" swimtime="00:03:34.18" resultid="102093" heatid="105192" lane="4" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.02" />
                    <SPLIT distance="100" swimtime="00:01:45.58" />
                    <SPLIT distance="150" swimtime="00:02:41.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="285" reactiontime="+99" swimtime="00:01:37.69" resultid="102094" heatid="105245" lane="1" entrytime="00:01:45.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="216" reactiontime="+102" swimtime="00:00:41.72" resultid="102095" heatid="105260" lane="9" entrytime="00:00:44.50" />
                <RESULT eventid="99409" points="307" reactiontime="+101" swimtime="00:00:43.67" resultid="102096" heatid="105346" lane="4" entrytime="00:00:45.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-02-06" firstname="Arkadiusz" gender="M" lastname="DOLIŃSKI" nation="POL" swrid="4992677" athleteid="102097">
              <RESULTS>
                <RESULT eventid="98798" points="384" reactiontime="+86" swimtime="00:00:28.76" resultid="102098" heatid="105130" lane="7" entrytime="00:00:32.00" />
                <RESULT eventid="98924" points="337" reactiontime="+91" swimtime="00:00:34.52" resultid="102099" heatid="105187" lane="0" entrytime="00:00:35.00" />
                <RESULT eventid="98988" points="372" reactiontime="+96" swimtime="00:01:05.21" resultid="102100" heatid="105219" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="275" reactiontime="+102" swimtime="00:00:34.47" resultid="102101" heatid="105265" lane="2" />
                <RESULT eventid="99186" points="315" reactiontime="+81" swimtime="00:01:16.26" resultid="102102" heatid="105285" lane="3" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="237" reactiontime="+88" swimtime="00:03:00.60" resultid="102103" heatid="105338" lane="6" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.75" />
                    <SPLIT distance="100" swimtime="00:01:27.55" />
                    <SPLIT distance="150" swimtime="00:02:15.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-02-16" firstname="Agnieszka" gender="F" lastname="KOSTYRA" nation="POL" swrid="4071714" athleteid="102104">
              <RESULTS>
                <RESULT eventid="98814" status="DNS" swimtime="00:00:00.00" resultid="102105" heatid="105145" lane="3" entrytime="00:03:15.00" />
                <RESULT eventid="98863" points="248" swimtime="00:13:05.30" resultid="102106" heatid="105405" lane="8" entrytime="00:12:50.00" />
                <RESULT eventid="98940" points="246" reactiontime="+87" swimtime="00:03:41.87" resultid="102107" heatid="105192" lane="2" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.23" />
                    <SPLIT distance="100" swimtime="00:01:47.35" />
                    <SPLIT distance="150" swimtime="00:02:43.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" status="DNS" swimtime="00:00:00.00" resultid="102108" heatid="105210" lane="6" entrytime="00:01:12.00" />
                <RESULT eventid="99202" status="DNS" swimtime="00:00:00.00" resultid="102109" heatid="105291" lane="1" entrytime="00:03:00.00" />
                <RESULT eventid="99266" points="258" reactiontime="+90" swimtime="00:07:01.50" resultid="102110" heatid="106046" lane="1" entrytime="00:07:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.11" />
                    <SPLIT distance="100" swimtime="00:01:47.20" />
                    <SPLIT distance="150" swimtime="00:02:43.78" />
                    <SPLIT distance="200" swimtime="00:03:37.39" />
                    <SPLIT distance="250" swimtime="00:04:32.98" />
                    <SPLIT distance="300" swimtime="00:05:28.90" />
                    <SPLIT distance="350" swimtime="00:06:15.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="284" reactiontime="+91" swimtime="00:03:08.71" resultid="102111" heatid="105333" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.34" />
                    <SPLIT distance="100" swimtime="00:01:34.38" />
                    <SPLIT distance="150" swimtime="00:02:22.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" status="WDR" swimtime="00:00:00.00" resultid="102112" entrytime="00:06:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-07-06" firstname="Andrzej" gender="M" lastname="SZUFARSKI" nation="POL" swrid="4754687" athleteid="102113">
              <RESULTS>
                <RESULT eventid="98830" points="139" reactiontime="+103" swimtime="00:03:39.99" resultid="102114" heatid="105150" lane="7" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.76" />
                    <SPLIT distance="100" swimtime="00:01:45.37" />
                    <SPLIT distance="150" swimtime="00:02:47.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="146" reactiontime="+119" swimtime="00:04:01.08" resultid="102115" heatid="105197" lane="4" entrytime="00:03:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.57" />
                    <SPLIT distance="100" swimtime="00:01:56.30" />
                    <SPLIT distance="150" swimtime="00:02:58.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="142" reactiontime="+115" swimtime="00:01:51.93" resultid="102116" heatid="105250" lane="2" entrytime="00:01:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="118" reactiontime="+118" swimtime="00:08:17.01" resultid="102117" heatid="106047" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.03" />
                    <SPLIT distance="100" swimtime="00:01:54.78" />
                    <SPLIT distance="150" swimtime="00:03:05.73" />
                    <SPLIT distance="200" swimtime="00:04:11.05" />
                    <SPLIT distance="250" swimtime="00:05:15.57" />
                    <SPLIT distance="300" swimtime="00:06:22.57" />
                    <SPLIT distance="350" swimtime="00:07:21.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="89" reactiontime="+118" swimtime="00:01:51.25" resultid="102118" heatid="105326" lane="1" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="140" reactiontime="+109" swimtime="00:00:51.30" resultid="102119" heatid="105352" lane="9" entrytime="00:00:49.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-05-05" firstname="Jarosław" gender="M" lastname="WYSOCKI" nation="POL" swrid="4992928" athleteid="102120">
              <RESULTS>
                <RESULT eventid="98830" points="127" reactiontime="+88" swimtime="00:03:46.62" resultid="102121" heatid="105150" lane="6" entrytime="00:03:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.65" />
                    <SPLIT distance="100" swimtime="00:01:44.14" />
                    <SPLIT distance="150" swimtime="00:02:46.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="182" reactiontime="+99" swimtime="00:03:43.87" resultid="102122" heatid="105198" lane="5" entrytime="00:03:42.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.58" />
                    <SPLIT distance="100" swimtime="00:01:49.37" />
                    <SPLIT distance="150" swimtime="00:02:47.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="196" reactiontime="+101" swimtime="00:01:40.48" resultid="102123" heatid="105251" lane="0" entrytime="00:01:40.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="230" reactiontime="+94" swimtime="00:00:43.52" resultid="102124" heatid="105354" lane="1" entrytime="00:00:43.34" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-03-03" firstname="Henryk" gender="M" lastname="ZIENTARA" nation="POL" swrid="4754680" athleteid="102125">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="102126" heatid="105124" lane="5" entrytime="00:00:41.30" />
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="102127" heatid="105149" lane="0" entrytime="00:04:18.25" />
                <RESULT eventid="98924" points="99" reactiontime="+79" swimtime="00:00:51.95" resultid="102128" heatid="105181" lane="3" entrytime="00:00:53.65" />
                <RESULT eventid="98956" points="105" reactiontime="+110" swimtime="00:04:29.15" resultid="102129" heatid="105196" lane="3" entrytime="00:04:21.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.89" />
                    <SPLIT distance="100" swimtime="00:02:05.48" />
                    <SPLIT distance="150" swimtime="00:03:18.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="111" reactiontime="+104" swimtime="00:02:01.48" resultid="102130" heatid="105249" lane="4" entrytime="00:01:54.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="62" reactiontime="+86" swimtime="00:02:11.02" resultid="102131" heatid="105281" lane="6" entrytime="00:02:05.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="139" reactiontime="+102" swimtime="00:00:51.39" resultid="102132" heatid="105352" lane="8" entrytime="00:00:48.21" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-08-21" firstname="Tomasz" gender="M" lastname="OSÓBKA" nation="POL" swrid="4992926" athleteid="102133">
              <RESULTS>
                <RESULT eventid="98798" points="35" reactiontime="+118" swimtime="00:01:03.48" resultid="102134" heatid="105123" lane="5" entrytime="00:00:59.58" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="102135" heatid="105213" lane="1" entrytime="00:02:45.25" />
                <RESULT eventid="99091" points="17" reactiontime="+126" swimtime="00:03:45.19" resultid="102136" heatid="105249" lane="1" entrytime="00:03:42.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:39.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="20" reactiontime="+113" swimtime="00:01:38.15" resultid="102137" heatid="105351" lane="8" entrytime="00:01:35.58" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-10-13" firstname="Edward" gender="M" lastname="KOROLKO" nation="POL" swrid="4754683" athleteid="102138">
              <RESULTS>
                <RESULT eventid="98798" points="137" reactiontime="+102" swimtime="00:00:40.55" resultid="102139" heatid="105124" lane="4" entrytime="00:00:40.25" />
                <RESULT eventid="98924" points="60" reactiontime="+85" swimtime="00:01:01.34" resultid="102140" heatid="105181" lane="8" entrytime="00:00:55.80" />
                <RESULT eventid="98988" points="98" reactiontime="+100" swimtime="00:01:41.64" resultid="102141" heatid="105214" lane="9" entrytime="00:01:36.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="52" reactiontime="+94" swimtime="00:02:19.10" resultid="102142" heatid="105281" lane="3" entrytime="00:02:05.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="102143" heatid="105336" lane="7" entrytime="00:04:40.12" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-03-07" firstname="Grzegorz" gender="M" lastname="ARENTEWICZ" nation="POL" swrid="4754686" athleteid="102144">
              <RESULTS>
                <RESULT eventid="98830" points="277" reactiontime="+89" swimtime="00:02:54.81" resultid="102145" heatid="105151" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                    <SPLIT distance="100" swimtime="00:01:23.47" />
                    <SPLIT distance="150" swimtime="00:02:15.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" status="DNS" swimtime="00:00:00.00" resultid="102146" heatid="105182" lane="3" entrytime="00:00:48.00" />
                <RESULT eventid="99020" points="188" reactiontime="+103" swimtime="00:03:14.53" resultid="102147" heatid="105234" lane="7" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.02" />
                    <SPLIT distance="100" swimtime="00:01:33.31" />
                    <SPLIT distance="150" swimtime="00:02:26.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="249" reactiontime="+101" swimtime="00:02:42.09" resultid="102148" heatid="105299" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                    <SPLIT distance="100" swimtime="00:01:14.29" />
                    <SPLIT distance="150" swimtime="00:01:57.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" status="DNS" swimtime="00:00:00.00" resultid="102149" heatid="106050" lane="6" entrytime="00:06:45.00" />
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="102150" heatid="105328" lane="9" entrytime="00:01:25.00" />
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="102151" entrytime="00:05:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-07-25" firstname="Sławomir" gender="M" lastname="PRĘDKI" nation="POL" swrid="4041308" athleteid="102152">
              <RESULTS>
                <RESULT eventid="98798" points="503" reactiontime="+83" swimtime="00:00:26.29" resultid="102153" heatid="105134" lane="1" entrytime="00:00:30.00" />
                <RESULT eventid="98830" points="532" reactiontime="+85" swimtime="00:02:20.61" resultid="102154" heatid="105152" lane="4" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                    <SPLIT distance="100" swimtime="00:01:05.74" />
                    <SPLIT distance="150" swimtime="00:01:47.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="497" swimtime="00:02:40.29" resultid="102155" heatid="105204" lane="7" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                    <SPLIT distance="100" swimtime="00:01:16.00" />
                    <SPLIT distance="150" swimtime="00:01:58.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="541" reactiontime="+75" swimtime="00:00:57.57" resultid="102156" heatid="105222" lane="9" entrytime="00:01:05.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="517" reactiontime="+92" swimtime="00:01:12.81" resultid="102157" heatid="105252" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="508" reactiontime="+79" swimtime="00:02:07.76" resultid="102158" heatid="105301" lane="9" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.26" />
                    <SPLIT distance="100" swimtime="00:01:02.36" />
                    <SPLIT distance="150" swimtime="00:01:35.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="526" reactiontime="+89" swimtime="00:00:33.03" resultid="102159" heatid="105352" lane="1" entrytime="00:00:48.10" />
                <RESULT eventid="99473" points="514" reactiontime="+71" swimtime="00:04:34.56" resultid="102160" heatid="106063" lane="8" entrytime="00:05:45.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                    <SPLIT distance="100" swimtime="00:01:04.00" />
                    <SPLIT distance="150" swimtime="00:01:38.80" />
                    <SPLIT distance="200" swimtime="00:02:14.33" />
                    <SPLIT distance="250" swimtime="00:02:49.75" />
                    <SPLIT distance="300" swimtime="00:03:25.66" />
                    <SPLIT distance="350" swimtime="00:04:00.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-07-04" firstname="Karol" gender="M" lastname="TWAROWSKI" nation="POL" swrid="4967387" athleteid="102161">
              <RESULTS>
                <RESULT eventid="98830" points="458" reactiontime="+87" swimtime="00:02:27.87" resultid="102162" heatid="105151" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.57" />
                    <SPLIT distance="100" swimtime="00:01:06.82" />
                    <SPLIT distance="150" swimtime="00:01:50.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="402" swimtime="00:19:39.47" resultid="102163" heatid="105421" lane="2" entrytime="00:21:00.00" />
                <RESULT eventid="98924" points="421" reactiontime="+84" swimtime="00:00:32.07" resultid="102164" heatid="105184" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="99020" points="346" reactiontime="+104" swimtime="00:02:38.79" resultid="102165" heatid="105231" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                    <SPLIT distance="100" swimtime="00:01:11.41" />
                    <SPLIT distance="150" swimtime="00:01:53.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="420" reactiontime="+79" swimtime="00:01:09.34" resultid="102166" heatid="105283" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="426" reactiontime="+97" swimtime="00:05:24.06" resultid="102167" heatid="106051" lane="0" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.78" />
                    <SPLIT distance="100" swimtime="00:01:10.74" />
                    <SPLIT distance="150" swimtime="00:01:52.89" />
                    <SPLIT distance="200" swimtime="00:02:34.29" />
                    <SPLIT distance="250" swimtime="00:03:20.20" />
                    <SPLIT distance="300" swimtime="00:04:06.78" />
                    <SPLIT distance="350" swimtime="00:04:46.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="102168" heatid="105327" lane="4" entrytime="00:01:25.00" />
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="102169" heatid="105338" lane="3" entrytime="00:03:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-01" firstname="Katarzyna" gender="F" lastname="WALENTA" nation="POL" swrid="4754689" athleteid="102170">
              <RESULTS>
                <RESULT eventid="98777" points="447" reactiontime="+100" swimtime="00:00:31.03" resultid="102171" heatid="105120" lane="1" entrytime="00:00:30.34" entrycourse="SCM" />
                <RESULT eventid="98814" points="409" reactiontime="+94" swimtime="00:02:49.91" resultid="102172" heatid="105146" lane="5" entrytime="00:02:56.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                    <SPLIT distance="100" swimtime="00:01:18.85" />
                    <SPLIT distance="150" swimtime="00:02:07.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="390" reactiontime="+84" swimtime="00:00:37.03" resultid="102173" heatid="105178" lane="7" entrytime="00:00:34.50" />
                <RESULT eventid="99004" points="232" reactiontime="+92" swimtime="00:03:18.13" resultid="102174" heatid="105230" lane="6" entrytime="00:03:10.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.23" />
                    <SPLIT distance="100" swimtime="00:01:28.11" />
                    <SPLIT distance="150" swimtime="00:02:21.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="405" reactiontime="+94" swimtime="00:00:33.88" resultid="102175" heatid="105263" lane="1" entrytime="00:00:34.20" />
                <RESULT eventid="99266" points="373" reactiontime="+96" swimtime="00:06:12.72" resultid="102176" heatid="106046" lane="3" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                    <SPLIT distance="100" swimtime="00:01:26.62" />
                    <SPLIT distance="150" swimtime="00:02:14.47" />
                    <SPLIT distance="200" swimtime="00:03:00.92" />
                    <SPLIT distance="250" swimtime="00:03:51.17" />
                    <SPLIT distance="300" swimtime="00:04:43.04" />
                    <SPLIT distance="350" swimtime="00:05:28.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="358" reactiontime="+91" swimtime="00:01:18.79" resultid="102177" heatid="105323" lane="0" entrytime="00:01:19.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="371" reactiontime="+84" swimtime="00:00:41.01" resultid="102178" heatid="105349" lane="9" entrytime="00:00:39.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-08-03" firstname="Artur" gender="M" lastname="KŁOSIŃSKI" nation="POL" swrid="4754685" athleteid="102179">
              <RESULTS>
                <RESULT eventid="98798" points="434" reactiontime="+88" swimtime="00:00:27.61" resultid="102180" heatid="105123" lane="0" />
                <RESULT eventid="98830" points="336" reactiontime="+80" swimtime="00:02:43.88" resultid="102181" heatid="105155" lane="7" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                    <SPLIT distance="100" swimtime="00:01:17.03" />
                    <SPLIT distance="150" swimtime="00:02:06.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="352" reactiontime="+79" swimtime="00:00:34.02" resultid="102182" heatid="105179" lane="5" />
                <RESULT eventid="98956" status="DNS" swimtime="00:00:00.00" resultid="102183" heatid="105202" lane="4" entrytime="00:03:00.00" />
                <RESULT eventid="99186" points="338" reactiontime="+85" swimtime="00:01:14.53" resultid="102184" heatid="105286" lane="3" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" status="DNS" swimtime="00:00:00.00" resultid="102185" heatid="106051" lane="4" entrytime="00:06:00.00" />
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="102186" heatid="105340" lane="2" entrytime="00:02:50.00" />
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="102187" entrytime="00:05:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-02-03" firstname="Maciej" gender="M" lastname="KURAS" nation="POL" swrid="4754691" athleteid="102188">
              <RESULTS>
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="102189" heatid="105271" lane="0" entrytime="00:00:32.49" />
                <RESULT eventid="99186" status="DNS" swimtime="00:00:00.00" resultid="102190" heatid="105285" lane="9" entrytime="00:01:18.23" />
                <RESULT eventid="99393" points="274" reactiontime="+93" swimtime="00:02:52.23" resultid="102191" heatid="105340" lane="5" entrytime="00:02:49.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.97" />
                    <SPLIT distance="100" swimtime="00:01:23.55" />
                    <SPLIT distance="150" swimtime="00:02:07.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-04-23" firstname="Krzysztof" gender="M" lastname="LIETZ" nation="POL" swrid="4754688" athleteid="102192">
              <RESULTS>
                <RESULT eventid="98798" points="279" reactiontime="+86" swimtime="00:00:31.98" resultid="102193" heatid="105129" lane="4" entrytime="00:00:32.50" />
                <RESULT eventid="98830" points="186" reactiontime="+89" swimtime="00:03:19.69" resultid="102194" heatid="105151" lane="3" entrytime="00:03:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                    <SPLIT distance="100" swimtime="00:01:42.01" />
                    <SPLIT distance="150" swimtime="00:02:38.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="267" reactiontime="+98" swimtime="00:01:12.76" resultid="102195" heatid="105218" lane="1" entrytime="00:01:11.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="230" reactiontime="+86" swimtime="00:00:36.58" resultid="102196" heatid="105268" lane="5" entrytime="00:00:35.80" />
                <RESULT eventid="99218" points="212" reactiontime="+88" swimtime="00:02:50.91" resultid="102197" heatid="105298" lane="6" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.73" />
                    <SPLIT distance="100" swimtime="00:01:24.59" />
                    <SPLIT distance="150" swimtime="00:02:11.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="175" reactiontime="+97" swimtime="00:01:29.03" resultid="102198" heatid="105327" lane="3" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="206" reactiontime="+113" swimtime="00:06:12.32" resultid="102199" heatid="106065" lane="5" entrytime="00:06:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.98" />
                    <SPLIT distance="100" swimtime="00:01:28.35" />
                    <SPLIT distance="150" swimtime="00:02:16.73" />
                    <SPLIT distance="200" swimtime="00:03:06.29" />
                    <SPLIT distance="250" swimtime="00:03:54.55" />
                    <SPLIT distance="300" swimtime="00:04:43.82" />
                    <SPLIT distance="350" swimtime="00:05:30.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-02-16" firstname="Maciej" gender="M" lastname="KUJAWA" nation="POL" swrid="4992927" athleteid="102200">
              <RESULTS>
                <RESULT eventid="98830" points="217" reactiontime="+99" swimtime="00:03:09.45" resultid="102201" heatid="105148" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                    <SPLIT distance="100" swimtime="00:01:29.37" />
                    <SPLIT distance="150" swimtime="00:02:23.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="239" reactiontime="+87" swimtime="00:03:24.41" resultid="102202" heatid="105196" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.17" />
                    <SPLIT distance="100" swimtime="00:01:33.93" />
                    <SPLIT distance="150" swimtime="00:02:28.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="267" reactiontime="+95" swimtime="00:01:30.68" resultid="102203" heatid="105249" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="284" reactiontime="+83" swimtime="00:00:40.55" resultid="102204" heatid="105351" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-19" firstname="Tomasz" gender="M" lastname="ZASADOWSKI" nation="POL" athleteid="102205">
              <RESULTS>
                <RESULT eventid="98798" points="373" reactiontime="+85" swimtime="00:00:29.03" resultid="102206" heatid="105123" lane="9" />
                <RESULT eventid="98924" points="308" reactiontime="+69" swimtime="00:00:35.57" resultid="102207" heatid="105180" lane="8" />
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="102208" heatid="105265" lane="0" />
                <RESULT eventid="99186" points="270" reactiontime="+81" swimtime="00:01:20.27" resultid="102209" heatid="105281" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="247" reactiontime="+89" swimtime="00:01:19.36" resultid="102210" heatid="105324" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-03-24" firstname="Dariusz" gender="M" lastname="PELA" nation="POL" swrid="4992925" athleteid="102211">
              <RESULTS>
                <RESULT eventid="98798" points="303" reactiontime="+96" swimtime="00:00:31.11" resultid="102212" heatid="105129" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="98988" points="242" reactiontime="+109" swimtime="00:01:15.21" resultid="102213" heatid="105217" lane="0" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="237" reactiontime="+91" swimtime="00:01:34.45" resultid="102214" heatid="105252" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="270" reactiontime="+99" swimtime="00:00:41.24" resultid="102215" heatid="105356" lane="2" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="99059" points="64" reactiontime="+80" swimtime="00:03:52.76" resultid="102218" heatid="105239" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.95" />
                    <SPLIT distance="100" swimtime="00:03:52.94" />
                    <SPLIT distance="150" swimtime="00:03:11.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102125" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="102133" number="2" reactiontime="+111" />
                    <RELAYPOSITION athleteid="102113" number="3" />
                    <RELAYPOSITION athleteid="102138" number="4" reactiontime="+89" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" points="79" reactiontime="+103" swimtime="00:03:17.47" resultid="102219" heatid="105309" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.64" />
                    <SPLIT distance="100" swimtime="00:01:48.33" />
                    <SPLIT distance="150" swimtime="00:02:35.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102138" number="1" reactiontime="+103" />
                    <RELAYPOSITION athleteid="102133" number="2" reactiontime="+79" />
                    <RELAYPOSITION athleteid="102125" number="3" reactiontime="+79" />
                    <RELAYPOSITION athleteid="102113" number="4" reactiontime="+94" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="99059" points="380" reactiontime="+80" swimtime="00:02:08.97" resultid="102220" heatid="105242" lane="6" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.91" />
                    <SPLIT distance="100" swimtime="00:01:05.46" />
                    <SPLIT distance="150" swimtime="00:01:41.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102161" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="102152" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="102192" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="102179" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" points="440" reactiontime="+65" swimtime="00:01:51.54" resultid="102221" heatid="105311" lane="8" entrytime="00:01:54.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.33" />
                    <SPLIT distance="100" swimtime="00:00:52.58" />
                    <SPLIT distance="150" swimtime="00:01:24.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102152" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="102161" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="102192" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="102179" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="99059" points="287" reactiontime="+80" swimtime="00:02:21.57" resultid="102222" heatid="105241" lane="1" entrytime="00:02:19.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                    <SPLIT distance="100" swimtime="00:01:16.63" />
                    <SPLIT distance="150" swimtime="00:01:52.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102097" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="102120" number="2" reactiontime="+67" />
                    <RELAYPOSITION athleteid="102200" number="3" reactiontime="+65" />
                    <RELAYPOSITION athleteid="102205" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="99250" status="DNS" swimtime="00:00:00.00" resultid="102223" heatid="105310" lane="0" entrytime="00:02:07.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102188" number="1" />
                    <RELAYPOSITION athleteid="102120" number="2" />
                    <RELAYPOSITION athleteid="102200" number="3" />
                    <RELAYPOSITION athleteid="102144" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="381" reactiontime="+104" swimtime="00:01:57.02" resultid="102216" heatid="105159" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                    <SPLIT distance="100" swimtime="00:01:00.46" />
                    <SPLIT distance="150" swimtime="00:01:30.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102090" number="1" reactiontime="+104" />
                    <RELAYPOSITION athleteid="102152" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="102170" number="3" reactiontime="+70" />
                    <RELAYPOSITION athleteid="102161" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" status="DNS" swimtime="00:00:00.00" resultid="102217" heatid="105365" lane="9" entrytime="00:02:18.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102090" number="1" />
                    <RELAYPOSITION athleteid="102152" number="2" />
                    <RELAYPOSITION athleteid="102170" number="3" />
                    <RELAYPOSITION athleteid="102161" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="102927" name="UJCM KRAKÓW">
          <ATHLETES>
            <ATHLETE birthdate="1992-08-23" firstname="Magdalena" gender="F" lastname="DRAB" nation="POL" swrid="4072271" athleteid="102928">
              <RESULTS>
                <RESULT eventid="98777" points="531" reactiontime="+98" swimtime="00:00:29.30" resultid="102996" heatid="105121" lane="0" entrytime="00:00:29.18" entrycourse="LCM" />
                <RESULT eventid="98814" points="578" reactiontime="+91" swimtime="00:02:31.38" resultid="102997" heatid="105147" lane="4" entrytime="00:02:35.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.42" />
                    <SPLIT distance="100" swimtime="00:01:12.19" />
                    <SPLIT distance="150" swimtime="00:01:55.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="441" reactiontime="+92" swimtime="00:03:02.67" resultid="102998" heatid="105194" lane="4" entrytime="00:02:59.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.10" />
                    <SPLIT distance="100" swimtime="00:01:26.19" />
                    <SPLIT distance="150" swimtime="00:02:14.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="592" swimtime="00:01:02.00" resultid="102999" heatid="105212" lane="7" entrytime="00:01:02.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="459" reactiontime="+91" swimtime="00:01:23.40" resultid="103000" heatid="105247" lane="4" entrytime="00:01:22.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="582" reactiontime="+96" swimtime="00:02:15.31" resultid="103001" heatid="105294" lane="3" entrytime="00:02:14.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                    <SPLIT distance="100" swimtime="00:01:05.78" />
                    <SPLIT distance="150" swimtime="00:01:41.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="550" reactiontime="+84" swimtime="00:00:35.96" resultid="103002" heatid="105349" lane="6" entrytime="00:00:36.92" />
                <RESULT eventid="99457" points="569" reactiontime="+92" swimtime="00:04:48.45" resultid="103003" heatid="106054" lane="5" entrytime="00:04:49.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                    <SPLIT distance="100" swimtime="00:01:08.27" />
                    <SPLIT distance="150" swimtime="00:01:45.32" />
                    <SPLIT distance="200" swimtime="00:02:22.53" />
                    <SPLIT distance="250" swimtime="00:03:00.36" />
                    <SPLIT distance="300" swimtime="00:03:38.03" />
                    <SPLIT distance="350" swimtime="00:04:14.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04514" nation="POL" region="MAZ" clubid="100410" name="UKS 307 Warszawa Mokotów">
          <CONTACT name="Ilczyszyn" />
          <ATHLETES>
            <ATHLETE birthdate="1978-02-03" firstname="Damian" gender="M" lastname="ZIÓŁKOWSKI" nation="POL" swrid="4992934" athleteid="100411">
              <RESULTS>
                <RESULT eventid="98798" points="385" reactiontime="+88" swimtime="00:00:28.74" resultid="100412" heatid="105139" lane="2" entrytime="00:00:27.50" />
                <RESULT eventid="99091" points="297" reactiontime="+81" swimtime="00:01:27.59" resultid="100413" heatid="105254" lane="9" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="345" reactiontime="+87" swimtime="00:00:31.96" resultid="100414" heatid="105272" lane="6" entrytime="00:00:31.00" />
                <RESULT eventid="99473" points="303" reactiontime="+85" swimtime="00:05:27.30" resultid="100415" heatid="106062" lane="6" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                    <SPLIT distance="100" swimtime="00:01:14.34" />
                    <SPLIT distance="150" swimtime="00:01:55.95" />
                    <SPLIT distance="200" swimtime="00:02:38.98" />
                    <SPLIT distance="250" swimtime="00:03:22.81" />
                    <SPLIT distance="300" swimtime="00:04:06.33" />
                    <SPLIT distance="350" swimtime="00:04:49.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00408" nation="POL" region="RZ" clubid="100150" name="UKS Delfin Masters Tarnobrzeg">
          <CONTACT city="TARNOBRZEG" email="piotr.michaliki-bs.pl" name="MICHALIK ANGELIKA" state="PODKA" street="SKALNA GÓRA 8/21" street2="TARNOBRZEG" zip="39-400" />
          <ATHLETES>
            <ATHLETE birthdate="1984-02-08" firstname="Adrian" gender="M" lastname="MARSZAŁEK" nation="POL" athleteid="100151">
              <RESULTS>
                <RESULT eventid="98798" points="367" reactiontime="+80" swimtime="00:00:29.19" resultid="100152" heatid="105140" lane="1" entrytime="00:00:27.00" />
                <RESULT eventid="98956" points="305" reactiontime="+83" swimtime="00:03:08.60" resultid="100153" heatid="105203" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.58" />
                    <SPLIT distance="100" swimtime="00:01:27.49" />
                    <SPLIT distance="150" swimtime="00:02:16.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="325" reactiontime="+95" swimtime="00:01:24.97" resultid="100154" heatid="105257" lane="0" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="396" reactiontime="+80" swimtime="00:00:36.31" resultid="100155" heatid="105361" lane="5" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-04-27" firstname="Kamil" gender="M" lastname="ZIELIŃSKI" nation="POL" swrid="4071551" athleteid="100156">
              <RESULTS>
                <RESULT eventid="98798" points="474" reactiontime="+76" swimtime="00:00:26.80" resultid="100157" heatid="105142" lane="2" entrytime="00:00:26.00" />
                <RESULT eventid="98830" points="453" reactiontime="+75" swimtime="00:02:28.42" resultid="100158" heatid="105157" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.45" />
                    <SPLIT distance="100" swimtime="00:01:12.77" />
                    <SPLIT distance="150" swimtime="00:01:52.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="568" reactiontime="+73" swimtime="00:02:33.33" resultid="100159" heatid="105204" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.15" />
                    <SPLIT distance="100" swimtime="00:01:13.84" />
                    <SPLIT distance="150" swimtime="00:01:54.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="621" reactiontime="+79" swimtime="00:01:08.50" resultid="100160" heatid="105258" lane="4" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="448" reactiontime="+80" swimtime="00:00:29.31" resultid="100161" heatid="105275" lane="1" entrytime="00:00:28.00" />
                <RESULT eventid="99425" points="653" reactiontime="+71" swimtime="00:00:30.73" resultid="100162" heatid="105362" lane="4" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-04-24" firstname="Renata" gender="F" lastname="OSMALA" nation="POL" swrid="4992935" athleteid="100163">
              <RESULTS>
                <RESULT eventid="98863" points="376" reactiontime="+65" swimtime="00:11:23.85" resultid="100164" heatid="105404" lane="9" entrytime="00:11:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.07" />
                    <SPLIT distance="100" swimtime="00:01:18.42" />
                    <SPLIT distance="150" swimtime="00:02:01.06" />
                    <SPLIT distance="200" swimtime="00:02:44.71" />
                    <SPLIT distance="250" swimtime="00:03:28.10" />
                    <SPLIT distance="300" swimtime="00:04:11.87" />
                    <SPLIT distance="350" swimtime="00:04:55.77" />
                    <SPLIT distance="400" swimtime="00:05:39.32" />
                    <SPLIT distance="450" swimtime="00:06:22.89" />
                    <SPLIT distance="500" swimtime="00:07:06.50" />
                    <SPLIT distance="550" swimtime="00:07:49.97" />
                    <SPLIT distance="600" swimtime="00:08:33.47" />
                    <SPLIT distance="650" swimtime="00:09:17.22" />
                    <SPLIT distance="700" swimtime="00:10:00.14" />
                    <SPLIT distance="750" swimtime="00:10:43.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="335" reactiontime="+71" swimtime="00:00:38.93" resultid="100165" heatid="105177" lane="6" entrytime="00:00:37.50" />
                <RESULT eventid="98940" points="344" swimtime="00:03:18.42" resultid="100166" heatid="105194" lane="0" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.23" />
                    <SPLIT distance="100" swimtime="00:01:34.05" />
                    <SPLIT distance="150" swimtime="00:02:25.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="366" reactiontime="+69" swimtime="00:01:29.91" resultid="100167" heatid="105247" lane="7" entrytime="00:01:28.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="336" reactiontime="+81" swimtime="00:01:23.58" resultid="100168" heatid="105280" lane="8" entrytime="00:01:21.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.27" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99377" points="363" reactiontime="+82" swimtime="00:02:53.88" resultid="100169" heatid="105334" lane="2" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                    <SPLIT distance="100" swimtime="00:01:25.67" />
                    <SPLIT distance="150" swimtime="00:02:10.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="368" reactiontime="+90" swimtime="00:00:41.13" resultid="100170" heatid="105348" lane="2" entrytime="00:00:41.55" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-01" firstname="Beata" gender="F" lastname="KACZMARCZYK" nation="POL" swrid="4992940" athleteid="100171">
              <RESULTS>
                <RESULT eventid="98777" points="272" reactiontime="+79" swimtime="00:00:36.62" resultid="100172" heatid="105117" lane="6" entrytime="00:00:34.69" entrycourse="SCM" />
                <RESULT eventid="98907" points="259" reactiontime="+73" swimtime="00:00:42.41" resultid="100173" heatid="105175" lane="0" entrytime="00:00:42.00" />
                <RESULT eventid="98972" points="260" reactiontime="+93" swimtime="00:01:21.48" resultid="100174" heatid="105207" lane="4" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="245" reactiontime="+94" swimtime="00:03:00.49" resultid="100175" heatid="105291" lane="7" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.29" />
                    <SPLIT distance="100" swimtime="00:01:24.86" />
                    <SPLIT distance="150" swimtime="00:02:12.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="260" reactiontime="+95" swimtime="00:06:14.67" resultid="100176" heatid="106056" lane="4" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.32" />
                    <SPLIT distance="100" swimtime="00:01:29.66" />
                    <SPLIT distance="150" swimtime="00:02:17.90" />
                    <SPLIT distance="200" swimtime="00:03:06.53" />
                    <SPLIT distance="250" swimtime="00:03:54.35" />
                    <SPLIT distance="300" swimtime="00:04:43.07" />
                    <SPLIT distance="350" swimtime="00:05:30.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-03-28" firstname="Agata" gender="F" lastname="MEKSUŁA" nation="POL" swrid="4992937" athleteid="100177">
              <RESULTS>
                <RESULT eventid="98777" points="396" reactiontime="+84" swimtime="00:00:32.30" resultid="100178" heatid="105119" lane="1" entrytime="00:00:31.86" entrycourse="SCM" />
                <RESULT eventid="98972" points="395" reactiontime="+100" swimtime="00:01:10.94" resultid="100179" heatid="105209" lane="5" entrytime="00:01:14.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="281" reactiontime="+95" swimtime="00:00:38.24" resultid="100180" heatid="105261" lane="2" entrytime="00:00:39.10" />
                <RESULT eventid="99202" points="344" reactiontime="+109" swimtime="00:02:41.09" resultid="100181" heatid="105293" lane="0" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.96" />
                    <SPLIT distance="100" swimtime="00:01:19.25" />
                    <SPLIT distance="150" swimtime="00:02:00.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="318" reactiontime="+89" swimtime="00:05:50.33" resultid="100182" heatid="106054" lane="9" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.14" />
                    <SPLIT distance="100" swimtime="00:01:22.54" />
                    <SPLIT distance="150" swimtime="00:02:08.18" />
                    <SPLIT distance="200" swimtime="00:02:53.94" />
                    <SPLIT distance="250" swimtime="00:03:39.57" />
                    <SPLIT distance="300" swimtime="00:04:24.48" />
                    <SPLIT distance="350" swimtime="00:05:09.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-07-14" firstname="Aneta" gender="F" lastname="MADEJ" nation="POL" athleteid="100183">
              <RESULTS>
                <RESULT eventid="98940" points="328" reactiontime="+106" swimtime="00:03:21.51" resultid="100184" heatid="105191" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.15" />
                    <SPLIT distance="100" swimtime="00:01:32.82" />
                    <SPLIT distance="150" swimtime="00:02:26.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="331" reactiontime="+98" swimtime="00:01:33.01" resultid="100185" heatid="105246" lane="0" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="334" reactiontime="+84" swimtime="00:00:42.46" resultid="100186" heatid="105347" lane="9" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-17" firstname="Sławomir" gender="M" lastname="KOWALSKI" nation="POL" swrid="4992948" athleteid="100187">
              <RESULTS>
                <RESULT eventid="98830" points="320" reactiontime="+89" swimtime="00:02:46.59" resultid="100188" heatid="105154" lane="3" entrytime="00:02:45.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                    <SPLIT distance="100" swimtime="00:01:18.77" />
                    <SPLIT distance="150" swimtime="00:02:05.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="340" swimtime="00:03:01.96" resultid="100189" heatid="105203" lane="7" entrytime="00:02:57.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.30" />
                    <SPLIT distance="100" swimtime="00:01:25.99" />
                    <SPLIT distance="150" swimtime="00:02:13.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="382" reactiontime="+98" swimtime="00:01:20.53" resultid="100190" heatid="105255" lane="1" entrytime="00:01:22.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="417" reactiontime="+87" swimtime="00:00:35.69" resultid="100191" heatid="105358" lane="4" entrytime="00:00:36.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-03-03" firstname="Patrycja" gender="F" lastname="URBANIAK" nation="POL" swrid="4072332" athleteid="100192">
              <RESULTS>
                <RESULT eventid="98972" status="DNS" swimtime="00:00:00.00" resultid="100193" heatid="105211" lane="6" entrytime="00:01:06.58" />
                <RESULT eventid="99004" points="255" reactiontime="+94" swimtime="00:03:11.97" resultid="100194" heatid="105230" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.21" />
                    <SPLIT distance="100" swimtime="00:01:24.07" />
                    <SPLIT distance="150" swimtime="00:02:16.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="416" reactiontime="+76" swimtime="00:00:33.58" resultid="100195" heatid="105264" lane="0" entrytime="00:00:32.73" />
                <RESULT eventid="99202" status="DNS" swimtime="00:00:00.00" resultid="100196" heatid="105293" lane="4" entrytime="00:02:28.50" />
                <RESULT eventid="99344" points="365" reactiontime="+66" swimtime="00:01:18.30" resultid="100197" heatid="105323" lane="8" entrytime="00:01:17.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-12" firstname="Maciej" gender="M" lastname="PŁANETA" nation="POL" swrid="4992944" athleteid="100198">
              <RESULTS>
                <RESULT eventid="98798" points="297" reactiontime="+77" swimtime="00:00:31.33" resultid="100199" heatid="105132" lane="4" entrytime="00:00:30.50" />
                <RESULT eventid="98988" points="287" reactiontime="+95" swimtime="00:01:11.04" resultid="100200" heatid="105220" lane="0" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="230" reactiontime="+89" swimtime="00:00:36.59" resultid="100201" heatid="105268" lane="4" entrytime="00:00:35.55" />
                <RESULT eventid="99218" points="248" reactiontime="+80" swimtime="00:02:42.25" resultid="100202" heatid="105300" lane="9" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.86" />
                    <SPLIT distance="100" swimtime="00:01:19.67" />
                    <SPLIT distance="150" swimtime="00:02:02.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="269" reactiontime="+92" swimtime="00:05:40.87" resultid="100203" heatid="106063" lane="5" entrytime="00:05:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                    <SPLIT distance="100" swimtime="00:01:19.13" />
                    <SPLIT distance="150" swimtime="00:02:02.83" />
                    <SPLIT distance="200" swimtime="00:02:48.09" />
                    <SPLIT distance="250" swimtime="00:03:32.50" />
                    <SPLIT distance="300" swimtime="00:04:17.41" />
                    <SPLIT distance="350" swimtime="00:05:01.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="270" swimtime="00:22:26.53" resultid="102069" heatid="105422" lane="8" entrytime="00:22:45.77" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-15" firstname="Paweł" gender="M" lastname="NOWAK" nation="POL" swrid="4992947" athleteid="100204">
              <RESULTS>
                <RESULT comment="04" eventid="98798" reactiontime="+69" status="DSQ" swimtime="00:00:00.00" resultid="100205" heatid="105134" lane="9" entrytime="00:00:30.00" />
                <RESULT eventid="98924" points="278" reactiontime="+78" swimtime="00:00:36.80" resultid="100206" heatid="105186" lane="3" entrytime="00:00:36.00" />
                <RESULT eventid="99170" points="283" reactiontime="+93" swimtime="00:00:34.15" resultid="100207" heatid="105267" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="99186" status="DNS" swimtime="00:00:00.00" resultid="100208" heatid="105284" lane="8" entrytime="00:01:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-23" firstname="Krzysztof" gender="M" lastname="ŚLĘCZKA" nation="POL" swrid="4992942" athleteid="100209">
              <RESULTS>
                <RESULT eventid="98798" points="420" reactiontime="+73" swimtime="00:00:27.92" resultid="100210" heatid="105139" lane="7" entrytime="00:00:27.50" />
                <RESULT eventid="98891" status="WDR" swimtime="00:00:00.00" resultid="100211" entrytime="00:21:00.00" />
                <RESULT eventid="98924" points="317" reactiontime="+77" swimtime="00:00:35.25" resultid="100212" heatid="105187" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="98988" points="436" reactiontime="+78" swimtime="00:01:01.85" resultid="100213" heatid="105223" lane="5" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="396" reactiontime="+80" swimtime="00:00:30.52" resultid="100214" heatid="105271" lane="3" entrytime="00:00:31.50" />
                <RESULT eventid="99218" points="356" reactiontime="+86" swimtime="00:02:23.83" resultid="100215" heatid="105301" lane="2" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                    <SPLIT distance="100" swimtime="00:01:09.53" />
                    <SPLIT distance="150" swimtime="00:01:47.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="296" reactiontime="+85" swimtime="00:01:14.68" resultid="100216" heatid="105329" lane="2" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="314" reactiontime="+84" swimtime="00:05:23.50" resultid="100217" heatid="106062" lane="0" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.55" />
                    <SPLIT distance="100" swimtime="00:01:13.97" />
                    <SPLIT distance="150" swimtime="00:01:54.82" />
                    <SPLIT distance="200" swimtime="00:02:36.56" />
                    <SPLIT distance="250" swimtime="00:03:18.61" />
                    <SPLIT distance="300" swimtime="00:04:01.24" />
                    <SPLIT distance="350" swimtime="00:04:43.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-25" firstname="Artur" gender="M" lastname="SZKLARZ" nation="POL" swrid="4992946" athleteid="100218">
              <RESULTS>
                <RESULT eventid="98798" points="332" reactiontime="+75" swimtime="00:00:30.19" resultid="100219" heatid="105137" lane="6" entrytime="00:00:28.50" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="100220" heatid="105222" lane="6" entrytime="00:01:04.50" />
                <RESULT eventid="99020" reactiontime="+85" status="DNF" swimtime="00:00:00.00" resultid="100221" heatid="105235" lane="0" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.14" />
                    <SPLIT distance="100" swimtime="00:01:26.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="325" reactiontime="+79" swimtime="00:00:32.62" resultid="100222" heatid="105272" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="100223" heatid="105300" lane="4" entrytime="00:02:30.00" />
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="100224" heatid="105329" lane="8" entrytime="00:01:13.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-08-01" firstname="Monika" gender="F" lastname="MACIĄG" nation="POL" swrid="4992938" athleteid="100231">
              <RESULTS>
                <RESULT eventid="98777" points="313" reactiontime="+92" swimtime="00:00:34.92" resultid="100232" heatid="105118" lane="8" entrytime="00:00:33.84" entrycourse="SCM" />
                <RESULT eventid="98863" points="307" swimtime="00:12:11.62" resultid="100233" heatid="105405" lane="1" entrytime="00:12:40.11" />
                <RESULT eventid="98907" points="277" swimtime="00:00:41.50" resultid="100234" heatid="105175" lane="6" entrytime="00:00:41.51" />
                <RESULT eventid="98972" status="DNS" swimtime="00:00:00.00" resultid="100235" heatid="105208" lane="4" entrytime="00:01:17.21" />
                <RESULT eventid="99314" points="288" reactiontime="+83" swimtime="00:01:28.00" resultid="100236" heatid="105279" lane="1" entrytime="00:01:27.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="291" reactiontime="+100" swimtime="00:02:50.42" resultid="100237" heatid="105291" lane="5" entrytime="00:02:54.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                    <SPLIT distance="100" swimtime="00:01:23.98" />
                    <SPLIT distance="150" swimtime="00:02:08.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="280" reactiontime="+87" swimtime="00:03:09.63" resultid="100238" heatid="105333" lane="4" entrytime="00:03:07.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.78" />
                    <SPLIT distance="100" swimtime="00:01:33.14" />
                    <SPLIT distance="150" swimtime="00:02:21.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="276" reactiontime="+107" swimtime="00:06:07.06" resultid="100239" heatid="106055" lane="3" entrytime="00:05:42.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.81" />
                    <SPLIT distance="100" swimtime="00:01:24.68" />
                    <SPLIT distance="150" swimtime="00:02:10.50" />
                    <SPLIT distance="200" swimtime="00:02:56.50" />
                    <SPLIT distance="250" swimtime="00:03:43.11" />
                    <SPLIT distance="300" swimtime="00:04:31.13" />
                    <SPLIT distance="350" swimtime="00:05:19.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-04-09" firstname="Zbigniew" gender="M" lastname="RAMOS" nation="POL" athleteid="100240">
              <RESULTS>
                <RESULT eventid="98798" points="328" reactiontime="+86" swimtime="00:00:30.31" resultid="100241" heatid="105132" lane="2" entrytime="00:00:30.90" />
                <RESULT eventid="98956" points="260" swimtime="00:03:18.84" resultid="100242" heatid="105200" lane="7" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.71" />
                    <SPLIT distance="100" swimtime="00:01:27.83" />
                    <SPLIT distance="150" swimtime="00:02:20.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="322" reactiontime="+86" swimtime="00:01:08.39" resultid="100243" heatid="105220" lane="8" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="318" reactiontime="+93" swimtime="00:01:25.60" resultid="100244" heatid="105253" lane="4" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="272" reactiontime="+84" swimtime="00:00:34.61" resultid="100245" heatid="105270" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="99361" reactiontime="+87" status="DNS" swimtime="00:00:00.00" resultid="100246" heatid="105327" lane="2" entrytime="00:01:28.00" />
                <RESULT eventid="99425" points="335" reactiontime="+91" swimtime="00:00:38.39" resultid="100247" heatid="105358" lane="3" entrytime="00:00:36.90" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99059" points="409" reactiontime="+77" swimtime="00:02:05.79" resultid="100254" heatid="105242" lane="7" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.33" />
                    <SPLIT distance="100" swimtime="00:01:06.23" />
                    <SPLIT distance="150" swimtime="00:01:38.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100151" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="100156" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="100218" number="3" reactiontime="+9" />
                    <RELAYPOSITION athleteid="100209" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" points="438" reactiontime="+78" swimtime="00:01:51.70" resultid="100256" heatid="105311" lane="2" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.59" />
                    <SPLIT distance="100" swimtime="00:00:55.79" />
                    <SPLIT distance="150" swimtime="00:01:23.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100156" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="100218" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="100209" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="100151" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="99059" points="322" reactiontime="+66" swimtime="00:02:16.27" resultid="100255" heatid="105241" lane="8" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                    <SPLIT distance="100" swimtime="00:01:12.35" />
                    <SPLIT distance="150" swimtime="00:01:45.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100204" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="100187" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="100240" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="100198" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" points="355" reactiontime="+95" swimtime="00:01:59.81" resultid="100257" heatid="105310" lane="3" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                    <SPLIT distance="100" swimtime="00:00:59.52" />
                    <SPLIT distance="150" swimtime="00:01:30.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100240" number="1" reactiontime="+95" />
                    <RELAYPOSITION athleteid="100187" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="100198" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="100204" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="99036" points="329" reactiontime="+74" swimtime="00:02:33.54" resultid="100252" heatid="105238" lane="8" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.98" />
                    <SPLIT distance="100" swimtime="00:01:20.43" />
                    <SPLIT distance="150" swimtime="00:01:59.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100163" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="100183" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="100177" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="100231" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99234" points="357" reactiontime="+77" swimtime="00:02:16.35" resultid="100253" heatid="105307" lane="1" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.98" />
                    <SPLIT distance="100" swimtime="00:01:08.33" />
                    <SPLIT distance="150" swimtime="00:01:44.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100163" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="100231" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="100171" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="100177" number="4" reactiontime="+74" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="279" reactiontime="+96" swimtime="00:02:09.72" resultid="100249" heatid="105160" lane="6" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                    <SPLIT distance="100" swimtime="00:01:05.16" />
                    <SPLIT distance="150" swimtime="00:01:40.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100231" number="1" reactiontime="+96" />
                    <RELAYPOSITION athleteid="100187" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="100171" number="3" reactiontime="+22" />
                    <RELAYPOSITION athleteid="100240" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="99441" points="337" reactiontime="+83" swimtime="00:02:14.21" resultid="100250" heatid="105365" lane="2" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.30" />
                    <SPLIT distance="100" swimtime="00:01:09.72" />
                    <SPLIT distance="150" swimtime="00:01:47.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100163" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="100156" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="100177" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="100209" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="98846" points="361" reactiontime="+90" swimtime="00:01:59.07" resultid="100248" heatid="105161" lane="8" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                    <SPLIT distance="100" swimtime="00:00:59.70" />
                    <SPLIT distance="150" swimtime="00:01:32.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100177" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="100209" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="100163" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="100156" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="99441" points="249" reactiontime="+91" swimtime="00:02:28.34" resultid="100251" heatid="105364" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.45" />
                    <SPLIT distance="100" swimtime="00:01:17.31" />
                    <SPLIT distance="150" swimtime="00:01:51.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100231" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="100187" number="2" reactiontime="+33" />
                    <RELAYPOSITION athleteid="100240" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="100171" number="4" reactiontime="+71" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="101502" name="UKS G-8 Bielany">
          <CONTACT name="Koszuta" phone="68345914" />
          <ATHLETES>
            <ATHLETE birthdate="1971-05-04" firstname="Wiater" gender="M" lastname="KRZYSTOF" nation="POL" athleteid="101503">
              <RESULTS>
                <RESULT eventid="98891" status="DNS" swimtime="00:00:00.00" resultid="104996" heatid="105422" lane="7" entrytime="00:22:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="MAL" clubid="100258" name="UKS SP 8 Chrzanów">
          <CONTACT city="Chrzanów" email="abalp@poczta.onet.pl" name="Zabrzański" phone="692076808" state="MAŁ" street="niepodległości 7/46" zip="32-500" />
          <ATHLETES>
            <ATHLETE birthdate="1954-05-12" firstname="Alfred" gender="M" lastname="ZABRZAŃSKI" nation="POL" swrid="4477631" athleteid="100268">
              <RESULTS>
                <RESULT eventid="98798" points="289" reactiontime="+92" swimtime="00:00:31.61" resultid="100269" heatid="105131" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="98891" status="DNS" swimtime="00:00:00.00" resultid="100270" heatid="105423" lane="0" entrytime="00:26:25.00" />
                <RESULT eventid="98924" points="194" reactiontime="+91" swimtime="00:00:41.50" resultid="100271" heatid="105184" lane="1" entrytime="00:00:41.00" />
                <RESULT eventid="98988" points="281" reactiontime="+99" swimtime="00:01:11.56" resultid="100272" heatid="105219" lane="0" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="225" reactiontime="+111" swimtime="00:02:47.60" resultid="100273" heatid="105298" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.49" />
                    <SPLIT distance="100" swimtime="00:01:19.40" />
                    <SPLIT distance="150" swimtime="00:02:03.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="100274" entrytime="00:06:03.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00111" nation="POL" region="SLA" clubid="100904" name="UKS TRÓJKA Częstochowa">
          <CONTACT city="Częstochowa" name="Gawda Jacek" phone="511181791" state="ŚL" zip="42-200" />
          <ATHLETES>
            <ATHLETE birthdate="1990-02-15" firstname="Manuela" gender="F" lastname="NAWROCKA" nation="POL" license="S00111100008" swrid="4806455" athleteid="100905">
              <RESULTS>
                <RESULT eventid="98814" points="403" reactiontime="+91" swimtime="00:02:50.70" resultid="100906" heatid="105147" lane="7" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                    <SPLIT distance="100" swimtime="00:01:19.61" />
                    <SPLIT distance="150" swimtime="00:02:10.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="388" reactiontime="+80" swimtime="00:00:37.07" resultid="100907" heatid="105177" lane="3" entrytime="00:00:36.50" />
                <RESULT eventid="98940" points="373" swimtime="00:03:13.16" resultid="100908" heatid="105194" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.22" />
                    <SPLIT distance="100" swimtime="00:01:31.05" />
                    <SPLIT distance="150" swimtime="00:02:21.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="389" reactiontime="+101" swimtime="00:01:28.13" resultid="100909" heatid="105247" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="332" reactiontime="+82" swimtime="00:01:23.90" resultid="100910" heatid="105280" lane="9" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="297" reactiontime="+94" swimtime="00:01:23.88" resultid="100911" heatid="105322" lane="4" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="367" reactiontime="+66" swimtime="00:00:41.17" resultid="100912" heatid="105349" lane="8" entrytime="00:00:39.80" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="UKS3" nation="POL" region="WIE" clubid="100082" name="UKS Trójka Oborniki">
          <CONTACT city="Oborniki" email="janwol@poczta.onet.pl" name="Wolniewicz" phone="791064667" state="WIE" street="Piłsudskiego 49/42" zip="64-600" />
          <ATHLETES>
            <ATHLETE birthdate="1948-12-22" firstname="Janusz" gender="M" lastname="WOLNIEWICZ" nation="POL" swrid="4754624" athleteid="100083">
              <RESULTS>
                <RESULT eventid="98798" points="197" reactiontime="+85" swimtime="00:00:35.93" resultid="100084" heatid="105127" lane="7" entrytime="00:00:35.08" entrycourse="SCM" />
                <RESULT eventid="98891" points="132" swimtime="00:28:27.26" resultid="100085" heatid="105424" lane="0" entrytime="00:28:22.00" entrycourse="SCM" />
                <RESULT eventid="98988" points="173" reactiontime="+96" swimtime="00:01:24.06" resultid="100086" heatid="105215" lane="4" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="100087" heatid="105266" lane="8" entrytime="00:00:46.00" entrycourse="SCM" />
                <RESULT eventid="99218" points="112" reactiontime="+112" swimtime="00:03:31.46" resultid="100088" heatid="105296" lane="3" entrytime="00:03:16.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.02" />
                    <SPLIT distance="100" swimtime="00:01:42.92" />
                    <SPLIT distance="150" swimtime="00:02:40.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="123" reactiontime="+98" swimtime="00:07:22.40" resultid="100089" heatid="106066" lane="5" entrytime="00:07:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.67" />
                    <SPLIT distance="100" swimtime="00:01:38.96" />
                    <SPLIT distance="150" swimtime="00:02:34.17" />
                    <SPLIT distance="200" swimtime="00:03:30.52" />
                    <SPLIT distance="250" swimtime="00:04:28.78" />
                    <SPLIT distance="300" swimtime="00:05:27.43" />
                    <SPLIT distance="350" swimtime="00:06:26.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WODKAT" nation="POL" region="SLA" clubid="102257" name="UKS Wodnik 29 Katowice">
          <CONTACT name="Skoczylas" phone="662297707" />
          <ATHLETES>
            <ATHLETE birthdate="1958-03-01" firstname="Jan" gender="M" lastname="WILCZEK" nation="POL" swrid="4992641" athleteid="102258">
              <RESULTS>
                <RESULT eventid="98798" points="360" reactiontime="+102" swimtime="00:00:29.38" resultid="102259" heatid="105135" lane="2" entrytime="00:00:29.40" />
                <RESULT eventid="98988" points="295" reactiontime="+96" swimtime="00:01:10.41" resultid="102260" heatid="105220" lane="4" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="343" reactiontime="+98" swimtime="00:00:32.03" resultid="102261" heatid="105271" lane="4" entrytime="00:00:31.40" />
                <RESULT eventid="99361" points="288" reactiontime="+94" swimtime="00:01:15.42" resultid="102262" heatid="105329" lane="9" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-28" firstname="Jerzy" gender="M" lastname="MROZIŃSKI" nation="POL" swrid="4877351" athleteid="102263">
              <RESULTS>
                <RESULT eventid="98798" points="289" reactiontime="+91" swimtime="00:00:31.60" resultid="102264" heatid="105132" lane="1" entrytime="00:00:31.00" />
                <RESULT comment="Rekord Polski Masters" eventid="98956" points="300" reactiontime="+84" swimtime="00:03:09.56" resultid="102265" heatid="105201" lane="8" entrytime="00:03:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.76" />
                    <SPLIT distance="100" swimtime="00:01:29.91" />
                    <SPLIT distance="150" swimtime="00:02:19.69" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99091" points="339" reactiontime="+97" swimtime="00:01:23.76" resultid="102266" heatid="105254" lane="2" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="102267" heatid="105298" lane="5" entrytime="00:02:45.00" />
                <RESULT comment="Rekord Polski Masters" eventid="99425" points="403" reactiontime="+77" swimtime="00:00:36.09" resultid="102268" heatid="105359" lane="7" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-26" firstname="Piotr" gender="M" lastname="KLEPACKI" nation="POL" swrid="4992638" athleteid="102269">
              <RESULTS>
                <RESULT eventid="98798" points="240" swimtime="00:00:33.64" resultid="102270" heatid="105125" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="98924" points="134" reactiontime="+68" swimtime="00:00:46.89" resultid="102271" heatid="105180" lane="5" entrytime="00:00:59.00" />
                <RESULT eventid="98988" points="167" reactiontime="+86" swimtime="00:01:25.16" resultid="102272" heatid="105214" lane="7" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="105086" heatid="105351" lane="5" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-12-05" firstname="Marcin" gender="M" lastname="SZCZYPIŃSKI" nation="POL" swrid="4060998" athleteid="102274">
              <RESULTS>
                <RESULT eventid="98798" points="578" reactiontime="+83" swimtime="00:00:25.10" resultid="102275" heatid="105143" lane="0" entrytime="00:00:25.00" />
                <RESULT comment="Rekord Polski Masters, Rekord Polski Masters" eventid="98891" points="509" swimtime="00:18:10.62" resultid="102276" heatid="105420" lane="3" entrytime="00:18:45.00" />
                <RESULT eventid="98924" points="498" reactiontime="+82" swimtime="00:00:30.31" resultid="102277" heatid="105190" lane="1" entrytime="00:00:29.70" />
                <RESULT eventid="98988" points="632" reactiontime="+83" swimtime="00:00:54.65" resultid="102278" heatid="105228" lane="1" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="591" reactiontime="+78" swimtime="00:00:26.72" resultid="102279" heatid="105276" lane="8" entrytime="00:00:27.00" />
                <RESULT eventid="99218" points="531" reactiontime="+79" swimtime="00:02:05.92" resultid="102280" heatid="105305" lane="8" entrytime="00:02:08.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.71" />
                    <SPLIT distance="100" swimtime="00:01:02.50" />
                    <SPLIT distance="150" swimtime="00:01:34.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="612" reactiontime="+83" swimtime="00:00:58.67" resultid="102281" heatid="105331" lane="6" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.51" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99473" points="557" reactiontime="+82" swimtime="00:04:27.47" resultid="102282" heatid="106059" lane="7" entrytime="00:04:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.33" />
                    <SPLIT distance="100" swimtime="00:01:01.84" />
                    <SPLIT distance="150" swimtime="00:01:35.92" />
                    <SPLIT distance="200" swimtime="00:02:10.70" />
                    <SPLIT distance="250" swimtime="00:02:46.04" />
                    <SPLIT distance="300" swimtime="00:03:21.00" />
                    <SPLIT distance="350" swimtime="00:03:55.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-07-10" firstname="Sandra" gender="F" lastname="PIETRZAK" nation="POL" swrid="4061017" athleteid="102283">
              <RESULTS>
                <RESULT eventid="98777" points="509" reactiontime="+79" swimtime="00:00:29.72" resultid="102284" heatid="105120" lane="6" entrytime="00:00:29.99" entrycourse="LCM" />
                <RESULT comment="Rekord Polski Masters" eventid="98863" points="514" reactiontime="+64" swimtime="00:10:16.22" resultid="102285" heatid="105404" lane="8" entrytime="00:11:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                    <SPLIT distance="100" swimtime="00:01:10.58" />
                    <SPLIT distance="150" swimtime="00:01:48.36" />
                    <SPLIT distance="200" swimtime="00:02:26.65" />
                    <SPLIT distance="250" swimtime="00:03:05.14" />
                    <SPLIT distance="300" swimtime="00:03:43.68" />
                    <SPLIT distance="350" swimtime="00:04:22.97" />
                    <SPLIT distance="400" swimtime="00:05:02.27" />
                    <SPLIT distance="450" swimtime="00:05:41.52" />
                    <SPLIT distance="500" swimtime="00:06:21.25" />
                    <SPLIT distance="550" swimtime="00:07:00.93" />
                    <SPLIT distance="600" swimtime="00:07:40.36" />
                    <SPLIT distance="650" swimtime="00:08:19.67" />
                    <SPLIT distance="700" swimtime="00:08:59.33" />
                    <SPLIT distance="750" swimtime="00:09:37.66" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="98972" points="558" reactiontime="+87" swimtime="00:01:03.23" resultid="102286" heatid="105211" lane="5" entrytime="00:01:06.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="528" reactiontime="+89" swimtime="00:02:19.78" resultid="102287" heatid="105294" lane="0" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                    <SPLIT distance="100" swimtime="00:01:07.22" />
                    <SPLIT distance="150" swimtime="00:01:43.57" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99457" points="524" reactiontime="+91" swimtime="00:04:56.55" resultid="102288" heatid="106054" lane="0" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                    <SPLIT distance="100" swimtime="00:01:09.30" />
                    <SPLIT distance="150" swimtime="00:01:46.06" />
                    <SPLIT distance="200" swimtime="00:02:23.29" />
                    <SPLIT distance="250" swimtime="00:03:01.35" />
                    <SPLIT distance="300" swimtime="00:03:39.59" />
                    <SPLIT distance="350" swimtime="00:04:18.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-15" firstname="Anna" gender="F" lastname="DUDA" nation="POL" swrid="4992966" athleteid="102289">
              <RESULTS>
                <RESULT eventid="98777" points="457" reactiontime="+87" swimtime="00:00:30.80" resultid="102290" heatid="105120" lane="3" entrytime="00:00:29.84" entrycourse="SCM" />
                <RESULT eventid="98972" points="416" reactiontime="+83" swimtime="00:01:09.71" resultid="102291" heatid="105211" lane="4" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="475" reactiontime="+92" swimtime="00:00:32.12" resultid="102292" heatid="105264" lane="1" entrytime="00:00:31.40" />
                <RESULT eventid="99344" status="DNS" swimtime="00:00:00.00" resultid="102293" heatid="105323" lane="7" entrytime="00:01:16.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="99059" points="351" reactiontime="+70" swimtime="00:02:12.42" resultid="102295" heatid="105240" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.72" />
                    <SPLIT distance="100" swimtime="00:01:07.89" />
                    <SPLIT distance="150" swimtime="00:01:39.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102274" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="102263" number="2" reactiontime="+65" />
                    <RELAYPOSITION athleteid="102258" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="102269" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" status="DNS" swimtime="00:00:00.00" resultid="102296" heatid="105309" lane="6" entrytime="00:02:15.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102258" number="1" />
                    <RELAYPOSITION athleteid="102269" number="2" />
                    <RELAYPOSITION athleteid="102263" number="3" />
                    <RELAYPOSITION athleteid="102274" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski Masters" eventid="98846" points="413" reactiontime="+86" swimtime="00:01:53.87" resultid="102294" heatid="105161" lane="2" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.43" />
                    <SPLIT distance="100" swimtime="00:01:00.24" />
                    <SPLIT distance="150" swimtime="00:01:29.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="102283" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="102289" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="102258" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="102274" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="031/05" nation="POL" region="LOD" clubid="100562" name="UTW Masters Zgierz">
          <CONTACT city="ZGIERZ" internet="roman.wiczel@gmail.com" name="WICZEL" phone="691-928-922" state="ŁÓDZK" street="ŁĘCZYCKA 24" zip="95-100" />
          <ATHLETES>
            <ATHLETE birthdate="1948-01-22" firstname="Roman" gender="M" lastname="WICZEL" nation="POL" license="503105200002" swrid="4876444" athleteid="100563">
              <RESULTS>
                <RESULT eventid="98798" points="182" reactiontime="+95" swimtime="00:00:36.87" resultid="100564" heatid="105126" lane="5" entrytime="00:00:36.00" entrycourse="LCM" />
                <RESULT eventid="98956" points="242" reactiontime="+114" swimtime="00:03:23.66" resultid="100565" heatid="105199" lane="5" entrytime="00:03:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.19" />
                    <SPLIT distance="100" swimtime="00:01:38.22" />
                    <SPLIT distance="150" swimtime="00:02:31.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="267" reactiontime="+100" swimtime="00:01:30.71" resultid="100566" heatid="105252" lane="6" entrytime="00:01:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="307" reactiontime="+106" swimtime="00:00:39.52" resultid="100567" heatid="105356" lane="3" entrytime="00:00:40.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-02-07" firstname="Krzysztof" gender="M" lastname="WOJCIECHOWSKI" nation="POL" license="503105200008" athleteid="100568">
              <RESULTS>
                <RESULT eventid="98798" points="209" reactiontime="+114" swimtime="00:00:35.19" resultid="100569" heatid="105126" lane="0" entrytime="00:00:37.00" entrycourse="LCM" />
                <RESULT eventid="99091" points="224" reactiontime="+115" swimtime="00:01:36.13" resultid="100570" heatid="105252" lane="0" entrytime="00:01:33.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="270" reactiontime="+114" swimtime="00:00:41.24" resultid="100571" heatid="105355" lane="0" entrytime="00:00:42.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-12-03" firstname="Zbigniew" gender="M" lastname="MACIEJCZYK" nation="POL" license="503105200001" swrid="4302705" athleteid="100572">
              <RESULTS>
                <RESULT eventid="98798" points="246" reactiontime="+103" swimtime="00:00:33.33" resultid="100573" heatid="105127" lane="3" entrytime="00:00:35.00" entrycourse="LCM" />
                <RESULT eventid="98988" points="221" reactiontime="+107" swimtime="00:01:17.54" resultid="100574" heatid="105216" lane="1" entrytime="00:01:17.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" status="DNS" swimtime="00:00:00.00" resultid="100575" heatid="105232" lane="5" entrytime="00:04:10.00" entrycourse="LCM" />
                <RESULT eventid="99170" points="208" reactiontime="+101" swimtime="00:00:37.82" resultid="100576" heatid="105268" lane="9" entrytime="00:00:37.00" entrycourse="LCM" />
                <RESULT eventid="99361" points="118" reactiontime="+110" swimtime="00:01:41.42" resultid="100577" heatid="105326" lane="0" entrytime="00:01:47.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-10-03" firstname="Agata" gender="F" lastname="GŁOWACKA" nation="POL" license="503105100007" athleteid="100578">
              <RESULTS>
                <RESULT eventid="98777" points="233" reactiontime="+147" swimtime="00:00:38.56" resultid="100579" heatid="105119" lane="0" entrytime="00:00:32.00" />
                <RESULT eventid="98814" points="152" reactiontime="+129" swimtime="00:03:56.12" resultid="100580" heatid="105146" lane="2" entrytime="00:03:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.38" />
                    <SPLIT distance="100" swimtime="00:01:47.24" />
                    <SPLIT distance="150" swimtime="00:03:00.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="233" reactiontime="+88" swimtime="00:00:43.92" resultid="100581" heatid="105176" lane="4" entrytime="00:00:39.00" entrycourse="LCM" />
                <RESULT eventid="98972" status="DNS" swimtime="00:00:00.00" resultid="100582" heatid="105210" lane="7" entrytime="00:01:12.00" entrycourse="LCM" />
                <RESULT eventid="99154" status="DNS" swimtime="00:00:00.00" resultid="100583" heatid="105260" lane="3" entrytime="00:00:40.00" entrycourse="LCM" />
                <RESULT eventid="99314" points="186" reactiontime="+100" swimtime="00:01:41.70" resultid="100584" heatid="105278" lane="4" entrytime="00:01:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="163" reactiontime="+106" swimtime="00:03:26.58" resultid="100585" heatid="105293" lane="6" entrytime="00:02:35.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.29" />
                    <SPLIT distance="100" swimtime="00:01:33.27" />
                    <SPLIT distance="150" swimtime="00:02:29.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-03" firstname="Urszula" gender="F" lastname="MRÓZ" nation="POL" license="503105100003" swrid="4754660" athleteid="100586">
              <RESULTS>
                <RESULT eventid="98777" points="301" reactiontime="+103" swimtime="00:00:35.40" resultid="100587" heatid="105117" lane="4" entrytime="00:00:34.17" entrycourse="LCM" />
                <RESULT eventid="98907" points="295" reactiontime="+83" swimtime="00:00:40.64" resultid="100588" heatid="105176" lane="7" entrytime="00:00:39.20" entrycourse="LCM" />
                <RESULT eventid="98972" status="DNS" swimtime="00:00:00.00" resultid="100589" heatid="105209" lane="6" entrytime="00:01:15.00" entrycourse="LCM" />
                <RESULT eventid="99154" points="283" reactiontime="+103" swimtime="00:00:38.18" resultid="100590" heatid="105262" lane="1" entrytime="00:00:37.00" entrycourse="LCM" />
                <RESULT eventid="99314" points="220" reactiontime="+83" swimtime="00:01:36.18" resultid="100591" heatid="105279" lane="0" entrytime="00:01:28.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="209" reactiontime="+99" swimtime="00:01:34.24" resultid="100592" heatid="105322" lane="3" entrytime="00:01:27.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="204" reactiontime="+82" swimtime="00:03:30.66" resultid="100593" heatid="105334" lane="7" entrytime="00:03:02.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.63" />
                    <SPLIT distance="100" swimtime="00:01:44.36" />
                    <SPLIT distance="150" swimtime="00:02:39.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-09-03" firstname="Arkadiusz" gender="M" lastname="BILSKI" nation="POL" license="503105200013" athleteid="100594">
              <RESULTS>
                <RESULT eventid="98830" points="347" reactiontime="+84" swimtime="00:02:42.08" resultid="100595" heatid="105157" lane="6" entrytime="00:02:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.78" />
                    <SPLIT distance="100" swimtime="00:01:16.11" />
                    <SPLIT distance="150" swimtime="00:02:01.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="416" reactiontime="+92" swimtime="00:02:50.10" resultid="100596" heatid="105204" lane="0" entrytime="00:02:44.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.37" />
                    <SPLIT distance="100" swimtime="00:01:20.11" />
                    <SPLIT distance="150" swimtime="00:02:04.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="447" reactiontime="+76" swimtime="00:01:16.43" resultid="100597" heatid="105258" lane="9" entrytime="00:01:13.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="450" reactiontime="+78" swimtime="00:00:34.78" resultid="100598" heatid="105362" lane="0" entrytime="00:00:32.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-05-12" firstname="Tadeusz" gender="M" lastname="OBIEDZIŃSKI" nation="POL" license="503105200011" swrid="4992722" athleteid="100599">
              <RESULTS>
                <RESULT eventid="98830" points="118" reactiontime="+102" swimtime="00:03:52.12" resultid="100600" heatid="105150" lane="3" entrytime="00:03:40.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.20" />
                    <SPLIT distance="100" swimtime="00:01:48.19" />
                    <SPLIT distance="150" swimtime="00:02:50.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="159" reactiontime="+115" swimtime="00:03:54.00" resultid="100601" heatid="105198" lane="3" entrytime="00:03:43.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.37" />
                    <SPLIT distance="100" swimtime="00:01:46.62" />
                    <SPLIT distance="150" swimtime="00:02:49.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" status="DNS" swimtime="00:00:00.00" resultid="100602" heatid="105233" lane="6" entrytime="00:03:43.83" entrycourse="LCM" />
                <RESULT eventid="99091" points="195" reactiontime="+103" swimtime="00:01:40.67" resultid="100603" heatid="105252" lane="9" entrytime="00:01:34.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="100604" heatid="105267" lane="7" entrytime="00:00:39.98" entrycourse="LCM" />
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="100605" heatid="105326" lane="7" entrytime="00:01:42.63" entrycourse="LCM" />
                <RESULT eventid="99425" points="250" reactiontime="+104" swimtime="00:00:42.31" resultid="100606" heatid="105356" lane="0" entrytime="00:00:40.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-12" firstname="Małgorzata" gender="F" lastname="ŚCIBIOREK" nation="POL" license="503105100005" swrid="4992745" athleteid="100607">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski Masters" eventid="98814" points="462" reactiontime="+88" swimtime="00:02:43.18" resultid="100608" heatid="105147" lane="5" entrytime="00:02:41.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                    <SPLIT distance="100" swimtime="00:01:15.62" />
                    <SPLIT distance="150" swimtime="00:02:03.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="378" reactiontime="+77" swimtime="00:00:37.42" resultid="100609" heatid="105178" lane="8" entrytime="00:00:35.00" entrycourse="LCM" />
                <RESULT eventid="99004" points="343" reactiontime="+95" swimtime="00:02:53.94" resultid="100610" heatid="105230" lane="4" entrytime="00:02:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                    <SPLIT distance="100" swimtime="00:01:14.01" />
                    <SPLIT distance="150" swimtime="00:01:59.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="476" reactiontime="+85" swimtime="00:00:32.10" resultid="100611" heatid="105264" lane="8" entrytime="00:00:31.50" entrycourse="LCM" />
                <RESULT comment="Rekord Polski Masters" eventid="99314" points="399" reactiontime="+84" swimtime="00:01:18.94" resultid="100612" heatid="105280" lane="3" entrytime="00:01:13.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.51" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99344" points="498" reactiontime="+95" swimtime="00:01:10.62" resultid="100613" heatid="105323" lane="3" entrytime="00:01:12.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1922-01-04" firstname="Kazimierz" gender="M" lastname="MRÓWCZYŃSKI" nation="POL" license="503105200015" swrid="4302706" athleteid="100614">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski Masters" eventid="98798" points="33" reactiontime="+107" swimtime="00:01:05.04" resultid="100615" heatid="105124" lane="9" entrytime="00:00:55.00" entrycourse="LCM" />
                <RESULT comment="Rekord Polski Masters" eventid="98988" points="29" reactiontime="+133" swimtime="00:02:31.56" resultid="100616" heatid="105213" lane="2" entrytime="00:02:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.39" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99218" points="29" reactiontime="+134" swimtime="00:05:30.88" resultid="100617" heatid="105295" lane="1" entrytime="00:04:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.55" />
                    <SPLIT distance="100" swimtime="00:02:43.00" />
                    <SPLIT distance="150" swimtime="00:04:09.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="100618" entrytime="00:10:00.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-09" firstname="Włodzimierz" gender="M" lastname="PRZYTULSKI" nation="POL" license="503105200006" swrid="4754657" athleteid="100619">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="100620" heatid="105133" lane="3" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT eventid="98830" points="292" reactiontime="+90" swimtime="00:02:51.73" resultid="100621" heatid="105153" lane="1" entrytime="00:02:57.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                    <SPLIT distance="100" swimtime="00:01:18.54" />
                    <SPLIT distance="150" swimtime="00:02:12.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="309" reactiontime="+91" swimtime="00:00:35.53" resultid="100622" heatid="105186" lane="2" entrytime="00:00:36.00" entrycourse="LCM" />
                <RESULT eventid="98988" points="354" reactiontime="+83" swimtime="00:01:06.28" resultid="100623" heatid="105221" lane="7" entrytime="00:01:07.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="270" reactiontime="+72" swimtime="00:01:20.31" resultid="100624" heatid="105284" lane="6" entrytime="00:01:19.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="100625" heatid="105300" lane="8" entrytime="00:02:32.00" entrycourse="LCM" />
                <RESULT eventid="99361" points="270" reactiontime="+93" swimtime="00:01:17.01" resultid="100626" heatid="105328" lane="5" entrytime="00:01:18.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="100627" heatid="105339" lane="4" entrytime="00:02:58.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-07" firstname="Ewa" gender="F" lastname="STĘPIEŃ" nation="POL" license="503105100004" swrid="4876443" athleteid="100628">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski Masters" eventid="98777" points="395" reactiontime="+66" swimtime="00:00:32.34" resultid="100629" heatid="105119" lane="7" entrytime="00:00:31.81" entrycourse="SCM" />
                <RESULT eventid="98972" points="343" reactiontime="+82" swimtime="00:01:14.33" resultid="100630" heatid="105209" lane="3" entrytime="00:01:14.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="382" reactiontime="+72" swimtime="00:01:28.68" resultid="100631" heatid="105247" lane="8" entrytime="00:01:29.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" status="DNS" swimtime="00:00:00.00" resultid="100632" heatid="105291" lane="6" entrytime="00:02:56.00" entrycourse="LCM" />
                <RESULT eventid="99409" points="392" swimtime="00:00:40.27" resultid="100633" heatid="105349" lane="1" entrytime="00:00:39.80" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="99059" points="245" reactiontime="+83" swimtime="00:02:29.24" resultid="100640" heatid="105240" lane="5" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                    <SPLIT distance="100" swimtime="00:01:16.07" />
                    <SPLIT distance="150" swimtime="00:01:55.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100619" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="100563" number="2" reactiontime="+28" />
                    <RELAYPOSITION athleteid="100572" number="3" reactiontime="+86" />
                    <RELAYPOSITION athleteid="100568" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" points="247" reactiontime="+111" swimtime="00:02:15.20" resultid="100641" heatid="105309" lane="2" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                    <SPLIT distance="100" swimtime="00:01:10.35" />
                    <SPLIT distance="150" swimtime="00:01:45.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100572" number="1" reactiontime="+111" />
                    <RELAYPOSITION athleteid="100599" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="100568" number="3" reactiontime="+62" />
                    <RELAYPOSITION athleteid="100619" number="4" reactiontime="+79" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="99036" points="334" reactiontime="+81" swimtime="00:02:32.74" resultid="100638" heatid="105238" lane="5" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.56" />
                    <SPLIT distance="100" swimtime="00:01:21.88" />
                    <SPLIT distance="150" swimtime="00:01:55.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100586" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="100628" number="2" reactiontime="+38" />
                    <RELAYPOSITION athleteid="100607" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="100578" number="4" reactiontime="+62" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99234" points="348" reactiontime="+95" swimtime="00:02:17.50" resultid="100639" heatid="105307" lane="6" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.33" />
                    <SPLIT distance="100" swimtime="00:01:12.93" />
                    <SPLIT distance="150" swimtime="00:01:45.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100586" number="1" reactiontime="+95" />
                    <RELAYPOSITION athleteid="100578" number="2" reactiontime="+84" />
                    <RELAYPOSITION athleteid="100628" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="100607" number="4" reactiontime="+62" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="318" reactiontime="+89" swimtime="00:02:04.28" resultid="100634" heatid="105161" lane="7" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                    <SPLIT distance="100" swimtime="00:01:00.93" />
                    <SPLIT distance="150" swimtime="00:01:33.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100607" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="100594" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="100628" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="100619" number="4" reactiontime="+69" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99441" points="330" reactiontime="+82" swimtime="00:02:15.19" resultid="100635" heatid="105365" lane="3" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                    <SPLIT distance="100" swimtime="00:01:10.64" />
                    <SPLIT distance="150" swimtime="00:01:42.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100619" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="100594" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="100607" number="3" reactiontime="+64" />
                    <RELAYPOSITION athleteid="100628" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="98846" points="224" reactiontime="+103" swimtime="00:02:19.62" resultid="100636" heatid="105160" lane="7" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                    <SPLIT distance="100" swimtime="00:01:08.16" />
                    <SPLIT distance="150" swimtime="00:01:42.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100572" number="1" reactiontime="+103" />
                    <RELAYPOSITION athleteid="100586" number="2" reactiontime="+85" />
                    <RELAYPOSITION athleteid="100568" number="3" reactiontime="+60" />
                    <RELAYPOSITION athleteid="100578" number="4" reactiontime="+78" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" points="206" reactiontime="+95" swimtime="00:02:37.99" resultid="100637" heatid="105364" lane="2" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.09" />
                    <SPLIT distance="100" swimtime="00:01:20.96" />
                    <SPLIT distance="150" swimtime="00:02:01.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100586" number="1" reactiontime="+95" />
                    <RELAYPOSITION athleteid="100563" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="100572" number="3" reactiontime="+88" />
                    <RELAYPOSITION athleteid="100578" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="UKR" clubid="101176" name="Ukraina">
          <CONTACT name="Lysenko" />
          <ATHLETES>
            <ATHLETE birthdate="1973-03-22" firstname="Andrii" gender="M" lastname="LYSENKO" nation="UKR" swrid="4776565" athleteid="101177">
              <RESULTS>
                <RESULT eventid="98830" points="409" reactiontime="+96" swimtime="00:02:33.50" resultid="101178" heatid="105157" lane="1" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                    <SPLIT distance="100" swimtime="00:01:12.11" />
                    <SPLIT distance="150" swimtime="00:01:57.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="390" reactiontime="+86" swimtime="00:00:32.90" resultid="101179" heatid="105189" lane="0" entrytime="00:00:32.00" />
                <RESULT eventid="98988" points="462" reactiontime="+99" swimtime="00:01:00.65" resultid="101180" heatid="105225" lane="2" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="425" reactiontime="+75" swimtime="00:01:09.06" resultid="101181" heatid="105286" lane="4" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="372" reactiontime="+106" swimtime="00:05:38.89" resultid="101182" heatid="106053" lane="0" entrytime="00:05:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                    <SPLIT distance="100" swimtime="00:01:16.00" />
                    <SPLIT distance="150" swimtime="00:01:59.68" />
                    <SPLIT distance="200" swimtime="00:02:43.18" />
                    <SPLIT distance="250" swimtime="00:03:31.73" />
                    <SPLIT distance="300" swimtime="00:04:20.93" />
                    <SPLIT distance="350" swimtime="00:05:00.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="394" reactiontime="+95" swimtime="00:02:32.64" resultid="101183" heatid="105342" lane="1" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.09" />
                    <SPLIT distance="100" swimtime="00:01:14.68" />
                    <SPLIT distance="150" swimtime="00:01:53.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="357" reactiontime="+96" swimtime="00:05:10.18" resultid="101184" heatid="106061" lane="2" entrytime="00:04:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                    <SPLIT distance="100" swimtime="00:01:15.20" />
                    <SPLIT distance="150" swimtime="00:01:54.84" />
                    <SPLIT distance="200" swimtime="00:02:34.79" />
                    <SPLIT distance="250" swimtime="00:03:13.26" />
                    <SPLIT distance="300" swimtime="00:03:53.07" />
                    <SPLIT distance="350" swimtime="00:04:32.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-05-05" firstname="Sergii" gender="M" lastname="BABKIN" nation="UKR" swrid="4776556" athleteid="101185">
              <RESULTS>
                <RESULT eventid="98798" points="454" reactiontime="+75" swimtime="00:00:27.20" resultid="101186" heatid="105140" lane="6" entrytime="00:00:27.00" />
                <RESULT eventid="98830" points="433" reactiontime="+82" swimtime="00:02:30.68" resultid="101187" heatid="105157" lane="0" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                    <SPLIT distance="100" swimtime="00:01:10.59" />
                    <SPLIT distance="150" swimtime="00:01:55.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="513" reactiontime="+74" swimtime="00:00:30.02" resultid="101188" heatid="105189" lane="3" entrytime="00:00:30.50" />
                <RESULT eventid="98988" points="481" reactiontime="+75" swimtime="00:00:59.86" resultid="101189" heatid="105225" lane="3" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="468" reactiontime="+76" swimtime="00:01:06.88" resultid="101190" heatid="105288" lane="0" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="424" reactiontime="+75" swimtime="00:02:15.74" resultid="101191" heatid="105304" lane="9" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                    <SPLIT distance="100" swimtime="00:01:08.87" />
                    <SPLIT distance="150" swimtime="00:01:43.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="425" reactiontime="+76" swimtime="00:02:28.77" resultid="101192" heatid="105342" lane="6" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.89" />
                    <SPLIT distance="100" swimtime="00:01:12.72" />
                    <SPLIT distance="150" swimtime="00:01:51.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="101193" entrytime="00:04:58.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-06-12" firstname="Andryi" gender="M" lastname="KHOMENKO" nation="UKR" swrid="4776894" athleteid="101194">
              <RESULTS>
                <RESULT eventid="98830" points="357" reactiontime="+87" swimtime="00:02:40.60" resultid="101195" heatid="105156" lane="9" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                    <SPLIT distance="100" swimtime="00:01:14.08" />
                    <SPLIT distance="150" swimtime="00:02:03.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="345" reactiontime="+79" swimtime="00:00:34.27" resultid="101196" heatid="105189" lane="8" entrytime="00:00:32.00" />
                <RESULT eventid="99186" points="345" reactiontime="+75" swimtime="00:01:13.99" resultid="101197" heatid="105287" lane="9" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="311" reactiontime="+98" swimtime="00:05:59.73" resultid="101198" heatid="106052" lane="6" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                    <SPLIT distance="100" swimtime="00:01:16.86" />
                    <SPLIT distance="150" swimtime="00:02:04.92" />
                    <SPLIT distance="200" swimtime="00:02:52.07" />
                    <SPLIT distance="250" swimtime="00:03:45.93" />
                    <SPLIT distance="300" swimtime="00:04:40.54" />
                    <SPLIT distance="350" swimtime="00:05:21.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="294" reactiontime="+89" swimtime="00:02:48.24" resultid="101199" heatid="105341" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                    <SPLIT distance="100" swimtime="00:01:22.88" />
                    <SPLIT distance="150" swimtime="00:02:07.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="101200" heatid="106061" lane="9" entrytime="00:05:01.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="URWAR" nation="POL" region="WAR" clubid="102495" name="Ursynów Masters">
          <CONTACT city="WARSZAWA" name="MICHAŁ NOWAK" />
          <ATHLETES>
            <ATHLETE birthdate="1985-05-26" firstname="Urszula" gender="F" lastname="GRYCZ" nation="POL" swrid="4992646" athleteid="102496">
              <RESULTS>
                <RESULT eventid="98863" points="254" swimtime="00:12:59.00" resultid="102497" heatid="105405" lane="7" entrytime="00:12:40.00" />
                <RESULT eventid="98972" points="321" reactiontime="+91" swimtime="00:01:16.03" resultid="102498" heatid="105209" lane="4" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="278" reactiontime="+89" swimtime="00:01:38.48" resultid="102499" heatid="105246" lane="8" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="275" reactiontime="+95" swimtime="00:02:53.65" resultid="102500" heatid="105291" lane="4" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.70" />
                    <SPLIT distance="100" swimtime="00:01:23.78" />
                    <SPLIT distance="150" swimtime="00:02:09.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="285" reactiontime="+96" swimtime="00:00:44.75" resultid="102501" heatid="105347" lane="0" entrytime="00:00:45.00" />
                <RESULT eventid="99457" points="272" reactiontime="+101" swimtime="00:06:09.07" resultid="102502" heatid="106055" lane="1" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.68" />
                    <SPLIT distance="100" swimtime="00:01:24.74" />
                    <SPLIT distance="150" swimtime="00:02:10.95" />
                    <SPLIT distance="200" swimtime="00:02:57.81" />
                    <SPLIT distance="250" swimtime="00:03:45.46" />
                    <SPLIT distance="300" swimtime="00:04:33.90" />
                    <SPLIT distance="350" swimtime="00:05:22.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-12-17" firstname="Michał" gender="M" lastname="NOWAK" nation="POL" swrid="4302652" athleteid="102503">
              <RESULTS>
                <RESULT eventid="98830" points="211" reactiontime="+98" swimtime="00:03:11.34" resultid="102504" heatid="105152" lane="0" entrytime="00:03:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.11" />
                    <SPLIT distance="100" swimtime="00:01:35.09" />
                    <SPLIT distance="150" swimtime="00:02:27.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="251" reactiontime="+93" swimtime="00:03:21.09" resultid="102505" heatid="105200" lane="3" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.65" />
                    <SPLIT distance="100" swimtime="00:01:37.39" />
                    <SPLIT distance="150" swimtime="00:02:29.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="294" reactiontime="+88" swimtime="00:01:27.82" resultid="102506" heatid="105253" lane="2" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="175" reactiontime="+80" swimtime="00:07:15.23" resultid="102507" heatid="106050" lane="8" entrytime="00:06:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.06" />
                    <SPLIT distance="100" swimtime="00:01:48.73" />
                    <SPLIT distance="150" swimtime="00:04:42.59" />
                    <SPLIT distance="200" swimtime="00:03:45.19" />
                    <SPLIT distance="300" swimtime="00:05:40.75" />
                    <SPLIT distance="350" swimtime="00:06:29.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="340" reactiontime="+85" swimtime="00:00:38.20" resultid="102508" heatid="105357" lane="5" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-01-23" firstname="Michał" gender="M" lastname="RYBARCZYK" nation="POL" swrid="4992648" athleteid="102509">
              <RESULTS>
                <RESULT eventid="98798" points="343" reactiontime="+87" swimtime="00:00:29.87" resultid="102510" heatid="105135" lane="5" entrytime="00:00:29.30" />
                <RESULT eventid="98924" points="95" reactiontime="+86" swimtime="00:00:52.68" resultid="102511" heatid="105184" lane="9" entrytime="00:00:42.00" />
                <RESULT eventid="98988" points="310" reactiontime="+84" swimtime="00:01:09.24" resultid="102512" heatid="105221" lane="4" entrytime="00:01:05.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="306" reactiontime="+85" swimtime="00:00:33.26" resultid="102513" heatid="105270" lane="4" entrytime="00:00:33.50" />
                <RESULT eventid="99218" points="287" reactiontime="+89" swimtime="00:02:34.54" resultid="102514" heatid="105300" lane="1" entrytime="00:02:31.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                    <SPLIT distance="100" swimtime="00:01:12.55" />
                    <SPLIT distance="150" swimtime="00:01:53.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="213" reactiontime="+82" swimtime="00:01:23.39" resultid="102515" heatid="105328" lane="6" entrytime="00:01:19.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="259" reactiontime="+83" swimtime="00:05:44.92" resultid="102516" heatid="106063" lane="4" entrytime="00:05:29.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.70" />
                    <SPLIT distance="100" swimtime="00:01:17.49" />
                    <SPLIT distance="150" swimtime="00:02:01.62" />
                    <SPLIT distance="200" swimtime="00:02:46.28" />
                    <SPLIT distance="250" swimtime="00:03:31.59" />
                    <SPLIT distance="300" swimtime="00:04:16.93" />
                    <SPLIT distance="350" swimtime="00:05:01.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1942-03-23" firstname="Ryszard" gender="M" lastname="RYBARCZYK" nation="POL" swrid="4992649" athleteid="102517">
              <RESULTS>
                <RESULT eventid="98798" points="131" reactiontime="+105" swimtime="00:00:41.11" resultid="102518" heatid="105125" lane="0" entrytime="00:00:40.00" />
                <RESULT comment="K12" eventid="98956" reactiontime="+114" status="DSQ" swimtime="00:00:00.00" resultid="102519" heatid="105197" lane="0" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.68" />
                    <SPLIT distance="100" swimtime="00:01:56.53" />
                    <SPLIT distance="150" swimtime="00:03:02.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="155" reactiontime="+119" swimtime="00:01:48.78" resultid="102520" heatid="105250" lane="1" entrytime="00:01:47.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="102521" heatid="105295" lane="7" entrytime="00:04:31.52" />
                <RESULT eventid="99425" points="182" reactiontime="+105" swimtime="00:00:46.98" resultid="102522" heatid="105352" lane="7" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="WAR" clubid="100416" name="Victory Masters Elblag">
          <CONTACT city="Elbląg" name="Latecki" street="Łokietka 45" zip="82-300" />
          <ATHLETES>
            <ATHLETE birthdate="1980-03-21" firstname="Tomasz" gender="M" lastname="WYSOCKI" nation="POL" swrid="4919378" athleteid="100423">
              <RESULTS>
                <RESULT eventid="98798" points="490" reactiontime="+93" swimtime="00:00:26.51" resultid="100424" heatid="105141" lane="5" entrytime="00:00:26.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-11-18" firstname="Danuta" gender="F" lastname="GOJLIK" nation="POL" athleteid="100425">
              <RESULTS>
                <RESULT eventid="98940" points="175" reactiontime="+112" swimtime="00:04:08.53" resultid="100426" heatid="105191" lane="3" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.31" />
                    <SPLIT distance="100" swimtime="00:02:01.96" />
                    <SPLIT distance="150" swimtime="00:03:06.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="163" reactiontime="+83" swimtime="00:01:57.62" resultid="100427" heatid="105245" lane="8" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" status="DNS" swimtime="00:00:00.00" resultid="100428" heatid="105259" lane="0" entrytime="00:00:58.00" />
                <RESULT eventid="99409" points="156" reactiontime="+101" swimtime="00:00:54.76" resultid="100429" heatid="105346" lane="2" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-08-31" firstname="Karolina" gender="F" lastname="KARAŚ" nation="POL" swrid="4992650" athleteid="100430">
              <RESULTS>
                <RESULT eventid="98777" points="124" reactiontime="+101" swimtime="00:00:47.56" resultid="100431" heatid="105114" lane="1" entrytime="00:00:42.54" entrycourse="SCM" />
                <RESULT eventid="98863" points="143" swimtime="00:15:42.63" resultid="100432" heatid="105405" lane="4" entrytime="00:12:00.00" />
                <RESULT eventid="98972" points="125" reactiontime="+95" swimtime="00:01:44.07" resultid="100433" heatid="105206" lane="6" entrytime="00:01:33.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="132" reactiontime="+99" swimtime="00:03:41.52" resultid="100434" heatid="105290" lane="7" entrytime="00:03:21.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.13" />
                    <SPLIT distance="100" swimtime="00:01:51.77" />
                    <SPLIT distance="150" swimtime="00:02:47.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="146" reactiontime="+101" swimtime="00:07:34.01" resultid="100435" heatid="106056" lane="1" entrytime="00:06:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.27" />
                    <SPLIT distance="100" swimtime="00:01:53.03" />
                    <SPLIT distance="150" swimtime="00:02:51.42" />
                    <SPLIT distance="200" swimtime="00:03:49.50" />
                    <SPLIT distance="250" swimtime="00:04:47.86" />
                    <SPLIT distance="300" swimtime="00:05:45.87" />
                    <SPLIT distance="350" swimtime="00:06:41.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-05-05" firstname="Beata" gender="F" lastname="KARAŚ" nation="POL" swrid="4992651" athleteid="100436">
              <RESULTS>
                <RESULT eventid="98863" points="167" swimtime="00:14:56.38" resultid="100437" heatid="105405" lane="0" entrytime="00:13:30.00" />
                <RESULT eventid="99004" points="119" reactiontime="+100" swimtime="00:04:07.55" resultid="100438" heatid="105230" lane="9" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.88" />
                    <SPLIT distance="100" swimtime="00:01:58.54" />
                    <SPLIT distance="150" swimtime="00:03:02.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99266" points="141" reactiontime="+120" swimtime="00:08:35.39" resultid="100439" heatid="106045" lane="5" entrytime="00:08:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.59" />
                    <SPLIT distance="100" swimtime="00:01:57.15" />
                    <SPLIT distance="150" swimtime="00:03:06.99" />
                    <SPLIT distance="200" swimtime="00:04:13.83" />
                    <SPLIT distance="250" swimtime="00:05:28.57" />
                    <SPLIT distance="300" swimtime="00:06:43.81" />
                    <SPLIT distance="350" swimtime="00:07:40.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="115" reactiontime="+109" swimtime="00:01:54.90" resultid="100440" heatid="105321" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="167" reactiontime="+114" swimtime="00:07:13.84" resultid="100441" heatid="106057" lane="4" entrytime="00:07:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.73" />
                    <SPLIT distance="100" swimtime="00:01:45.46" />
                    <SPLIT distance="150" swimtime="00:02:40.92" />
                    <SPLIT distance="200" swimtime="00:03:36.73" />
                    <SPLIT distance="250" swimtime="00:04:31.92" />
                    <SPLIT distance="300" swimtime="00:05:27.83" />
                    <SPLIT distance="350" swimtime="00:06:22.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-02-04" firstname="Ewa" gender="F" lastname="KERNER MATEUSIAK" nation="POL" swrid="4992652" athleteid="100442">
              <RESULTS>
                <RESULT eventid="98777" points="93" reactiontime="+191" swimtime="00:00:52.22" resultid="100443" heatid="105113" lane="2" entrytime="00:00:49.73" entrycourse="SCM" />
                <RESULT eventid="98863" points="81" swimtime="00:18:59.19" resultid="100444" heatid="105406" lane="3" entrytime="00:16:00.00" />
                <RESULT eventid="98907" points="81" reactiontime="+103" swimtime="00:01:02.39" resultid="100445" heatid="105172" lane="3" entrytime="00:01:25.00" />
                <RESULT eventid="98940" status="DNS" swimtime="00:00:00.00" resultid="100446" heatid="105191" lane="8" entrytime="00:06:00.00" />
                <RESULT eventid="99089" points="59" reactiontime="+126" swimtime="00:02:44.42" resultid="100447" heatid="105243" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="61" reactiontime="+175" swimtime="00:02:27.33" resultid="100448" heatid="105277" lane="1" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="57" reactiontime="+168" swimtime="00:01:16.59" resultid="100449" heatid="105344" lane="1" entrytime="00:01:07.00" />
                <RESULT eventid="99457" points="76" reactiontime="+139" swimtime="00:09:23.17" resultid="100450" heatid="106057" lane="1" entrytime="00:09:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.74" />
                    <SPLIT distance="100" swimtime="00:02:09.41" />
                    <SPLIT distance="150" swimtime="00:03:21.77" />
                    <SPLIT distance="200" swimtime="00:04:35.30" />
                    <SPLIT distance="250" swimtime="00:05:48.02" />
                    <SPLIT distance="300" swimtime="00:07:00.66" />
                    <SPLIT distance="350" swimtime="00:08:13.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-06-06" firstname="Andrzej" gender="M" lastname="PASIECZNY" nation="POL" swrid="4605096" athleteid="100451">
              <RESULTS>
                <RESULT eventid="98798" points="377" reactiontime="+99" swimtime="00:00:28.94" resultid="100452" heatid="105135" lane="3" entrytime="00:00:29.35" />
                <RESULT eventid="99020" points="423" reactiontime="+89" swimtime="00:02:28.50" resultid="100453" heatid="105236" lane="7" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="100" swimtime="00:01:09.44" />
                    <SPLIT distance="150" swimtime="00:01:47.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="439" reactiontime="+95" swimtime="00:02:14.18" resultid="100454" heatid="105303" lane="1" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.82" />
                    <SPLIT distance="100" swimtime="00:01:06.17" />
                    <SPLIT distance="150" swimtime="00:01:40.52" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="04" eventid="99361" reactiontime="+72" status="DSQ" swimtime="00:00:00.00" resultid="100455" heatid="105330" lane="6" entrytime="00:01:05.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="437" reactiontime="+96" swimtime="00:04:49.86" resultid="100456" heatid="106060" lane="9" entrytime="00:04:50.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                    <SPLIT distance="100" swimtime="00:01:09.67" />
                    <SPLIT distance="150" swimtime="00:01:46.79" />
                    <SPLIT distance="200" swimtime="00:02:23.94" />
                    <SPLIT distance="250" swimtime="00:03:00.72" />
                    <SPLIT distance="300" swimtime="00:03:38.36" />
                    <SPLIT distance="350" swimtime="00:04:14.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-03-12" firstname="Grzegorz" gender="M" lastname="LATECKI" nation="POL" swrid="4754637" athleteid="100457">
              <RESULTS>
                <RESULT eventid="98798" points="389" reactiontime="+86" swimtime="00:00:28.64" resultid="100458" heatid="105137" lane="3" entrytime="00:00:28.50" />
                <RESULT eventid="98924" points="367" reactiontime="+83" swimtime="00:00:33.57" resultid="100459" heatid="105188" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="99170" points="395" reactiontime="+90" swimtime="00:00:30.55" resultid="100460" heatid="105274" lane="0" entrytime="00:00:29.90" />
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="100461" heatid="105340" lane="4" entrytime="00:02:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1938-02-09" firstname="Krystyna" gender="F" lastname="OPALIŃSKA" nation="POL" athleteid="100462">
              <RESULTS>
                <RESULT eventid="98777" points="27" reactiontime="+135" swimtime="00:01:18.94" resultid="100463" heatid="105113" lane="9" entrytime="00:01:15.00" />
                <RESULT eventid="98907" points="47" reactiontime="+126" swimtime="00:01:14.68" resultid="100464" heatid="105172" lane="4" entrytime="00:01:10.00" />
                <RESULT eventid="99314" status="DNS" swimtime="00:00:00.00" resultid="100465" heatid="105277" lane="7" entrytime="00:02:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-12-25" firstname="Waldemar" gender="M" lastname="MACIESZA" nation="POL" athleteid="100466">
              <RESULTS>
                <RESULT eventid="99091" points="180" reactiontime="+101" swimtime="00:01:43.41" resultid="100467" heatid="105251" lane="8" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="202" reactiontime="+114" swimtime="00:00:45.42" resultid="100468" heatid="105353" lane="6" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-01" firstname="Tomasz" gender="M" lastname="GLEB" nation="POL" athleteid="105077">
              <RESULTS>
                <RESULT eventid="98798" points="318" reactiontime="+82" swimtime="00:00:30.63" resultid="105078" heatid="105131" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="98891" points="289" swimtime="00:21:56.48" resultid="105079" heatid="105422" lane="4" entrytime="00:22:01.00" />
                <RESULT eventid="98956" points="298" reactiontime="+82" swimtime="00:03:10.12" resultid="105080" heatid="105200" lane="8" entrytime="00:03:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.12" />
                    <SPLIT distance="100" swimtime="00:01:31.28" />
                    <SPLIT distance="150" swimtime="00:02:21.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="350" reactiontime="+93" swimtime="00:01:06.53" resultid="105081" heatid="105221" lane="5" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="244" reactiontime="+106" swimtime="00:06:30.21" resultid="105082" heatid="106049" lane="4" entrytime="00:07:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.68" />
                    <SPLIT distance="100" swimtime="00:01:40.78" />
                    <SPLIT distance="150" swimtime="00:02:35.46" />
                    <SPLIT distance="200" swimtime="00:03:30.67" />
                    <SPLIT distance="250" swimtime="00:04:22.36" />
                    <SPLIT distance="300" swimtime="00:05:13.47" />
                    <SPLIT distance="350" swimtime="00:05:53.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="306" reactiontime="+98" swimtime="00:05:26.56" resultid="105083" heatid="106062" lane="7" entrytime="00:05:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                    <SPLIT distance="100" swimtime="00:01:15.78" />
                    <SPLIT distance="150" swimtime="00:01:57.55" />
                    <SPLIT distance="200" swimtime="00:02:39.95" />
                    <SPLIT distance="250" swimtime="00:03:23.16" />
                    <SPLIT distance="300" swimtime="00:04:06.30" />
                    <SPLIT distance="350" swimtime="00:04:47.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="104986" name="WOPR Kutno">
          <ATHLETES>
            <ATHLETE birthdate="1932-03-11" firstname="Kazimierz" gender="M" lastname="FROM" nation="POL" athleteid="104987">
              <RESULTS>
                <RESULT eventid="98798" points="40" reactiontime="+134" swimtime="00:01:01.03" resultid="104988" heatid="105123" lane="4" entrytime="00:00:58.00" />
                <RESULT eventid="98924" points="30" reactiontime="+100" swimtime="00:01:17.00" resultid="104989" heatid="105180" lane="6" entrytime="00:01:16.00" />
                <RESULT eventid="99186" points="25" reactiontime="+109" swimtime="00:02:56.73" resultid="104990" heatid="105281" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="26" reactiontime="+102" swimtime="00:06:14.02" resultid="104991" heatid="105336" lane="9" entrytime="00:05:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.07" />
                    <SPLIT distance="100" swimtime="00:03:05.22" />
                    <SPLIT distance="150" swimtime="00:04:40.53" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters, Rekord Polski Masters" eventid="98891" points="25" swimtime="00:49:31.63" resultid="104992" heatid="105425" lane="7" entrytime="00:50:00.00" />
                <RESULT eventid="98988" points="33" reactiontime="+126" swimtime="00:02:25.24" resultid="104993" heatid="105213" lane="7" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="29" reactiontime="+132" swimtime="00:05:31.74" resultid="104994" heatid="105295" lane="8" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.25" />
                    <SPLIT distance="100" swimtime="00:02:36.47" />
                    <SPLIT distance="150" swimtime="00:04:10.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="27" reactiontime="+136" swimtime="00:12:10.35" resultid="104995" heatid="106067" lane="5" entrytime="00:12:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.15" />
                    <SPLIT distance="100" swimtime="00:02:47.36" />
                    <SPLIT distance="150" swimtime="00:04:21.71" />
                    <SPLIT distance="200" swimtime="00:05:58.47" />
                    <SPLIT distance="250" swimtime="00:07:32.01" />
                    <SPLIT distance="300" swimtime="00:09:06.35" />
                    <SPLIT distance="350" swimtime="00:10:39.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="101163" name="WOPR Tczew">
          <CONTACT name="Hebel Aleksanrda" />
          <ATHLETES>
            <ATHLETE birthdate="1987-06-22" firstname="Aleksandra" gender="F" lastname="HEBEL" nation="POL" swrid="4754694" athleteid="101164">
              <RESULTS>
                <RESULT eventid="98777" points="344" reactiontime="+115" swimtime="00:00:33.85" resultid="101165" heatid="105117" lane="0" entrytime="00:00:35.08" entrycourse="SCM" />
                <RESULT eventid="98907" points="232" reactiontime="+98" swimtime="00:00:44.00" resultid="101166" heatid="105175" lane="8" entrytime="00:00:42.00" />
                <RESULT eventid="98972" points="291" reactiontime="+115" swimtime="00:01:18.49" resultid="101167" heatid="105209" lane="0" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="234" reactiontime="+111" swimtime="00:01:34.31" resultid="101168" heatid="105278" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="257" reactiontime="+113" swimtime="00:02:57.52" resultid="101169" heatid="105291" lane="3" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                    <SPLIT distance="100" swimtime="00:01:24.75" />
                    <SPLIT distance="150" swimtime="00:02:12.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="232" reactiontime="+132" swimtime="00:03:21.76" resultid="101170" heatid="105333" lane="5" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.16" />
                    <SPLIT distance="100" swimtime="00:01:37.75" />
                    <SPLIT distance="150" swimtime="00:02:30.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-10-28" firstname="Andrzej" gender="M" lastname="GOŁEMBIEWSKI" nation="POL" athleteid="101171">
              <RESULTS>
                <RESULT eventid="98956" points="400" reactiontime="+88" swimtime="00:02:52.36" resultid="101172" heatid="105203" lane="1" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.49" />
                    <SPLIT distance="100" swimtime="00:01:22.82" />
                    <SPLIT distance="150" swimtime="00:02:08.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="449" reactiontime="+85" swimtime="00:01:16.30" resultid="101173" heatid="105256" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="345" reactiontime="+89" swimtime="00:02:25.43" resultid="101174" heatid="105301" lane="8" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.47" />
                    <SPLIT distance="100" swimtime="00:01:07.43" />
                    <SPLIT distance="150" swimtime="00:01:46.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="468" reactiontime="+97" swimtime="00:00:34.33" resultid="101175" heatid="105360" lane="4" entrytime="00:00:34.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WMT" nation="POL" region="MAZ" clubid="101571" name="Warsaw Masters Team">
          <CONTACT city="Warszawa" email="wojciech.kaluzynski@gmail.com" name="KAŁUŻYŃSKI Wojciech" phone="607 45 4444" />
          <ATHLETES>
            <ATHLETE birthdate="1935-06-16" firstname="Elżbieta" gender="F" lastname="JANIK" nation="POL" swrid="4270351" athleteid="101572">
              <RESULTS>
                <RESULT eventid="98907" points="45" reactiontime="+95" swimtime="00:01:15.58" resultid="101573" heatid="105172" lane="5" entrytime="00:01:10.00" />
                <RESULT eventid="99314" points="48" reactiontime="+101" swimtime="00:02:39.24" resultid="101574" heatid="105277" lane="2" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="47" reactiontime="+102" swimtime="00:05:43.12" resultid="101575" heatid="105332" lane="1" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.34" />
                    <SPLIT distance="100" swimtime="00:02:48.76" />
                    <SPLIT distance="150" swimtime="00:04:16.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Mirosław" gender="M" lastname="WARCHOŁ" nation="POL" swrid="4222718" athleteid="101576">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski Masters" eventid="98830" points="341" reactiontime="+95" swimtime="00:02:43.04" resultid="101577" heatid="105153" lane="0" entrytime="00:02:57.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.03" />
                    <SPLIT distance="100" swimtime="00:01:16.26" />
                    <SPLIT distance="150" swimtime="00:02:06.80" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="98988" points="400" reactiontime="+85" swimtime="00:01:03.62" resultid="101578" heatid="105220" lane="7" entrytime="00:01:08.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="328" reactiontime="+81" swimtime="00:01:15.30" resultid="101579" heatid="105284" lane="5" entrytime="00:01:18.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.08" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99393" points="324" reactiontime="+89" swimtime="00:02:42.84" resultid="101580" heatid="105340" lane="1" entrytime="00:02:54.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.95" />
                    <SPLIT distance="100" swimtime="00:01:18.49" />
                    <SPLIT distance="150" swimtime="00:02:00.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-10-03" firstname="Ryszard" gender="M" lastname="SIELSKI" nation="POL" swrid="4129765" athleteid="101581">
              <RESULTS>
                <RESULT eventid="98830" points="57" reactiontime="+124" swimtime="00:04:55.79" resultid="101582" heatid="105148" lane="3" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.58" />
                    <SPLIT distance="100" swimtime="00:02:33.39" />
                    <SPLIT distance="150" swimtime="00:03:49.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98891" points="52" swimtime="00:38:48.00" resultid="101583" heatid="105425" lane="2" entrytime="00:40:00.00" />
                <RESULT eventid="98924" points="30" reactiontime="+88" swimtime="00:01:16.99" resultid="101584" heatid="105180" lane="3" entrytime="00:00:59.00" />
                <RESULT eventid="98956" points="58" reactiontime="+120" swimtime="00:05:26.79" resultid="101585" heatid="105196" lane="6" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.15" />
                    <SPLIT distance="100" swimtime="00:02:38.21" />
                    <SPLIT distance="150" swimtime="00:04:03.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="101586" heatid="105249" lane="7" entrytime="00:02:20.00" />
                <RESULT eventid="99282" status="DNS" swimtime="00:00:00.00" resultid="101587" heatid="106049" lane="9" entrytime="00:08:00.00" />
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="101588" heatid="105325" lane="9" entrytime="00:02:40.00" />
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="101589" heatid="105336" lane="8" entrytime="00:05:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-21" firstname="Marianna" gender="F" lastname="GAJDUS" nation="POL" swrid="4992655" athleteid="101590">
              <RESULTS>
                <RESULT eventid="98814" points="293" swimtime="00:03:09.90" resultid="101591" heatid="105146" lane="7" entrytime="00:03:03.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.04" />
                    <SPLIT distance="100" swimtime="00:01:30.76" />
                    <SPLIT distance="150" swimtime="00:02:26.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="325" reactiontime="+77" swimtime="00:01:15.66" resultid="101592" heatid="105209" lane="1" entrytime="00:01:15.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="361" reactiontime="+73" swimtime="00:00:35.20" resultid="101593" heatid="105262" lane="6" entrytime="00:00:35.83" />
                <RESULT eventid="99202" points="317" reactiontime="+71" swimtime="00:02:45.56" resultid="101594" heatid="105292" lane="6" entrytime="00:02:45.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                    <SPLIT distance="100" swimtime="00:01:21.24" />
                    <SPLIT distance="150" swimtime="00:02:05.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="307" reactiontime="+64" swimtime="00:01:22.97" resultid="101595" heatid="105323" lane="9" entrytime="00:01:21.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="301" reactiontime="+76" swimtime="00:05:56.53" resultid="101596" heatid="106055" lane="0" entrytime="00:05:55.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.14" />
                    <SPLIT distance="100" swimtime="00:01:24.46" />
                    <SPLIT distance="150" swimtime="00:02:10.41" />
                    <SPLIT distance="200" swimtime="00:02:56.42" />
                    <SPLIT distance="250" swimtime="00:03:42.34" />
                    <SPLIT distance="300" swimtime="00:04:28.18" />
                    <SPLIT distance="350" swimtime="00:05:14.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-05" firstname="Bartłomiej" gender="M" lastname="PAWŁOWSKI" nation="POL" swrid="4992755" athleteid="101597">
              <RESULTS>
                <RESULT eventid="98798" points="359" reactiontime="+89" swimtime="00:00:29.41" resultid="101598" heatid="105137" lane="1" entrytime="00:00:28.50" />
                <RESULT eventid="98988" points="365" reactiontime="+82" swimtime="00:01:05.62" resultid="101599" heatid="105213" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="334" reactiontime="+82" swimtime="00:01:24.22" resultid="101600" heatid="105256" lane="9" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="101601" heatid="105295" lane="0" />
                <RESULT eventid="99425" points="418" reactiontime="+83" swimtime="00:00:35.65" resultid="101602" heatid="105360" lane="5" entrytime="00:00:34.78" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-05-14" firstname="Sebastian" gender="M" lastname="WOJCIECHOWSKI" nation="POL" athleteid="101603">
              <RESULTS>
                <RESULT eventid="98891" points="180" swimtime="00:25:42.42" resultid="101604" heatid="105422" lane="2" entrytime="00:22:30.00" />
                <RESULT eventid="99218" points="184" reactiontime="+90" swimtime="00:02:59.21" resultid="101605" heatid="105297" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.37" />
                    <SPLIT distance="100" swimtime="00:01:23.90" />
                    <SPLIT distance="150" swimtime="00:02:13.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="187" reactiontime="+97" swimtime="00:06:24.35" resultid="101606" heatid="106065" lane="2" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.09" />
                    <SPLIT distance="100" swimtime="00:01:24.83" />
                    <SPLIT distance="150" swimtime="00:02:13.53" />
                    <SPLIT distance="200" swimtime="00:03:03.51" />
                    <SPLIT distance="250" swimtime="00:03:54.13" />
                    <SPLIT distance="300" swimtime="00:04:45.52" />
                    <SPLIT distance="350" swimtime="00:05:35.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-06-17" firstname="Leszek" gender="M" lastname="MADEJ" nation="POL" swrid="4183799" athleteid="101607">
              <RESULTS>
                <RESULT eventid="98798" points="442" reactiontime="+78" swimtime="00:00:27.45" resultid="101608" heatid="105139" lane="5" entrytime="00:00:27.43" />
                <RESULT eventid="98956" points="374" reactiontime="+87" swimtime="00:02:56.25" resultid="101609" heatid="105203" lane="2" entrytime="00:02:57.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.54" />
                    <SPLIT distance="100" swimtime="00:01:25.49" />
                    <SPLIT distance="150" swimtime="00:02:11.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="486" reactiontime="+77" swimtime="00:00:59.64" resultid="101610" heatid="105226" lane="7" entrytime="00:00:59.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.46" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99091" points="405" reactiontime="+82" swimtime="00:01:18.97" resultid="101611" heatid="105255" lane="4" entrytime="00:01:21.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="443" reactiontime="+76" swimtime="00:02:13.71" resultid="101612" heatid="105304" lane="8" entrytime="00:02:12.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                    <SPLIT distance="100" swimtime="00:01:07.30" />
                    <SPLIT distance="150" swimtime="00:01:41.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="429" reactiontime="+74" swimtime="00:00:35.36" resultid="101613" heatid="105359" lane="9" entrytime="00:00:36.56" />
                <RESULT comment="Rekord Polski Masters" eventid="99473" points="439" reactiontime="+78" swimtime="00:04:49.39" resultid="101614" heatid="106061" lane="6" entrytime="00:04:57.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                    <SPLIT distance="100" swimtime="00:01:10.68" />
                    <SPLIT distance="150" swimtime="00:01:48.14" />
                    <SPLIT distance="200" swimtime="00:02:26.17" />
                    <SPLIT distance="250" swimtime="00:03:02.86" />
                    <SPLIT distance="300" swimtime="00:03:39.03" />
                    <SPLIT distance="350" swimtime="00:04:14.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-05-11" firstname="Sara" gender="F" lastname="DEBEVEC" nation="POL" athleteid="101615">
              <RESULTS>
                <RESULT eventid="98777" status="DNS" swimtime="00:00:00.00" resultid="101616" heatid="105115" lane="7" entrytime="00:00:39.00" />
                <RESULT eventid="98863" status="WDR" swimtime="00:00:00.00" resultid="101617" entrytime="00:13:50.00" />
                <RESULT eventid="99154" points="167" reactiontime="+94" swimtime="00:00:45.48" resultid="101618" heatid="105261" lane="9" entrytime="00:00:40.00" />
                <RESULT comment="04" eventid="99202" reactiontime="+87" status="DSQ" swimtime="00:00:00.00" resultid="101619" heatid="105290" lane="6" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.63" />
                    <SPLIT distance="100" swimtime="00:01:30.90" />
                    <SPLIT distance="150" swimtime="00:02:22.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="160" reactiontime="+148" swimtime="00:01:43.01" resultid="101620" heatid="105322" lane="0" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="202" reactiontime="+122" swimtime="00:06:47.00" resultid="101621" heatid="106057" lane="6" entrytime="00:07:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.56" />
                    <SPLIT distance="100" swimtime="00:01:35.30" />
                    <SPLIT distance="150" swimtime="00:02:27.18" />
                    <SPLIT distance="200" swimtime="00:03:20.04" />
                    <SPLIT distance="250" swimtime="00:04:12.92" />
                    <SPLIT distance="300" swimtime="00:05:05.94" />
                    <SPLIT distance="350" swimtime="00:05:57.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-05-20" firstname="Anna" gender="F" lastname="STANISŁAWSKA" nation="POL" swrid="4992660" athleteid="101622">
              <RESULTS>
                <RESULT eventid="98777" points="282" reactiontime="+105" swimtime="00:00:36.17" resultid="101623" heatid="105116" lane="7" entrytime="00:00:36.40" entrycourse="SCM" />
                <RESULT eventid="98972" points="254" reactiontime="+113" swimtime="00:01:22.21" resultid="101624" heatid="105205" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99004" points="180" reactiontime="+109" swimtime="00:03:35.42" resultid="101625" heatid="105230" lane="8" entrytime="00:03:53.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.42" />
                    <SPLIT distance="100" swimtime="00:01:41.35" />
                    <SPLIT distance="150" swimtime="00:02:39.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="208" reactiontime="+106" swimtime="00:00:42.30" resultid="101626" heatid="105260" lane="1" entrytime="00:00:43.03" />
                <RESULT eventid="99202" points="215" reactiontime="+104" swimtime="00:03:08.54" resultid="101627" heatid="105291" lane="9" entrytime="00:03:12.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.51" />
                    <SPLIT distance="100" swimtime="00:01:31.17" />
                    <SPLIT distance="150" swimtime="00:02:21.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99344" points="169" reactiontime="+114" swimtime="00:01:41.24" resultid="101628" heatid="105321" lane="5" entrytime="00:01:52.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="206" reactiontime="+117" swimtime="00:06:44.69" resultid="101629" heatid="106056" lane="0" entrytime="00:06:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.53" />
                    <SPLIT distance="100" swimtime="00:01:36.07" />
                    <SPLIT distance="150" swimtime="00:02:28.72" />
                    <SPLIT distance="200" swimtime="00:03:21.68" />
                    <SPLIT distance="250" swimtime="00:04:12.17" />
                    <SPLIT distance="300" swimtime="00:05:03.65" />
                    <SPLIT distance="350" swimtime="00:05:54.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-05-15" firstname="Jerzy" gender="M" lastname="LESZCZYŃSKI" nation="POL" athleteid="101630">
              <RESULTS>
                <RESULT eventid="98798" points="335" reactiontime="+69" swimtime="00:00:30.09" resultid="101631" heatid="105135" lane="8" entrytime="00:00:29.60" />
                <RESULT eventid="98830" points="276" reactiontime="+84" swimtime="00:02:54.93" resultid="101632" heatid="105153" lane="2" entrytime="00:02:55.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                    <SPLIT distance="100" swimtime="00:01:23.98" />
                    <SPLIT distance="150" swimtime="00:02:14.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="296" reactiontime="+81" swimtime="00:03:10.53" resultid="101633" heatid="105201" lane="4" entrytime="00:03:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.57" />
                    <SPLIT distance="100" swimtime="00:01:29.46" />
                    <SPLIT distance="150" swimtime="00:02:19.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="333" reactiontime="+76" swimtime="00:01:07.67" resultid="101634" heatid="105220" lane="6" entrytime="00:01:08.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="321" reactiontime="+73" swimtime="00:01:25.35" resultid="101635" heatid="105254" lane="6" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="101636" heatid="105299" lane="5" entrytime="00:02:35.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-11-07" firstname="Andrzej" gender="M" lastname="LEWANDOWSKI" nation="POL" swrid="4992668" athleteid="101637">
              <RESULTS>
                <RESULT eventid="98798" points="260" reactiontime="+78" swimtime="00:00:32.73" resultid="101638" heatid="105131" lane="8" entrytime="00:00:31.54" />
                <RESULT eventid="98956" points="253" reactiontime="+88" swimtime="00:03:20.74" resultid="101639" heatid="105201" lane="3" entrytime="00:03:09.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.38" />
                    <SPLIT distance="100" swimtime="00:01:33.24" />
                    <SPLIT distance="150" swimtime="00:02:26.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="220" reactiontime="+93" swimtime="00:01:17.61" resultid="101640" heatid="105218" lane="2" entrytime="00:01:10.95" />
                <RESULT eventid="99091" points="285" reactiontime="+85" swimtime="00:01:28.83" resultid="101641" heatid="105254" lane="7" entrytime="00:01:24.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="213" reactiontime="+91" swimtime="00:00:37.52" resultid="101642" heatid="105269" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="99425" points="354" reactiontime="+91" swimtime="00:00:37.67" resultid="101643" heatid="105359" lane="5" entrytime="00:00:35.95" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-08-02" firstname="Tomasz" gender="M" lastname="JĄKALSKI" nation="POL" swrid="4992693" athleteid="101644">
              <RESULTS>
                <RESULT eventid="98924" points="465" reactiontime="+63" swimtime="00:00:31.03" resultid="101645" heatid="105190" lane="7" entrytime="00:00:29.70" />
                <RESULT eventid="99186" points="412" reactiontime="+76" swimtime="00:01:09.79" resultid="101646" heatid="105287" lane="5" entrytime="00:01:08.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="218" reactiontime="+74" swimtime="00:03:05.73" resultid="101647" heatid="105342" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.58" />
                    <SPLIT distance="100" swimtime="00:01:30.08" />
                    <SPLIT distance="150" swimtime="00:02:15.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="303" reactiontime="+99" swimtime="00:06:02.77" resultid="103025" heatid="106051" lane="5" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.75" />
                    <SPLIT distance="100" swimtime="00:01:14.42" />
                    <SPLIT distance="150" swimtime="00:02:01.30" />
                    <SPLIT distance="200" swimtime="00:02:48.67" />
                    <SPLIT distance="250" swimtime="00:03:39.27" />
                    <SPLIT distance="300" swimtime="00:04:30.70" />
                    <SPLIT distance="350" swimtime="00:05:16.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-05-14" firstname="Wojciech" gender="M" lastname="KAŁUŻYŃSKI" nation="POL" swrid="4992656" athleteid="101648">
              <RESULTS>
                <RESULT eventid="98798" points="321" reactiontime="+83" swimtime="00:00:30.53" resultid="101649" heatid="105132" lane="7" entrytime="00:00:30.99" />
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="101650" heatid="105148" lane="7" />
                <RESULT eventid="98924" points="252" reactiontime="+89" swimtime="00:00:38.02" resultid="101651" heatid="105185" lane="5" entrytime="00:00:38.00" />
                <RESULT eventid="98988" points="332" reactiontime="+90" swimtime="00:01:07.68" resultid="101652" heatid="105220" lane="3" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="246" reactiontime="+83" swimtime="00:00:35.77" resultid="101653" heatid="105268" lane="8" entrytime="00:00:37.00" />
                <RESULT eventid="99218" points="292" reactiontime="+92" swimtime="00:02:33.58" resultid="101654" heatid="105299" lane="3" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                    <SPLIT distance="100" swimtime="00:01:12.41" />
                    <SPLIT distance="150" swimtime="00:01:52.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="276" reactiontime="+92" swimtime="00:05:37.95" resultid="101655" heatid="106063" lane="3" entrytime="00:05:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                    <SPLIT distance="100" swimtime="00:01:18.83" />
                    <SPLIT distance="150" swimtime="00:02:01.56" />
                    <SPLIT distance="200" swimtime="00:02:45.71" />
                    <SPLIT distance="250" swimtime="00:03:29.27" />
                    <SPLIT distance="300" swimtime="00:04:13.62" />
                    <SPLIT distance="350" swimtime="00:04:56.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-10-02" firstname="Andrzej" gender="M" lastname="WISZNIEWSKI" nation="POL" swrid="4967430" athleteid="101656">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="101657" heatid="105125" lane="9" entrytime="00:00:40.00" />
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="101658" heatid="105150" lane="0" entrytime="00:03:50.20" />
                <RESULT eventid="98956" status="DNS" swimtime="00:00:00.00" resultid="101659" heatid="105197" lane="3" entrytime="00:03:54.20" />
                <RESULT eventid="99020" status="DNS" swimtime="00:00:00.00" resultid="101660" heatid="105233" lane="0" entrytime="00:03:59.60" />
                <RESULT eventid="99186" status="DNS" swimtime="00:00:00.00" resultid="101661" heatid="105282" lane="8" entrytime="00:01:54.30" />
                <RESULT eventid="99282" status="DNS" swimtime="00:00:00.00" resultid="101662" heatid="106048" lane="6" entrytime="00:08:30.20" />
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="101663" heatid="105325" lane="4" entrytime="00:01:55.40" />
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="101664" heatid="105337" lane="6" entrytime="00:03:45.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-03" firstname="Robert" gender="M" lastname="SUTOWSKI" nation="POL" swrid="4992657" athleteid="101665">
              <RESULTS>
                <RESULT eventid="98798" points="140" reactiontime="+124" swimtime="00:00:40.20" resultid="101666" heatid="105125" lane="3" entrytime="00:00:38.79" />
                <RESULT eventid="98830" points="112" reactiontime="+118" swimtime="00:03:55.85" resultid="101667" heatid="105148" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.07" />
                    <SPLIT distance="100" swimtime="00:01:59.50" />
                    <SPLIT distance="150" swimtime="00:03:10.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="89" reactiontime="+96" swimtime="00:00:53.82" resultid="101668" heatid="105181" lane="5" entrytime="00:00:53.46" />
                <RESULT eventid="98988" points="155" reactiontime="+124" swimtime="00:01:27.16" resultid="101669" heatid="105214" lane="4" entrytime="00:01:27.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="107" reactiontime="+118" swimtime="00:00:47.20" resultid="101670" heatid="105266" lane="0" entrytime="00:00:47.45" />
                <RESULT eventid="99218" points="146" reactiontime="+109" swimtime="00:03:13.52" resultid="101671" heatid="105297" lane="9" entrytime="00:03:09.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.87" />
                    <SPLIT distance="100" swimtime="00:01:33.62" />
                    <SPLIT distance="150" swimtime="00:02:25.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="167" reactiontime="+120" swimtime="00:06:39.46" resultid="101672" heatid="106067" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.14" />
                    <SPLIT distance="100" swimtime="00:01:33.73" />
                    <SPLIT distance="150" swimtime="00:02:24.82" />
                    <SPLIT distance="200" swimtime="00:03:16.69" />
                    <SPLIT distance="250" swimtime="00:04:08.97" />
                    <SPLIT distance="300" swimtime="00:05:01.00" />
                    <SPLIT distance="350" swimtime="00:05:51.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-18" firstname="Łukasz" gender="M" lastname="KUBISZEWSKI-JAKUBIAK" nation="POL" athleteid="101673">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="101674" heatid="105127" lane="5" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-03-04" firstname="Stefan" gender="M" lastname="BORODZIUK" nation="POL" athleteid="101675">
              <RESULTS>
                <RESULT eventid="98798" points="180" reactiontime="+97" swimtime="00:00:37.02" resultid="101676" heatid="105125" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="98891" points="91" swimtime="00:32:11.00" resultid="101677" heatid="105425" lane="5" entrytime="00:30:15.00" />
                <RESULT eventid="98924" points="110" reactiontime="+78" swimtime="00:00:50.13" resultid="101678" heatid="105182" lane="7" entrytime="00:00:49.00" />
                <RESULT eventid="98988" points="167" reactiontime="+92" swimtime="00:01:25.09" resultid="101679" heatid="105214" lane="5" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="98" reactiontime="+73" swimtime="00:01:52.41" resultid="101680" heatid="105282" lane="7" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="124" reactiontime="+98" swimtime="00:03:24.19" resultid="101681" heatid="105296" lane="7" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.46" />
                    <SPLIT distance="100" swimtime="00:01:38.84" />
                    <SPLIT distance="150" swimtime="00:02:33.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="101682" heatid="105336" lane="3" entrytime="00:04:20.00" />
                <RESULT eventid="99473" points="114" reactiontime="+108" swimtime="00:07:33.40" resultid="101683" heatid="106066" lane="3" entrytime="00:07:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.41" />
                    <SPLIT distance="100" swimtime="00:01:38.78" />
                    <SPLIT distance="150" swimtime="00:02:35.46" />
                    <SPLIT distance="200" swimtime="00:03:34.02" />
                    <SPLIT distance="250" swimtime="00:04:32.98" />
                    <SPLIT distance="300" swimtime="00:05:33.63" />
                    <SPLIT distance="350" swimtime="00:06:35.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-08-28" firstname="Katarzyna" gender="F" lastname="DOBCZYŃSKA" nation="POL" swrid="4754752" athleteid="101684">
              <RESULTS>
                <RESULT eventid="98777" points="238" reactiontime="+111" swimtime="00:00:38.29" resultid="101685" heatid="105115" lane="5" entrytime="00:00:37.89" entrycourse="SCM" />
                <RESULT eventid="98907" points="215" reactiontime="+100" swimtime="00:00:45.12" resultid="101686" heatid="105174" lane="7" entrytime="00:00:45.00" />
                <RESULT eventid="98972" points="240" reactiontime="+110" swimtime="00:01:23.74" resultid="101687" heatid="105207" lane="1" entrytime="00:01:23.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="229" reactiontime="+102" swimtime="00:01:34.96" resultid="101688" heatid="105278" lane="6" entrytime="00:01:33.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="219" reactiontime="+108" swimtime="00:03:07.33" resultid="101689" heatid="105291" lane="8" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.92" />
                    <SPLIT distance="100" swimtime="00:01:30.43" />
                    <SPLIT distance="150" swimtime="00:02:20.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="238" reactiontime="+103" swimtime="00:03:20.12" resultid="101690" heatid="105333" lane="9" entrytime="00:03:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.38" />
                    <SPLIT distance="100" swimtime="00:01:39.23" />
                    <SPLIT distance="150" swimtime="00:02:31.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-01" firstname="Paweł" gender="M" lastname="KOWALEWSKI" nation="POL" athleteid="101691">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski Masters" eventid="98891" points="410" swimtime="00:19:32.04" resultid="101692" heatid="105420" lane="1" entrytime="00:19:30.00" />
                <RESULT eventid="99218" points="386" reactiontime="+90" swimtime="00:02:20.07" resultid="101693" heatid="105303" lane="0" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                    <SPLIT distance="100" swimtime="00:01:07.54" />
                    <SPLIT distance="150" swimtime="00:01:43.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="424" reactiontime="+84" swimtime="00:04:52.84" resultid="101694" heatid="106060" lane="8" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                    <SPLIT distance="100" swimtime="00:01:11.07" />
                    <SPLIT distance="150" swimtime="00:01:48.62" />
                    <SPLIT distance="200" swimtime="00:02:26.97" />
                    <SPLIT distance="250" swimtime="00:03:04.28" />
                    <SPLIT distance="300" swimtime="00:03:41.18" />
                    <SPLIT distance="350" swimtime="00:04:17.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-05" firstname="Rafał" gender="M" lastname="SKOŚKIEWICZ" nation="POL" swrid="4183802" athleteid="101695">
              <RESULTS>
                <RESULT eventid="98798" points="387" reactiontime="+95" swimtime="00:00:28.69" resultid="101696" heatid="105136" lane="2" entrytime="00:00:29.00" />
                <RESULT eventid="98830" points="380" reactiontime="+86" swimtime="00:02:37.26" resultid="101697" heatid="105155" lane="6" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                    <SPLIT distance="100" swimtime="00:01:13.08" />
                    <SPLIT distance="150" swimtime="00:02:01.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="400" reactiontime="+89" swimtime="00:00:32.61" resultid="101698" heatid="105188" lane="8" entrytime="00:00:33.00" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="101699" heatid="105225" lane="9" entrytime="00:01:01.01" />
                <RESULT eventid="99186" points="386" reactiontime="+97" swimtime="00:01:11.28" resultid="101700" heatid="105287" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="307" reactiontime="+93" swimtime="00:02:45.82" resultid="101701" heatid="105341" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.43" />
                    <SPLIT distance="100" swimtime="00:01:22.40" />
                    <SPLIT distance="150" swimtime="00:02:05.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-28" firstname="Monika" gender="F" lastname="FIGURA" nation="POL" athleteid="101702">
              <RESULTS>
                <RESULT eventid="98907" points="312" reactiontime="+81" swimtime="00:00:39.89" resultid="101703" heatid="105176" lane="5" entrytime="00:00:39.00" />
                <RESULT eventid="98972" points="303" reactiontime="+75" swimtime="00:01:17.45" resultid="101704" heatid="105209" lane="9" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" status="DNS" swimtime="00:00:00.00" resultid="101705" heatid="105279" lane="5" entrytime="00:01:25.00" />
                <RESULT eventid="99377" points="260" reactiontime="+85" swimtime="00:03:14.30" resultid="101706" heatid="105333" lane="3" entrytime="00:03:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.63" />
                    <SPLIT distance="100" swimtime="00:01:33.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-02-23" firstname="Joanna" gender="F" lastname="GOŁĘBIOWSKA" nation="POL" swrid="4060381" athleteid="101707">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="98972" points="586" reactiontime="+81" swimtime="00:01:02.21" resultid="101708" heatid="105212" lane="3" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="515" reactiontime="+80" swimtime="00:00:31.27" resultid="101709" heatid="105264" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="99344" points="565" reactiontime="+78" swimtime="00:01:07.69" resultid="101710" heatid="105323" lane="4" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-04-28" firstname="Paweł" gender="M" lastname="ROGOSZ" nation="POL" swrid="4270348" athleteid="101711">
              <RESULTS>
                <RESULT eventid="98798" points="326" reactiontime="+100" swimtime="00:00:30.38" resultid="101712" heatid="105131" lane="7" entrytime="00:00:31.50" />
                <RESULT eventid="98830" points="353" reactiontime="+98" swimtime="00:02:41.21" resultid="101713" heatid="105154" lane="7" entrytime="00:02:51.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                    <SPLIT distance="100" swimtime="00:01:19.64" />
                    <SPLIT distance="150" swimtime="00:02:04.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="285" reactiontime="+104" swimtime="00:02:49.29" resultid="101714" heatid="105235" lane="9" entrytime="00:02:55.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.17" />
                    <SPLIT distance="100" swimtime="00:01:20.42" />
                    <SPLIT distance="150" swimtime="00:02:04.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="338" reactiontime="+112" swimtime="00:05:49.74" resultid="101715" heatid="106052" lane="0" entrytime="00:05:59.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.92" />
                    <SPLIT distance="100" swimtime="00:01:18.70" />
                    <SPLIT distance="150" swimtime="00:02:08.62" />
                    <SPLIT distance="200" swimtime="00:02:58.98" />
                    <SPLIT distance="250" swimtime="00:03:44.42" />
                    <SPLIT distance="300" swimtime="00:04:31.85" />
                    <SPLIT distance="350" swimtime="00:05:11.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="309" reactiontime="+108" swimtime="00:01:13.67" resultid="101716" heatid="105328" lane="3" entrytime="00:01:19.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="257" reactiontime="+92" swimtime="00:02:55.99" resultid="101717" heatid="105339" lane="5" entrytime="00:02:58.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.25" />
                    <SPLIT distance="100" swimtime="00:01:25.68" />
                    <SPLIT distance="150" swimtime="00:02:11.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-06-07" firstname="Olga" gender="F" lastname="KRYSIAK" nation="POL" swrid="4072533" athleteid="101718">
              <RESULTS>
                <RESULT eventid="98777" status="DNS" swimtime="00:00:00.00" resultid="101719" heatid="105121" lane="9" entrytime="00:00:29.20" entrycourse="LCM" />
                <RESULT eventid="98972" status="DNS" swimtime="00:00:00.00" resultid="101720" heatid="105212" lane="8" entrytime="00:01:03.90" />
                <RESULT eventid="99154" status="DNS" swimtime="00:00:00.00" resultid="101721" heatid="105263" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="99202" status="DNS" swimtime="00:00:00.00" resultid="101722" heatid="105294" lane="9" entrytime="00:02:26.50" />
                <RESULT eventid="99457" status="WDR" swimtime="00:00:00.00" resultid="101723" entrytime="00:05:20.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-12-11" firstname="Igor" gender="M" lastname="RĘBAS" nation="POL" swrid="4251117" athleteid="101724">
              <RESULTS>
                <RESULT eventid="98798" points="483" reactiontime="+82" swimtime="00:00:26.64" resultid="101725" heatid="105142" lane="0" entrytime="00:00:26.20" />
                <RESULT eventid="98988" points="523" reactiontime="+79" swimtime="00:00:58.21" resultid="101726" heatid="105227" lane="2" entrytime="00:00:57.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="522" reactiontime="+83" swimtime="00:00:27.85" resultid="101727" heatid="105275" lane="3" entrytime="00:00:27.50" />
                <RESULT eventid="99361" points="495" reactiontime="+69" swimtime="00:01:02.94" resultid="101728" heatid="105331" lane="7" entrytime="00:01:01.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98830" points="437" reactiontime="+86" swimtime="00:02:30.22" resultid="103022" heatid="105156" lane="2" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.34" />
                    <SPLIT distance="100" swimtime="00:01:10.10" />
                    <SPLIT distance="150" swimtime="00:01:55.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" status="DNS" swimtime="00:00:00.00" resultid="103023" heatid="105236" lane="2" entrytime="00:02:30.00" />
                <RESULT eventid="99282" points="369" reactiontime="+87" swimtime="00:05:39.88" resultid="104384" heatid="106051" lane="3" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.46" />
                    <SPLIT distance="100" swimtime="00:01:07.45" />
                    <SPLIT distance="150" swimtime="00:01:53.65" />
                    <SPLIT distance="200" swimtime="00:02:39.15" />
                    <SPLIT distance="250" swimtime="00:03:29.80" />
                    <SPLIT distance="300" swimtime="00:04:21.26" />
                    <SPLIT distance="350" swimtime="00:05:01.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-06-16" firstname="Paweł" gender="M" lastname="WITKOWSKI" nation="POL" athleteid="101729">
              <RESULTS>
                <RESULT eventid="98956" points="427" reactiontime="+88" swimtime="00:02:48.58" resultid="101730" heatid="105202" lane="6" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.42" />
                    <SPLIT distance="100" swimtime="00:01:20.47" />
                    <SPLIT distance="150" swimtime="00:02:04.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="460" reactiontime="+90" swimtime="00:01:15.73" resultid="101731" heatid="105255" lane="6" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="298" reactiontime="+83" swimtime="00:01:17.72" resultid="101732" heatid="105284" lane="7" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="517" reactiontime="+91" swimtime="00:00:33.22" resultid="101733" heatid="105359" lane="3" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-09-01" firstname="Andrzej" gender="M" lastname="CIEŚLIŃSKI" nation="POL" athleteid="101734">
              <RESULTS>
                <RESULT eventid="98798" points="237" reactiontime="+89" swimtime="00:00:33.77" resultid="101735" heatid="105129" lane="9" entrytime="00:00:33.20" />
                <RESULT eventid="98988" points="206" reactiontime="+76" swimtime="00:01:19.31" resultid="101736" heatid="105216" lane="8" entrytime="00:01:18.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.21" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="04" eventid="99218" reactiontime="+65" status="DSQ" swimtime="00:00:00.00" resultid="101737" heatid="105298" lane="7" entrytime="00:02:50.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.58" />
                    <SPLIT distance="100" swimtime="00:01:30.34" />
                    <SPLIT distance="150" swimtime="00:02:24.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-02-29" firstname="Jan" gender="M" lastname="BOBOLI" nation="POL" swrid="4754700" athleteid="101738">
              <RESULTS>
                <RESULT eventid="98798" points="179" reactiontime="+95" swimtime="00:00:37.07" resultid="101739" heatid="105126" lane="3" entrytime="00:00:36.00" />
                <RESULT eventid="98924" points="62" reactiontime="+84" swimtime="00:01:00.50" resultid="101740" heatid="105182" lane="9" entrytime="00:00:50.00" />
                <RESULT eventid="98988" points="130" reactiontime="+96" swimtime="00:01:32.41" resultid="101741" heatid="105214" lane="3" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="140" reactiontime="+88" swimtime="00:00:43.15" resultid="101742" heatid="105267" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="99425" points="47" reactiontime="+114" swimtime="00:01:13.61" resultid="101743" heatid="105351" lane="2" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-08-01" firstname="Edyta" gender="F" lastname="OLSZEWSKA" nation="POL" swrid="4754701" athleteid="101744">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="98940" points="367" swimtime="00:03:14.13" resultid="101745" heatid="105194" lane="7" entrytime="00:03:12.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.46" />
                    <SPLIT distance="100" swimtime="00:01:33.57" />
                    <SPLIT distance="150" swimtime="00:02:23.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="354" reactiontime="+81" swimtime="00:01:30.95" resultid="101746" heatid="105247" lane="1" entrytime="00:01:28.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="278" swimtime="00:02:52.99" resultid="101747" heatid="105292" lane="7" entrytime="00:02:47.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                    <SPLIT distance="100" swimtime="00:01:25.54" />
                    <SPLIT distance="150" swimtime="00:02:10.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="330" reactiontime="+82" swimtime="00:00:42.63" resultid="101748" heatid="105349" lane="7" entrytime="00:00:39.76" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-02-17" firstname="Piotr" gender="M" lastname="BARSKI" nation="POL" swrid="4595751" athleteid="101749">
              <RESULTS>
                <RESULT eventid="98798" points="431" reactiontime="+87" swimtime="00:00:27.67" resultid="101750" heatid="105142" lane="1" entrytime="00:00:26.00" />
                <RESULT eventid="98956" points="386" reactiontime="+86" swimtime="00:02:54.39" resultid="101751" heatid="105196" lane="4" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.07" />
                    <SPLIT distance="100" swimtime="00:01:25.25" />
                    <SPLIT distance="150" swimtime="00:02:10.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="459" reactiontime="+87" swimtime="00:01:00.81" resultid="101752" heatid="105227" lane="0" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="422" reactiontime="+89" swimtime="00:01:17.89" resultid="101753" heatid="105258" lane="0" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="445" reactiontime="+64" swimtime="00:00:34.92" resultid="101754" heatid="105362" lane="8" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-08-05" firstname="Tomasz" gender="M" lastname="BIELAN" nation="POL" athleteid="101755">
              <RESULTS>
                <RESULT eventid="98988" points="234" reactiontime="+96" swimtime="00:01:16.12" resultid="101756" heatid="105216" lane="5" entrytime="00:01:15.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="223" reactiontime="+84" swimtime="00:00:36.96" resultid="101757" heatid="105268" lane="6" entrytime="00:00:36.38" />
                <RESULT eventid="99218" points="184" reactiontime="+93" swimtime="00:02:59.05" resultid="101758" heatid="105297" lane="7" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                    <SPLIT distance="100" swimtime="00:01:25.37" />
                    <SPLIT distance="150" swimtime="00:02:14.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-13" firstname="Stanisław" gender="M" lastname="KOZAK" nation="POL" swrid="4992669" athleteid="101759">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="101760" heatid="105130" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="98956" points="468" reactiontime="+84" swimtime="00:02:43.48" resultid="101761" heatid="105204" lane="8" entrytime="00:02:40.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.38" />
                    <SPLIT distance="100" swimtime="00:01:18.46" />
                    <SPLIT distance="150" swimtime="00:02:01.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="573" reactiontime="+77" swimtime="00:01:10.38" resultid="101762" heatid="105258" lane="8" entrytime="00:01:10.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="101763" heatid="105274" lane="8" entrytime="00:00:29.84" />
                <RESULT eventid="99425" points="602" reactiontime="+92" swimtime="00:00:31.57" resultid="101764" heatid="105362" lane="3" entrytime="00:00:31.21" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-10-04" firstname="Maciej" gender="M" lastname="SZYMAŃSKI" nation="POL" athleteid="101765">
              <RESULTS>
                <RESULT eventid="98798" points="574" reactiontime="+77" swimtime="00:00:25.15" resultid="101766" heatid="105143" lane="7" entrytime="00:00:24.99" />
                <RESULT eventid="98891" status="WDR" swimtime="00:00:00.00" resultid="101767" entrytime="00:21:00.00" />
                <RESULT eventid="99170" points="507" reactiontime="+83" swimtime="00:00:28.12" resultid="101768" heatid="105276" lane="9" entrytime="00:00:27.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-10-17" firstname="Waldemar" gender="M" lastname="DE MAKAY" nation="POL" athleteid="101769">
              <RESULTS>
                <RESULT eventid="98798" points="262" reactiontime="+113" swimtime="00:00:32.64" resultid="101770" heatid="105130" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="98891" points="240" swimtime="00:23:20.89" resultid="101771" heatid="105422" lane="0" entrytime="00:22:52.00" />
                <RESULT eventid="98924" points="198" swimtime="00:00:41.24" resultid="101772" heatid="105185" lane="9" entrytime="00:00:40.00" />
                <RESULT eventid="98988" points="262" reactiontime="+112" swimtime="00:01:13.25" resultid="101773" heatid="105218" lane="0" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="221" reactiontime="+106" swimtime="00:02:48.51" resultid="101774" heatid="105299" lane="9" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                    <SPLIT distance="100" swimtime="00:01:19.00" />
                    <SPLIT distance="150" swimtime="00:02:04.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="172" reactiontime="+77" swimtime="00:03:20.89" resultid="101775" heatid="105338" lane="5" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.57" />
                    <SPLIT distance="100" swimtime="00:01:38.98" />
                    <SPLIT distance="150" swimtime="00:02:30.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="234" reactiontime="+120" swimtime="00:05:56.70" resultid="101776" heatid="106063" lane="1" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.65" />
                    <SPLIT distance="100" swimtime="00:01:23.82" />
                    <SPLIT distance="150" swimtime="00:02:09.52" />
                    <SPLIT distance="200" swimtime="00:02:56.24" />
                    <SPLIT distance="250" swimtime="00:03:42.43" />
                    <SPLIT distance="300" swimtime="00:04:29.04" />
                    <SPLIT distance="350" swimtime="00:05:14.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-10" firstname="Michał" gender="M" lastname="RUDZIŃSKI" nation="POL" swrid="4934041" athleteid="101777">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="101778" heatid="105126" lane="1" entrytime="00:00:36.84" />
                <RESULT eventid="98830" points="148" reactiontime="+101" swimtime="00:03:35.47" resultid="101779" heatid="105150" lane="8" entrytime="00:03:47.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.67" />
                    <SPLIT distance="100" swimtime="00:01:48.82" />
                    <SPLIT distance="150" swimtime="00:02:44.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98956" points="219" reactiontime="+118" swimtime="00:03:30.68" resultid="101780" heatid="105199" lane="6" entrytime="00:03:31.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.62" />
                    <SPLIT distance="100" swimtime="00:01:39.07" />
                    <SPLIT distance="150" swimtime="00:02:35.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" status="DNS" swimtime="00:00:00.00" resultid="101781" heatid="105231" lane="3" />
                <RESULT eventid="99091" points="225" reactiontime="+108" swimtime="00:01:36.07" resultid="101782" heatid="105251" lane="7" entrytime="00:01:38.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="144" reactiontime="+133" swimtime="00:07:44.40" resultid="101783" heatid="106047" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.45" />
                    <SPLIT distance="100" swimtime="00:01:55.56" />
                    <SPLIT distance="150" swimtime="00:03:04.15" />
                    <SPLIT distance="200" swimtime="00:04:09.50" />
                    <SPLIT distance="250" swimtime="00:05:04.06" />
                    <SPLIT distance="300" swimtime="00:05:59.67" />
                    <SPLIT distance="350" swimtime="00:06:53.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="94" reactiontime="+109" swimtime="00:01:49.37" resultid="101784" heatid="105325" lane="6" entrytime="00:01:58.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="235" reactiontime="+98" swimtime="00:00:43.20" resultid="101785" heatid="105354" lane="9" entrytime="00:00:44.32" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-10-23" firstname="Agata" gender="F" lastname="NYKOWSKA" nation="POL" athleteid="101786">
              <RESULTS>
                <RESULT eventid="98907" points="155" reactiontime="+94" swimtime="00:00:50.36" resultid="101787" heatid="105174" lane="8" entrytime="00:00:47.00" />
                <RESULT eventid="98972" points="229" swimtime="00:01:25.00" resultid="101788" heatid="105207" lane="8" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="142" reactiontime="+83" swimtime="00:01:51.15" resultid="101789" heatid="105278" lane="8" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="196" reactiontime="+102" swimtime="00:06:51.31" resultid="101790" heatid="106056" lane="2" entrytime="00:06:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.94" />
                    <SPLIT distance="100" swimtime="00:01:36.21" />
                    <SPLIT distance="150" swimtime="00:02:28.94" />
                    <SPLIT distance="200" swimtime="00:03:21.99" />
                    <SPLIT distance="250" swimtime="00:04:13.96" />
                    <SPLIT distance="300" swimtime="00:05:07.05" />
                    <SPLIT distance="350" swimtime="00:06:00.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-04" firstname="Jan" gender="M" lastname="GROCHOWICZ" nation="POL" athleteid="101791">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="101792" heatid="105134" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="98988" points="281" reactiontime="+97" swimtime="00:01:11.60" resultid="101793" heatid="105218" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="101794" heatid="105265" lane="7" />
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="101795" heatid="105298" lane="9" entrytime="00:02:55.00" />
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="101796" entrytime="00:06:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-30" firstname="Monika" gender="F" lastname="JARECKA-SKORYKOW" nation="POL" swrid="4992672" athleteid="101797">
              <RESULTS>
                <RESULT eventid="98777" points="445" reactiontime="+84" swimtime="00:00:31.08" resultid="101798" heatid="105119" lane="5" entrytime="00:00:31.46" entrycourse="SCM" />
                <RESULT eventid="98814" points="348" reactiontime="+88" swimtime="00:02:59.25" resultid="101799" heatid="105145" lane="5" entrytime="00:03:12.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                    <SPLIT distance="100" swimtime="00:01:26.01" />
                    <SPLIT distance="150" swimtime="00:02:15.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="368" reactiontime="+81" swimtime="00:03:14.09" resultid="101800" heatid="105194" lane="1" entrytime="00:03:13.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.61" />
                    <SPLIT distance="100" swimtime="00:01:31.15" />
                    <SPLIT distance="150" swimtime="00:02:22.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="393" reactiontime="+78" swimtime="00:01:27.78" resultid="101801" heatid="105247" lane="9" entrytime="00:01:29.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="378" reactiontime="+74" swimtime="00:00:34.67" resultid="101802" heatid="105263" lane="9" entrytime="00:00:34.98" />
                <RESULT eventid="99409" points="427" reactiontime="+88" swimtime="00:00:39.12" resultid="101803" heatid="105349" lane="2" entrytime="00:00:39.66" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-05-15" firstname="Michał" gender="M" lastname="WETOSZKA" nation="POL" athleteid="101804">
              <RESULTS>
                <RESULT eventid="98924" points="159" reactiontime="+79" swimtime="00:00:44.33" resultid="101805" heatid="105184" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="98988" points="193" reactiontime="+85" swimtime="00:01:21.13" resultid="101806" heatid="105217" lane="9" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="170" reactiontime="+95" swimtime="00:00:40.47" resultid="101807" heatid="105266" lane="5" entrytime="00:00:42.00" />
                <RESULT eventid="99218" points="160" reactiontime="+97" swimtime="00:03:07.66" resultid="101808" heatid="105297" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.72" />
                    <SPLIT distance="100" swimtime="00:01:26.58" />
                    <SPLIT distance="150" swimtime="00:02:18.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-08-12" firstname="Jakub" gender="M" lastname="SZULC" nation="POL" swrid="4992670" athleteid="101809">
              <RESULTS>
                <RESULT eventid="98988" points="421" reactiontime="+79" swimtime="00:01:02.57" resultid="101810" heatid="105221" lane="6" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="409" reactiontime="+86" swimtime="00:00:30.21" resultid="101811" heatid="105269" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="99218" points="349" reactiontime="+80" swimtime="00:02:24.79" resultid="101812" heatid="105300" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                    <SPLIT distance="100" swimtime="00:01:10.84" />
                    <SPLIT distance="150" swimtime="00:01:48.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="101813" entrytime="00:05:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-12-16" firstname="Przemysław" gender="M" lastname="WOŁOSZ" nation="POL" swrid="4992659" athleteid="101814">
              <RESULTS>
                <RESULT eventid="98924" status="DNS" swimtime="00:00:00.00" resultid="101815" heatid="105180" lane="9" />
                <RESULT eventid="99091" points="277" reactiontime="+81" swimtime="00:01:29.68" resultid="101816" heatid="105253" lane="8" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="273" reactiontime="+93" swimtime="00:00:34.55" resultid="101817" heatid="105267" lane="5" entrytime="00:00:39.00" />
                <RESULT eventid="99186" points="170" reactiontime="+85" swimtime="00:01:33.63" resultid="101818" heatid="105283" lane="4" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="203" reactiontime="+100" swimtime="00:01:24.72" resultid="101819" heatid="105324" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-09" firstname="Tomasz" gender="M" lastname="MAKOMASKI" nation="POL" swrid="4992665" athleteid="101820">
              <RESULTS>
                <RESULT eventid="98798" points="432" reactiontime="+89" swimtime="00:00:27.66" resultid="101821" heatid="105139" lane="3" entrytime="00:00:27.44" />
                <RESULT eventid="98956" points="357" reactiontime="+91" swimtime="00:02:59.00" resultid="101822" heatid="105203" lane="3" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.44" />
                    <SPLIT distance="100" swimtime="00:01:27.49" />
                    <SPLIT distance="150" swimtime="00:02:14.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="418" reactiontime="+75" swimtime="00:01:02.70" resultid="101823" heatid="105224" lane="9" entrytime="00:01:02.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="423" reactiontime="+77" swimtime="00:01:17.82" resultid="101824" heatid="105257" lane="7" entrytime="00:01:16.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="351" reactiontime="+82" swimtime="00:00:31.77" resultid="101825" heatid="105271" lane="6" entrytime="00:00:31.55" />
                <RESULT eventid="99361" points="312" reactiontime="+91" swimtime="00:01:13.41" resultid="101826" heatid="105330" lane="0" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="467" reactiontime="+78" swimtime="00:00:34.36" resultid="101827" heatid="105360" lane="9" entrytime="00:00:35.07" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-04-17" firstname="Andrzej" gender="M" lastname="SKORYKOW" nation="POL" swrid="4270349" athleteid="101828">
              <RESULTS>
                <RESULT eventid="98798" points="458" reactiontime="+79" swimtime="00:00:27.11" resultid="101829" heatid="105139" lane="1" entrytime="00:00:27.50" />
                <RESULT eventid="98830" points="446" reactiontime="+87" swimtime="00:02:29.14" resultid="101830" heatid="105156" lane="4" entrytime="00:02:32.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                    <SPLIT distance="100" swimtime="00:01:09.56" />
                    <SPLIT distance="150" swimtime="00:01:55.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="472" reactiontime="+67" swimtime="00:00:30.86" resultid="101831" heatid="105189" lane="6" entrytime="00:00:30.80" />
                <RESULT eventid="99020" points="427" reactiontime="+92" swimtime="00:02:28.04" resultid="101832" heatid="105236" lane="6" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                    <SPLIT distance="100" swimtime="00:01:10.03" />
                    <SPLIT distance="150" swimtime="00:01:48.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="477" reactiontime="+70" swimtime="00:00:28.69" resultid="101833" heatid="105275" lane="9" entrytime="00:00:28.20" />
                <RESULT eventid="99218" points="450" reactiontime="+88" swimtime="00:02:13.09" resultid="101834" heatid="105304" lane="0" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                    <SPLIT distance="100" swimtime="00:01:06.47" />
                    <SPLIT distance="150" swimtime="00:01:40.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="471" reactiontime="+75" swimtime="00:01:04.01" resultid="101835" heatid="105330" lane="4" entrytime="00:01:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" status="DNS" swimtime="00:00:00.00" resultid="101836" heatid="106060" lane="7" entrytime="00:04:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-07-26" firstname="Anna" gender="F" lastname="SZEMBERG" nation="POL" swrid="4302692" athleteid="101837">
              <RESULTS>
                <RESULT eventid="98777" points="85" swimtime="00:00:53.88" resultid="101838" heatid="105114" lane="7" entrytime="00:00:42.47" entrycourse="LCM" />
                <RESULT eventid="98863" points="105" swimtime="00:17:25.67" resultid="101839" heatid="105406" lane="6" entrytime="00:17:59.00" />
                <RESULT eventid="98907" status="DNS" swimtime="00:00:00.00" resultid="101840" heatid="105172" lane="6" entrytime="00:01:59.00" />
                <RESULT eventid="98972" points="82" swimtime="00:01:59.40" resultid="101841" heatid="105206" lane="0" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="81" swimtime="00:04:20.61" resultid="101842" heatid="105289" lane="2" entrytime="00:04:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.75" />
                    <SPLIT distance="100" swimtime="00:02:08.27" />
                    <SPLIT distance="150" swimtime="00:03:16.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="93" swimtime="00:08:46.12" resultid="101843" heatid="106057" lane="7" entrytime="00:08:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.69" />
                    <SPLIT distance="100" swimtime="00:02:05.29" />
                    <SPLIT distance="150" swimtime="00:03:13.31" />
                    <SPLIT distance="200" swimtime="00:04:21.33" />
                    <SPLIT distance="250" swimtime="00:05:28.93" />
                    <SPLIT distance="300" swimtime="00:06:36.32" />
                    <SPLIT distance="350" swimtime="00:07:42.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-05-31" firstname="Katharina" gender="F" lastname="THUMEYER" nation="POL" athleteid="101844">
              <RESULTS>
                <RESULT eventid="98777" points="230" reactiontime="+93" swimtime="00:00:38.73" resultid="101845" heatid="105115" lane="2" entrytime="00:00:39.00" />
                <RESULT eventid="98863" status="DNS" swimtime="00:00:00.00" resultid="101846" heatid="105406" lane="5" entrytime="00:15:00.00" />
                <RESULT eventid="98907" status="DNS" swimtime="00:00:00.00" resultid="101847" heatid="105174" lane="9" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-13" firstname="Agnieszka" gender="F" lastname="MAZURKIEWICZ" nation="POL" swrid="4992662" athleteid="101848">
              <RESULTS>
                <RESULT eventid="98777" points="318" reactiontime="+97" swimtime="00:00:34.74" resultid="101849" heatid="105116" lane="5" entrytime="00:00:35.89" entrycourse="SCM" />
                <RESULT eventid="98972" points="286" reactiontime="+97" swimtime="00:01:18.95" resultid="101850" heatid="105207" lane="3" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="304" reactiontime="+94" swimtime="00:00:37.27" resultid="101851" heatid="105261" lane="1" entrytime="00:00:39.57" />
                <RESULT eventid="99202" points="272" reactiontime="+97" swimtime="00:02:54.36" resultid="101852" heatid="105291" lane="2" entrytime="00:02:58.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.48" />
                    <SPLIT distance="100" swimtime="00:01:25.11" />
                    <SPLIT distance="150" swimtime="00:02:11.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="248" reactiontime="+90" swimtime="00:06:20.42" resultid="101853" heatid="106056" lane="6" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.84" />
                    <SPLIT distance="100" swimtime="00:01:31.44" />
                    <SPLIT distance="150" swimtime="00:02:20.05" />
                    <SPLIT distance="200" swimtime="00:03:08.85" />
                    <SPLIT distance="250" swimtime="00:03:57.82" />
                    <SPLIT distance="300" swimtime="00:04:46.60" />
                    <SPLIT distance="350" swimtime="00:05:35.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-24" firstname="Jan" gender="M" lastname="PFITZNER" nation="POL" swrid="4992671" athleteid="101854">
              <RESULTS>
                <RESULT eventid="98798" points="473" reactiontime="+73" swimtime="00:00:26.83" resultid="101855" heatid="105142" lane="9" entrytime="00:00:26.49" />
                <RESULT eventid="98924" points="438" reactiontime="+88" swimtime="00:00:31.64" resultid="101856" heatid="105180" lane="0" />
                <RESULT eventid="98988" points="503" reactiontime="+78" swimtime="00:00:58.96" resultid="101857" heatid="105226" lane="1" entrytime="00:00:59.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="462" reactiontime="+76" swimtime="00:00:29.01" resultid="101858" heatid="105274" lane="4" entrytime="00:00:28.49" />
                <RESULT eventid="99218" points="378" reactiontime="+73" swimtime="00:02:21.07" resultid="101859" heatid="105304" lane="7" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.84" />
                    <SPLIT distance="100" swimtime="00:01:09.12" />
                    <SPLIT distance="150" swimtime="00:01:45.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="377" reactiontime="+87" swimtime="00:05:04.40" resultid="101860" heatid="106060" lane="3" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                    <SPLIT distance="100" swimtime="00:01:13.66" />
                    <SPLIT distance="150" swimtime="00:01:53.44" />
                    <SPLIT distance="200" swimtime="00:02:33.53" />
                    <SPLIT distance="250" swimtime="00:03:11.00" />
                    <SPLIT distance="300" swimtime="00:03:49.16" />
                    <SPLIT distance="350" swimtime="00:04:26.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="5">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="99059" points="529" reactiontime="+85" swimtime="00:01:55.51" resultid="101872" heatid="105242" lane="4" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                    <SPLIT distance="100" swimtime="00:01:03.37" />
                    <SPLIT distance="150" swimtime="00:01:31.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101854" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="101759" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="101724" number="3" reactiontime="+16" />
                    <RELAYPOSITION athleteid="101765" number="4" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="6">
              <RESULTS>
                <RESULT eventid="99059" points="461" reactiontime="+85" swimtime="00:02:00.92" resultid="101873" heatid="105242" lane="3" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                    <SPLIT distance="100" swimtime="00:01:04.83" />
                    <SPLIT distance="150" swimtime="00:01:34.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101695" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="101729" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="101828" number="3" reactiontime="+72" />
                    <RELAYPOSITION athleteid="101749" number="4" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="7">
              <RESULTS>
                <RESULT eventid="99059" points="417" reactiontime="+71" swimtime="00:02:05.05" resultid="101874" heatid="105242" lane="9" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                    <SPLIT distance="100" swimtime="00:01:04.31" />
                    <SPLIT distance="150" swimtime="00:01:34.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101644" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="101820" number="2" />
                    <RELAYPOSITION athleteid="101809" number="3" reactiontime="+64" />
                    <RELAYPOSITION athleteid="101791" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="9">
              <RESULTS>
                <RESULT eventid="99250" points="544" reactiontime="+85" swimtime="00:01:43.92" resultid="101876" heatid="105311" lane="4" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.82" />
                    <SPLIT distance="100" swimtime="00:00:51.48" />
                    <SPLIT distance="150" swimtime="00:01:17.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101765" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="101759" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="101724" number="3" reactiontime="+9" />
                    <RELAYPOSITION athleteid="101854" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="10">
              <RESULTS>
                <RESULT eventid="99250" points="446" reactiontime="+93" swimtime="00:01:51.03" resultid="101877" heatid="105311" lane="3" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.72" />
                    <SPLIT distance="100" swimtime="00:00:55.66" />
                    <SPLIT distance="150" swimtime="00:01:24.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101695" number="1" reactiontime="+93" />
                    <RELAYPOSITION athleteid="101820" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="101597" number="3" reactiontime="+28" />
                    <RELAYPOSITION athleteid="101828" number="4" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="11">
              <RESULTS>
                <RESULT comment="04/ 2 zmiana" eventid="99250" reactiontime="+83" status="DSQ" swimtime="00:00:00.00" resultid="101878" heatid="105309" lane="5" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.93" />
                    <SPLIT distance="100" swimtime="00:01:04.67" />
                    <SPLIT distance="150" swimtime="00:01:40.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101630" number="1" reactiontime="+83" status="DSQ" />
                    <RELAYPOSITION athleteid="101734" number="2" reactiontime="-7" status="DSQ" />
                    <RELAYPOSITION athleteid="101738" number="3" reactiontime="+5" status="DSQ" />
                    <RELAYPOSITION athleteid="101804" number="4" reactiontime="+72" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="15">
              <RESULTS>
                <RESULT eventid="99059" status="DNS" swimtime="00:00:00.00" resultid="101882" heatid="105240" lane="3" entrytime="00:02:30.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101675" number="1" />
                    <RELAYPOSITION athleteid="101711" number="2" />
                    <RELAYPOSITION athleteid="101738" number="3" />
                    <RELAYPOSITION athleteid="101630" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="3">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="99036" points="407" reactiontime="+81" swimtime="00:02:23.02" resultid="101870" heatid="105238" lane="4" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.78" />
                    <SPLIT distance="100" swimtime="00:01:18.53" />
                    <SPLIT distance="150" swimtime="00:01:49.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101702" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="101797" number="2" reactiontime="+73" />
                    <RELAYPOSITION athleteid="101707" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="101590" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" number="4">
              <RESULTS>
                <RESULT eventid="99036" points="235" reactiontime="+90" swimtime="00:02:51.80" resultid="101871" heatid="105237" lane="4" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.82" />
                    <SPLIT distance="100" swimtime="00:01:37.41" />
                    <SPLIT distance="150" swimtime="00:02:15.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101786" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="101844" number="2" reactiontime="+30" />
                    <RELAYPOSITION athleteid="101848" number="3" reactiontime="+71" />
                    <RELAYPOSITION athleteid="101622" number="4" reactiontime="+75" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="8">
              <RESULTS>
                <RESULT eventid="99234" points="425" reactiontime="+87" swimtime="00:02:08.68" resultid="101875" heatid="105307" lane="5" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                    <SPLIT distance="100" swimtime="00:01:07.35" />
                    <SPLIT distance="150" swimtime="00:01:40.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101797" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="101848" number="2" reactiontime="+90" />
                    <RELAYPOSITION athleteid="101590" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="101707" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="289" reactiontime="+90" swimtime="00:02:08.33" resultid="101868" heatid="105160" lane="1" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.76" />
                    <SPLIT distance="100" swimtime="00:01:06.36" />
                    <SPLIT distance="150" swimtime="00:01:41.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101648" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="101622" number="2" reactiontime="+73" />
                    <RELAYPOSITION athleteid="101848" number="3" />
                    <RELAYPOSITION athleteid="101820" number="4" reactiontime="+65" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="98846" points="391" reactiontime="+75" swimtime="00:01:55.99" resultid="101869" heatid="105161" lane="4" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.15" />
                    <SPLIT distance="100" swimtime="00:01:05.53" />
                    <SPLIT distance="150" swimtime="00:01:31.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101590" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="101797" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="101854" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="101765" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="12">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="99441" points="414" reactiontime="+88" swimtime="00:02:05.27" resultid="101879" heatid="105365" lane="4" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                    <SPLIT distance="100" swimtime="00:01:03.80" />
                    <SPLIT distance="150" swimtime="00:01:34.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101854" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="101759" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="101707" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="101797" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="13">
              <RESULTS>
                <RESULT eventid="99441" points="329" reactiontime="+71" swimtime="00:02:15.24" resultid="101880" heatid="105365" lane="8" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                    <SPLIT distance="100" swimtime="00:01:04.80" />
                    <SPLIT distance="150" swimtime="00:01:40.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101644" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="101820" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="101590" number="3" />
                    <RELAYPOSITION athleteid="101848" number="4" reactiontime="+65" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="14">
              <RESULTS>
                <RESULT eventid="98846" points="213" reactiontime="+100" swimtime="00:02:21.97" resultid="101881" heatid="105159" lane="6" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.80" />
                    <SPLIT distance="100" swimtime="00:01:08.51" />
                    <SPLIT distance="150" swimtime="00:01:46.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101673" number="1" reactiontime="+100" />
                    <RELAYPOSITION athleteid="101615" number="2" reactiontime="+65" />
                    <RELAYPOSITION athleteid="101844" number="3" reactiontime="+4" />
                    <RELAYPOSITION athleteid="101738" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="SLA" clubid="100667" name="Weteran  Zabrze">
          <CONTACT city="ZABRZE" email="WETERANZABRZE@OP.PL" name="BOSOWSKI  WŁODZIMIERZ" street="ŚW.JANA  4AI4" zip="41803" />
          <ATHLETES>
            <ATHLETE birthdate="1950-10-05" firstname="Barbara" gender="F" lastname="BRENDLER" nation="POL" license="502611100005" swrid="4269850" athleteid="100668">
              <RESULTS>
                <RESULT eventid="98777" points="200" reactiontime="+94" swimtime="00:00:40.52" resultid="100669" heatid="105114" lane="5" entrytime="00:00:40.17" entrycourse="LCM" />
                <RESULT eventid="98972" points="160" reactiontime="+99" swimtime="00:01:35.76" resultid="100670" heatid="105206" lane="5" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" status="DNS" swimtime="00:00:00.00" resultid="100671" heatid="105289" lane="4" entrytime="00:03:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-11" firstname="Jan" gender="M" lastname="BARUCHA" nation="POL" license="502611200008" athleteid="100672">
              <RESULTS>
                <RESULT eventid="98924" reactiontime="+87" status="DNS" swimtime="00:00:00.00" resultid="100673" heatid="105185" lane="0" entrytime="00:00:39.80" />
                <RESULT eventid="99186" status="DNS" swimtime="00:00:00.00" resultid="100674" heatid="105284" lane="1" entrytime="00:01:24.00" />
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="100675" heatid="105338" lane="4" entrytime="00:03:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-02-25" firstname="Bernard" gender="M" lastname="POLOCZEK" nation="POL" license="502611200004" swrid="4792004" athleteid="100676">
              <RESULTS>
                <RESULT eventid="98924" points="173" reactiontime="+69" swimtime="00:00:43.09" resultid="100677" heatid="105183" lane="5" entrytime="00:00:42.41" />
                <RESULT eventid="99186" points="141" reactiontime="+72" swimtime="00:01:39.58" resultid="100678" heatid="105282" lane="3" entrytime="00:01:40.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="128" reactiontime="+74" swimtime="00:03:41.78" resultid="100679" heatid="105337" lane="2" entrytime="00:03:46.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.90" />
                    <SPLIT distance="100" swimtime="00:01:45.52" />
                    <SPLIT distance="150" swimtime="00:02:43.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-05-27" firstname="Dawid" gender="M" lastname="MUSZALA" nation="POL" swrid="4954168" athleteid="100680">
              <RESULTS>
                <RESULT eventid="98891" points="180" swimtime="00:25:40.81" resultid="100681" heatid="105421" lane="8" entrytime="00:21:20.00" />
                <RESULT eventid="99218" points="226" reactiontime="+62" swimtime="00:02:47.44" resultid="100682" heatid="105299" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.07" />
                    <SPLIT distance="100" swimtime="00:01:17.90" />
                    <SPLIT distance="150" swimtime="00:02:03.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="208" reactiontime="+68" swimtime="00:06:11.20" resultid="100683" heatid="106063" lane="7" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.26" />
                    <SPLIT distance="100" swimtime="00:01:22.95" />
                    <SPLIT distance="150" swimtime="00:02:07.28" />
                    <SPLIT distance="200" swimtime="00:02:54.13" />
                    <SPLIT distance="250" swimtime="00:03:43.01" />
                    <SPLIT distance="300" swimtime="00:04:32.70" />
                    <SPLIT distance="350" swimtime="00:05:23.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-12-02" firstname="Renata" gender="F" lastname="BASTEK" nation="POL" license="502611100001" swrid="4223066" athleteid="100684">
              <RESULTS>
                <RESULT eventid="98777" points="278" reactiontime="+87" swimtime="00:00:36.32" resultid="100685" heatid="105118" lane="2" entrytime="00:00:33.06" entrycourse="LCM" />
                <RESULT eventid="98907" points="214" reactiontime="+77" swimtime="00:00:45.18" resultid="100686" heatid="105175" lane="9" entrytime="00:00:43.00" />
                <RESULT eventid="98972" points="237" reactiontime="+91" swimtime="00:01:24.06" resultid="100687" heatid="105207" lane="2" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="186" reactiontime="+71" swimtime="00:01:41.67" resultid="100688" heatid="105278" lane="9" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.39" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99377" points="167" reactiontime="+76" swimtime="00:03:44.90" resultid="100689" heatid="105332" lane="3" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.75" />
                    <SPLIT distance="100" swimtime="00:01:50.83" />
                    <SPLIT distance="150" swimtime="00:02:49.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-07-16" firstname="Ewald" gender="M" lastname="BASTEK" nation="POL" license="502611200001" swrid="4188447" athleteid="100690">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="98891" points="164" swimtime="00:26:28.80" resultid="100691" heatid="105424" lane="1" entrytime="00:28:00.00" />
                <RESULT comment="Rekord Polski Masters" eventid="99218" points="155" reactiontime="+115" swimtime="00:03:09.81" resultid="100692" heatid="105296" lane="5" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.30" />
                    <SPLIT distance="100" swimtime="00:01:33.11" />
                    <SPLIT distance="150" swimtime="00:02:22.73" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99473" points="177" reactiontime="+110" swimtime="00:06:31.82" resultid="100693" heatid="106066" lane="4" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.76" />
                    <SPLIT distance="100" swimtime="00:01:33.72" />
                    <SPLIT distance="150" swimtime="00:02:23.88" />
                    <SPLIT distance="200" swimtime="00:03:14.82" />
                    <SPLIT distance="250" swimtime="00:04:04.16" />
                    <SPLIT distance="300" swimtime="00:04:54.57" />
                    <SPLIT distance="350" swimtime="00:05:45.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-28" firstname="Wiesław" gender="M" lastname="KORNICKI" nation="POL" license="502611200007" swrid="4137183" athleteid="100694">
              <RESULTS>
                <RESULT eventid="98798" points="265" reactiontime="+66" swimtime="00:00:32.55" resultid="100695" heatid="105131" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="98988" points="236" reactiontime="+83" swimtime="00:01:15.87" resultid="100696" heatid="105218" lane="9" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="243" reactiontime="+88" swimtime="00:00:35.91" resultid="100697" heatid="105269" lane="5" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-11-02" firstname="Beata" gender="F" lastname="SULEWSKA" nation="POL" license="502611100009" swrid="4792005" athleteid="100698">
              <RESULTS>
                <RESULT eventid="98814" status="DNS" swimtime="00:00:00.00" resultid="100699" heatid="105147" lane="6" entrytime="00:02:49.50" />
                <RESULT eventid="98863" points="445" reactiontime="+97" swimtime="00:10:46.64" resultid="100700" heatid="105404" lane="2" entrytime="00:10:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.46" />
                    <SPLIT distance="100" swimtime="00:01:13.97" />
                    <SPLIT distance="150" swimtime="00:01:53.48" />
                    <SPLIT distance="200" swimtime="00:02:33.67" />
                    <SPLIT distance="250" swimtime="00:03:14.03" />
                    <SPLIT distance="300" swimtime="00:03:54.87" />
                    <SPLIT distance="350" swimtime="00:04:35.84" />
                    <SPLIT distance="400" swimtime="00:05:16.97" />
                    <SPLIT distance="450" swimtime="00:05:58.00" />
                    <SPLIT distance="500" swimtime="00:06:39.43" />
                    <SPLIT distance="550" swimtime="00:07:20.94" />
                    <SPLIT distance="600" swimtime="00:08:02.54" />
                    <SPLIT distance="650" swimtime="00:08:44.24" />
                    <SPLIT distance="700" swimtime="00:09:25.35" />
                    <SPLIT distance="750" swimtime="00:10:06.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98940" points="406" reactiontime="+94" swimtime="00:03:07.78" resultid="100701" heatid="105194" lane="6" entrytime="00:03:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.89" />
                    <SPLIT distance="100" swimtime="00:01:29.90" />
                    <SPLIT distance="150" swimtime="00:02:18.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="402" reactiontime="+97" swimtime="00:01:27.15" resultid="100702" heatid="105247" lane="2" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.12" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99266" points="422" reactiontime="+98" swimtime="00:05:57.81" resultid="100703" heatid="106046" lane="5" entrytime="00:06:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                    <SPLIT distance="100" swimtime="00:01:19.44" />
                    <SPLIT distance="150" swimtime="00:02:10.67" />
                    <SPLIT distance="200" swimtime="00:02:59.09" />
                    <SPLIT distance="250" swimtime="00:03:47.54" />
                    <SPLIT distance="300" swimtime="00:04:37.34" />
                    <SPLIT distance="350" swimtime="00:05:18.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="442" reactiontime="+89" swimtime="00:05:13.93" resultid="100704" heatid="106054" lane="1" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                    <SPLIT distance="100" swimtime="00:01:14.35" />
                    <SPLIT distance="150" swimtime="00:01:53.96" />
                    <SPLIT distance="200" swimtime="00:02:33.95" />
                    <SPLIT distance="250" swimtime="00:03:14.00" />
                    <SPLIT distance="300" swimtime="00:03:54.49" />
                    <SPLIT distance="350" swimtime="00:04:34.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-11-29" firstname="Daniel" gender="M" lastname="FECICA" nation="POL" license="502611200002" swrid="4102523" athleteid="100705">
              <RESULTS>
                <RESULT eventid="98956" points="203" reactiontime="+112" swimtime="00:03:35.87" resultid="100706" heatid="105199" lane="2" entrytime="00:03:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.78" />
                    <SPLIT distance="100" swimtime="00:01:44.06" />
                    <SPLIT distance="150" swimtime="00:02:39.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="201" reactiontime="+102" swimtime="00:01:39.69" resultid="100707" heatid="105251" lane="2" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="126" reactiontime="+95" swimtime="00:00:44.73" resultid="100708" heatid="105266" lane="4" entrytime="00:00:42.00" />
                <RESULT eventid="99425" points="184" reactiontime="+107" swimtime="00:00:46.85" resultid="100709" heatid="105354" lane="2" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-03-12" firstname="Krystyna" gender="F" lastname="FECICA" nation="POL" license="502611100002" swrid="4102524" athleteid="100710">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="98940" points="183" reactiontime="+116" swimtime="00:04:04.68" resultid="100711" heatid="105192" lane="1" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.27" />
                    <SPLIT distance="100" swimtime="00:01:58.27" />
                    <SPLIT distance="150" swimtime="00:03:01.61" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="99089" points="187" reactiontime="+105" swimtime="00:01:52.37" resultid="100712" heatid="105244" lane="3" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="109" reactiontime="+115" swimtime="00:00:52.46" resultid="100713" heatid="105259" lane="2" entrytime="00:00:50.00" />
                <RESULT comment="Rekord Polski Masters" eventid="99409" points="183" reactiontime="+99" swimtime="00:00:51.87" resultid="100714" heatid="105345" lane="7" entrytime="00:00:52.50" />
                <RESULT comment="Rekord Polski Masters" eventid="99457" points="126" reactiontime="+108" swimtime="00:07:56.44" resultid="100715" heatid="106057" lane="2" entrytime="00:08:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.04" />
                    <SPLIT distance="100" swimtime="00:01:53.06" />
                    <SPLIT distance="150" swimtime="00:02:54.21" />
                    <SPLIT distance="200" swimtime="00:03:56.19" />
                    <SPLIT distance="250" swimtime="00:04:56.32" />
                    <SPLIT distance="300" swimtime="00:05:56.82" />
                    <SPLIT distance="350" swimtime="00:06:57.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-05-22" firstname="Włodzimierz" gender="M" lastname="BOSOWSKI" nation="POL" license="502611200005" swrid="4129761" athleteid="100716">
              <RESULTS>
                <RESULT eventid="98798" points="155" reactiontime="+100" swimtime="00:00:38.89" resultid="100717" heatid="105126" lane="9" entrytime="00:00:37.85" />
                <RESULT eventid="99170" points="93" reactiontime="+99" swimtime="00:00:49.34" resultid="100718" heatid="105267" lane="8" entrytime="00:00:40.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-05-21" firstname="Marek" gender="M" lastname="ROTHER" nation="POL" license="502611200009" swrid="4351633" athleteid="100719">
              <RESULTS>
                <RESULT eventid="98830" points="422" reactiontime="+82" swimtime="00:02:31.94" resultid="100720" heatid="105155" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                    <SPLIT distance="100" swimtime="00:01:09.94" />
                    <SPLIT distance="150" swimtime="00:01:55.77" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters, Rekord Polski Masters" eventid="98924" points="497" reactiontime="+70" swimtime="00:00:30.33" resultid="100721" heatid="105189" lane="4" entrytime="00:00:30.50" />
                <RESULT eventid="99186" points="500" reactiontime="+64" swimtime="00:01:05.42" resultid="100722" heatid="105288" lane="8" entrytime="00:01:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="100723" heatid="105303" lane="8" entrytime="00:02:15.00" />
                <RESULT eventid="99393" points="472" reactiontime="+72" swimtime="00:02:23.65" resultid="100724" heatid="105343" lane="1" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.76" />
                    <SPLIT distance="100" swimtime="00:01:10.49" />
                    <SPLIT distance="150" swimtime="00:01:47.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-05-03" firstname="Marta" gender="F" lastname="FRANK" nation="POL" license="502611100008" swrid="4967439" athleteid="100725">
              <RESULTS>
                <RESULT eventid="98777" points="401" reactiontime="+79" swimtime="00:00:32.16" resultid="100726" heatid="105118" lane="3" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="98907" points="420" reactiontime="+67" swimtime="00:00:36.11" resultid="100727" heatid="105178" lane="9" entrytime="00:00:35.90" />
                <RESULT eventid="99314" points="409" reactiontime="+71" swimtime="00:01:18.28" resultid="100728" heatid="105280" lane="7" entrytime="00:01:17.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="356" reactiontime="+71" swimtime="00:02:54.92" resultid="100729" heatid="105334" lane="6" entrytime="00:02:53.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.64" />
                    <SPLIT distance="100" swimtime="00:01:24.41" />
                    <SPLIT distance="150" swimtime="00:02:11.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="4">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="99059" points="176" reactiontime="+76" swimtime="00:02:46.42" resultid="100733" heatid="105240" lane="1" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.91" />
                    <SPLIT distance="100" swimtime="00:01:30.71" />
                    <SPLIT distance="150" swimtime="00:02:08.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100676" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="100705" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="100694" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="100690" number="4" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="6">
              <RESULTS>
                <RESULT eventid="99250" points="250" reactiontime="+91" swimtime="00:02:14.55" resultid="100735" heatid="105309" lane="1" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.59" />
                    <SPLIT distance="100" swimtime="00:01:15.65" />
                    <SPLIT distance="150" swimtime="00:01:43.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100676" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="100716" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="100719" number="3" reactiontime="+73" />
                    <RELAYPOSITION athleteid="100694" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="F" number="3">
              <RESULTS>
                <RESULT eventid="99036" points="214" reactiontime="+71" swimtime="00:02:57.06" resultid="100732" heatid="105238" lane="0" entrytime="00:02:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                    <SPLIT distance="100" swimtime="00:01:27.65" />
                    <SPLIT distance="150" swimtime="00:02:16.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100725" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="100710" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="100684" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="100668" number="4" reactiontime="+68" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="F" number="5">
              <RESULTS>
                <RESULT eventid="99234" points="225" reactiontime="+98" swimtime="00:02:38.93" resultid="100734" heatid="105306" lane="5" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.54" />
                    <SPLIT distance="100" swimtime="00:01:28.57" />
                    <SPLIT distance="150" swimtime="00:02:06.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100668" number="1" reactiontime="+98" />
                    <RELAYPOSITION athleteid="100710" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="100684" number="3" reactiontime="+74" />
                    <RELAYPOSITION athleteid="100725" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="146" reactiontime="+116" swimtime="00:02:40.96" resultid="100730" heatid="105159" lane="5" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                    <SPLIT distance="100" swimtime="00:01:24.16" />
                    <SPLIT distance="150" swimtime="00:02:02.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100684" number="1" reactiontime="+116" />
                    <RELAYPOSITION athleteid="100710" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="100705" number="3" reactiontime="+62" />
                    <RELAYPOSITION athleteid="100716" number="4" reactiontime="+87" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="98846" points="199" reactiontime="+97" swimtime="00:02:25.18" resultid="100731" heatid="105159" lane="3" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.19" />
                    <SPLIT distance="100" swimtime="00:01:17.65" />
                    <SPLIT distance="150" swimtime="00:01:51.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100668" number="1" reactiontime="+97" />
                    <RELAYPOSITION athleteid="100690" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="100725" number="3" reactiontime="+60" />
                    <RELAYPOSITION athleteid="100694" number="4" reactiontime="+66" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" number="7">
              <RESULTS>
                <RESULT eventid="99441" points="144" reactiontime="+73" swimtime="00:02:58.13" resultid="100736" heatid="105363" lane="5" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.01" />
                    <SPLIT distance="100" swimtime="00:01:37.12" />
                    <SPLIT distance="150" swimtime="00:02:21.63" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="100676" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="100710" number="2" reactiontime="+33" />
                    <RELAYPOSITION athleteid="100705" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="100684" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="LBS" clubid="101232" name="ZKS Drzonków">
          <CONTACT city="Świdnica" email="horbacz.marcin@wp.pl" name="Horbacz Marcin" phone="603672717" state="LBS" street="Buchałów 12c" zip="66-008" />
          <ATHLETES>
            <ATHLETE birthdate="1971-01-01" firstname="Piotr" gender="M" lastname="Barta" nation="POL" athleteid="101233">
              <RESULTS>
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="101234" heatid="105156" lane="7" entrytime="00:02:35.00" entrycourse="LCM" />
                <RESULT comment="Rekord Polski Masters" eventid="98956" points="479" reactiontime="+85" swimtime="00:02:42.30" resultid="101235" heatid="105204" lane="9" entrytime="00:02:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                    <SPLIT distance="100" swimtime="00:01:16.46" />
                    <SPLIT distance="150" swimtime="00:01:58.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="501" reactiontime="+92" swimtime="00:01:13.58" resultid="101236" heatid="105257" lane="2" entrytime="00:01:16.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" status="DNS" swimtime="00:00:00.00" resultid="101237" heatid="106053" lane="9" entrytime="00:05:40.00" entrycourse="LCM" />
                <RESULT eventid="99425" points="467" reactiontime="+77" swimtime="00:00:34.37" resultid="101238" heatid="105361" lane="8" entrytime="00:00:34.34" entrycourse="LCM" />
                <RESULT eventid="99473" points="440" reactiontime="+108" swimtime="00:04:49.27" resultid="101239" heatid="106061" lane="3" entrytime="00:04:57.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                    <SPLIT distance="100" swimtime="00:01:10.20" />
                    <SPLIT distance="150" swimtime="00:01:46.78" />
                    <SPLIT distance="200" swimtime="00:02:23.69" />
                    <SPLIT distance="250" swimtime="00:03:00.13" />
                    <SPLIT distance="300" swimtime="00:03:36.87" />
                    <SPLIT distance="350" swimtime="00:04:13.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="INDYWID." nation="POL" clubid="100963" name="Zawodnik niezrzeszony" shortname="niezrzeszony">
          <CONTACT name="ch" />
          <ATHLETES>
            <ATHLETE birthdate="1974-11-19" firstname="Judyta" gender="F" lastname="SOŁTYK" nation="POL" athleteid="100964">
              <RESULTS>
                <RESULT eventid="98814" points="370" reactiontime="+94" swimtime="00:02:55.57" resultid="100965" heatid="105144" lane="0" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.00" />
                    <SPLIT distance="100" swimtime="00:01:21.57" />
                    <SPLIT distance="150" swimtime="00:02:13.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98863" points="424" reactiontime="+101" swimtime="00:10:57.22" resultid="100966" heatid="105404" lane="1" entrytime="00:10:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                    <SPLIT distance="100" swimtime="00:01:14.82" />
                    <SPLIT distance="150" swimtime="00:01:54.78" />
                    <SPLIT distance="200" swimtime="00:02:35.71" />
                    <SPLIT distance="250" swimtime="00:03:16.86" />
                    <SPLIT distance="300" swimtime="00:03:58.59" />
                    <SPLIT distance="350" swimtime="00:04:40.20" />
                    <SPLIT distance="400" swimtime="00:05:22.37" />
                    <SPLIT distance="450" swimtime="00:06:04.40" />
                    <SPLIT distance="500" swimtime="00:06:46.63" />
                    <SPLIT distance="550" swimtime="00:07:28.68" />
                    <SPLIT distance="600" swimtime="00:08:10.98" />
                    <SPLIT distance="650" swimtime="00:08:53.01" />
                    <SPLIT distance="700" swimtime="00:09:35.06" />
                    <SPLIT distance="750" swimtime="00:10:16.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="380" reactiontime="+86" swimtime="00:00:34.59" resultid="100967" heatid="105263" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="99202" points="389" reactiontime="+90" swimtime="00:02:34.74" resultid="100968" heatid="105293" lane="5" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                    <SPLIT distance="100" swimtime="00:01:14.01" />
                    <SPLIT distance="150" swimtime="00:01:54.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-27" firstname="Michał" gender="M" lastname="KLUPA" nation="POL" swrid="4071939" athleteid="100969">
              <RESULTS>
                <RESULT eventid="98830" points="484" reactiontime="+80" swimtime="00:02:25.16" resultid="100970" heatid="105157" lane="5" entrytime="00:02:29.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.90" />
                    <SPLIT distance="100" swimtime="00:01:06.74" />
                    <SPLIT distance="150" swimtime="00:01:52.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="522" reactiontime="+70" swimtime="00:00:29.84" resultid="100971" heatid="105189" lane="1" entrytime="00:00:31.86" />
                <RESULT eventid="99186" points="500" reactiontime="+72" swimtime="00:01:05.44" resultid="100972" heatid="105287" lane="2" entrytime="00:01:09.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="470" reactiontime="+73" swimtime="00:02:23.92" resultid="100973" heatid="105342" lane="3" entrytime="00:02:31.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.87" />
                    <SPLIT distance="100" swimtime="00:01:10.56" />
                    <SPLIT distance="150" swimtime="00:01:47.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-06-11" firstname="Leszek" gender="M" lastname="SZYSZKA" nation="POL" athleteid="100974">
              <RESULTS>
                <RESULT eventid="98798" points="196" reactiontime="+124" swimtime="00:00:35.94" resultid="100975" heatid="105134" lane="7" entrytime="00:00:30.00" />
                <RESULT eventid="98988" points="189" reactiontime="+130" swimtime="00:01:21.69" resultid="100976" heatid="105217" lane="4" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-09-19" firstname="Zygmunt" gender="M" lastname="LEWANDOWSKI" nation="POL" swrid="4186953" athleteid="100977">
              <RESULTS>
                <RESULT eventid="98798" points="131" reactiontime="+93" swimtime="00:00:41.16" resultid="100978" heatid="105125" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="98891" points="99" swimtime="00:31:17.98" resultid="100979" heatid="105425" lane="4" entrytime="00:30:00.00" />
                <RESULT eventid="98988" points="116" reactiontime="+98" swimtime="00:01:36.14" resultid="100980" heatid="105214" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="108" reactiontime="+102" swimtime="00:07:40.99" resultid="100982" heatid="106066" lane="7" entrytime="00:07:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.71" />
                    <SPLIT distance="100" swimtime="00:01:47.58" />
                    <SPLIT distance="150" swimtime="00:02:48.84" />
                    <SPLIT distance="200" swimtime="00:03:49.07" />
                    <SPLIT distance="250" swimtime="00:04:48.81" />
                    <SPLIT distance="300" swimtime="00:05:47.75" />
                    <SPLIT distance="350" swimtime="00:06:46.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="101" reactiontime="+104" swimtime="00:03:38.67" resultid="104385" heatid="105296" lane="9" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.94" />
                    <SPLIT distance="100" swimtime="00:01:45.49" />
                    <SPLIT distance="150" swimtime="00:02:43.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-11-22" firstname="Marek" gender="M" lastname="PAŁYSA" nation="POL" swrid="4992690" athleteid="100983">
              <RESULTS>
                <RESULT eventid="98956" points="245" reactiontime="+99" swimtime="00:03:22.93" resultid="100984" heatid="105201" lane="0" entrytime="00:03:11.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.75" />
                    <SPLIT distance="100" swimtime="00:01:32.44" />
                    <SPLIT distance="150" swimtime="00:02:25.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="292" reactiontime="+84" swimtime="00:01:28.10" resultid="100985" heatid="105255" lane="7" entrytime="00:01:22.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="294" reactiontime="+88" swimtime="00:00:33.72" resultid="100986" heatid="105270" lane="8" entrytime="00:00:34.60" />
                <RESULT eventid="99425" points="337" reactiontime="+91" swimtime="00:00:38.30" resultid="100987" heatid="105360" lane="7" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-02-18" firstname="Kazimierz" gender="M" lastname="SINICKI" nation="POL" swrid="4754753" athleteid="100988">
              <RESULTS>
                <RESULT eventid="98798" points="341" reactiontime="+86" swimtime="00:00:29.91" resultid="100989" heatid="105133" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="98988" points="313" reactiontime="+83" swimtime="00:01:09.03" resultid="100990" heatid="105221" lane="9" entrytime="00:01:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="236" reactiontime="+90" swimtime="00:00:36.25" resultid="100991" heatid="105269" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="100992" heatid="105299" lane="2" entrytime="00:02:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-03-01" firstname="Marcin" gender="M" lastname="GÓRKA" nation="POL" swrid="4060962" athleteid="101001">
              <RESULTS>
                <RESULT eventid="98924" points="514" reactiontime="+78" swimtime="00:00:30.01" resultid="101002" heatid="105190" lane="0" entrytime="00:00:30.00" />
                <RESULT eventid="99170" points="554" reactiontime="+89" swimtime="00:00:27.30" resultid="101003" heatid="105275" lane="5" entrytime="00:00:27.50" />
                <RESULT eventid="99186" points="516" reactiontime="+64" swimtime="00:01:04.74" resultid="101004" heatid="105288" lane="7" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="525" reactiontime="+87" swimtime="00:01:01.74" resultid="101005" heatid="105331" lane="0" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="452" reactiontime="+49" swimtime="00:02:25.82" resultid="101006" heatid="105343" lane="0" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                    <SPLIT distance="100" swimtime="00:01:11.93" />
                    <SPLIT distance="150" swimtime="00:01:48.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-02" firstname="Janusz" gender="M" lastname="PLONKA" nation="POL" swrid="4754750" athleteid="101014">
              <RESULTS>
                <RESULT eventid="98830" points="62" reactiontime="+110" swimtime="00:04:47.61" resultid="101015" heatid="105148" lane="5" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.66" />
                    <SPLIT distance="100" swimtime="00:02:25.00" />
                    <SPLIT distance="150" swimtime="00:03:48.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="66" reactiontime="+85" swimtime="00:00:59.29" resultid="101016" heatid="105181" lane="0" entrytime="00:00:57.00" />
                <RESULT eventid="99020" points="35" reactiontime="+107" swimtime="00:05:40.87" resultid="101017" heatid="105231" lane="4" entrytime="00:05:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.24" />
                    <SPLIT distance="100" swimtime="00:02:33.88" />
                    <SPLIT distance="150" swimtime="00:04:10.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="62" reactiontime="+122" swimtime="00:00:56.50" resultid="101018" heatid="105265" lane="4" entrytime="00:00:53.00" />
                <RESULT eventid="99282" points="48" reactiontime="+115" swimtime="00:11:08.50" resultid="101019" heatid="106047" lane="4" entrytime="00:10:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.45" />
                    <SPLIT distance="100" swimtime="00:02:29.00" />
                    <SPLIT distance="150" swimtime="00:04:13.43" />
                    <SPLIT distance="200" swimtime="00:05:43.62" />
                    <SPLIT distance="250" swimtime="00:07:17.51" />
                    <SPLIT distance="300" swimtime="00:08:49.18" />
                    <SPLIT distance="350" swimtime="00:10:02.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="49" reactiontime="+118" swimtime="00:02:15.43" resultid="101020" heatid="105325" lane="0" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="84" reactiontime="+119" swimtime="00:01:00.82" resultid="101021" heatid="105351" lane="1" entrytime="00:01:02.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-04-24" firstname="Włodzimierz" gender="M" lastname="ZIELEZIŃSKI" nation="POL" swrid="4992697" athleteid="101026">
              <RESULTS>
                <RESULT eventid="98798" points="225" reactiontime="+110" swimtime="00:00:34.33" resultid="101027" heatid="105128" lane="8" entrytime="00:00:34.50" />
                <RESULT comment="Rekord Polski Masters" eventid="98891" status="DNS" swimtime="00:00:00.00" resultid="101028" heatid="105424" lane="2" entrytime="00:27:00.00" />
                <RESULT eventid="98924" points="187" reactiontime="+84" swimtime="00:00:41.98" resultid="101029" heatid="105183" lane="7" entrytime="00:00:43.00" />
                <RESULT eventid="98988" points="201" reactiontime="+121" swimtime="00:01:20.02" resultid="101030" heatid="105216" lane="2" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="156" reactiontime="+103" swimtime="00:01:36.44" resultid="101031" heatid="105283" lane="1" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="184" reactiontime="+106" swimtime="00:02:59.04" resultid="101032" heatid="105297" lane="8" entrytime="00:03:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                    <SPLIT distance="100" swimtime="00:01:24.28" />
                    <SPLIT distance="150" swimtime="00:02:12.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="147" reactiontime="+85" swimtime="00:03:31.85" resultid="101033" heatid="105337" lane="5" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.49" />
                    <SPLIT distance="100" swimtime="00:01:40.30" />
                    <SPLIT distance="150" swimtime="00:02:37.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="177" reactiontime="+118" swimtime="00:06:31.55" resultid="101034" heatid="106065" lane="4" entrytime="00:06:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.48" />
                    <SPLIT distance="100" swimtime="00:01:27.59" />
                    <SPLIT distance="150" swimtime="00:02:16.67" />
                    <SPLIT distance="200" swimtime="00:03:07.61" />
                    <SPLIT distance="250" swimtime="00:03:59.69" />
                    <SPLIT distance="300" swimtime="00:04:52.09" />
                    <SPLIT distance="350" swimtime="00:05:43.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-03-04" firstname="Wiktor" gender="M" lastname="DĘBSKI" nation="POL" swrid="4992887" athleteid="101035">
              <RESULTS>
                <RESULT eventid="98798" points="402" reactiontime="+97" swimtime="00:00:28.32" resultid="101036" heatid="105135" lane="0" entrytime="00:00:29.90" />
                <RESULT eventid="98924" points="347" reactiontime="+80" swimtime="00:00:34.20" resultid="101037" heatid="105186" lane="4" entrytime="00:00:35.50" />
                <RESULT eventid="99091" points="409" reactiontime="+108" swimtime="00:01:18.72" resultid="101038" heatid="105255" lane="5" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="460" reactiontime="+99" swimtime="00:00:34.53" resultid="101039" heatid="105359" lane="2" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-21" firstname="Maksym" gender="M" lastname="BABENKO" nation="POL" athleteid="101040">
              <RESULTS>
                <RESULT eventid="98956" status="DNS" swimtime="00:00:00.00" resultid="101041" heatid="105204" lane="6" entrytime="00:02:35.00" />
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="101042" heatid="105257" lane="5" entrytime="00:01:14.00" />
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="101043" heatid="105342" lane="9" entrytime="00:02:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-05-13" firstname="Michał" gender="M" lastname="WITKOWSKI" nation="POL" swrid="4180262" athleteid="101044">
              <RESULTS>
                <RESULT eventid="98798" points="449" reactiontime="+77" swimtime="00:00:27.29" resultid="101045" heatid="105140" lane="0" entrytime="00:00:27.07" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="101046" heatid="105224" lane="4" entrytime="00:01:01.15" />
                <RESULT eventid="99170" points="471" reactiontime="+70" swimtime="00:00:28.82" resultid="101047" heatid="105274" lane="6" entrytime="00:00:29.01" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-07-27" firstname="Bartosz" gender="M" lastname="BELDYGA" nation="POL" athleteid="101048">
              <RESULTS>
                <RESULT eventid="98798" points="371" reactiontime="+92" swimtime="00:00:29.10" resultid="101049" heatid="105136" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="98891" status="WDR" swimtime="00:00:00.00" resultid="101050" />
                <RESULT eventid="98988" points="407" swimtime="00:01:03.26" resultid="101051" heatid="105219" lane="7" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="352" reactiontime="+84" swimtime="00:00:31.74" resultid="101052" heatid="105273" lane="7" entrytime="00:00:30.00" />
                <RESULT eventid="99218" points="350" reactiontime="+84" swimtime="00:02:24.65" resultid="101053" heatid="105302" lane="7" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                    <SPLIT distance="100" swimtime="00:01:08.76" />
                    <SPLIT distance="150" swimtime="00:01:47.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="286" swimtime="00:01:15.59" resultid="101054" heatid="105328" lane="2" entrytime="00:01:20.00" />
                <RESULT eventid="99473" points="292" reactiontime="+89" swimtime="00:05:31.55" resultid="101055" heatid="106065" lane="9" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.38" />
                    <SPLIT distance="100" swimtime="00:01:14.39" />
                    <SPLIT distance="150" swimtime="00:01:56.91" />
                    <SPLIT distance="200" swimtime="00:02:40.64" />
                    <SPLIT distance="250" swimtime="00:03:24.64" />
                    <SPLIT distance="300" swimtime="00:04:09.03" />
                    <SPLIT distance="350" swimtime="00:04:53.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-05-05" firstname="Bogdan" gender="M" lastname="DUBIŃSKI" nation="POL" swrid="4992696" athleteid="101056">
              <RESULTS>
                <RESULT eventid="98798" points="241" reactiontime="+81" swimtime="00:00:33.56" resultid="101057" heatid="105130" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="98891" points="167" swimtime="00:26:19.97" resultid="101058" heatid="105423" lane="9" entrytime="00:26:30.00" />
                <RESULT eventid="98924" points="212" reactiontime="+81" swimtime="00:00:40.29" resultid="101059" heatid="105185" lane="1" entrytime="00:00:39.00" />
                <RESULT eventid="99020" points="97" reactiontime="+92" swimtime="00:04:01.94" resultid="101060" heatid="105233" lane="9" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.73" />
                    <SPLIT distance="100" swimtime="00:01:50.56" />
                    <SPLIT distance="150" swimtime="00:02:54.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="169" reactiontime="+91" swimtime="00:01:33.91" resultid="101061" heatid="105282" lane="2" entrytime="00:01:30.00" />
                <RESULT eventid="99282" points="146" reactiontime="+106" swimtime="00:07:42.67" resultid="101062" heatid="106048" lane="4" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.04" />
                    <SPLIT distance="100" swimtime="00:01:59.49" />
                    <SPLIT distance="150" swimtime="00:03:00.75" />
                    <SPLIT distance="200" swimtime="00:03:58.77" />
                    <SPLIT distance="250" swimtime="00:05:07.03" />
                    <SPLIT distance="300" swimtime="00:06:12.75" />
                    <SPLIT distance="350" swimtime="00:06:59.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="145" reactiontime="+101" swimtime="00:03:32.98" resultid="101063" heatid="105337" lane="3" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.24" />
                    <SPLIT distance="100" swimtime="00:01:46.64" />
                    <SPLIT distance="150" swimtime="00:02:41.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="196" reactiontime="+110" swimtime="00:06:18.59" resultid="101064" heatid="106064" lane="1" entrytime="00:06:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                    <SPLIT distance="100" swimtime="00:01:26.56" />
                    <SPLIT distance="150" swimtime="00:02:16.44" />
                    <SPLIT distance="200" swimtime="00:03:06.62" />
                    <SPLIT distance="250" swimtime="00:03:56.54" />
                    <SPLIT distance="300" swimtime="00:04:46.40" />
                    <SPLIT distance="350" swimtime="00:05:35.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-02-06" firstname="Bartosz" gender="M" lastname="PIERUCKI" nation="POL" athleteid="101065">
              <RESULTS>
                <RESULT eventid="98798" points="283" reactiontime="+81" swimtime="00:00:31.82" resultid="101066" heatid="105128" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="99170" points="246" reactiontime="+96" swimtime="00:00:35.76" resultid="101068" heatid="105268" lane="3" entrytime="00:00:36.00" />
                <RESULT eventid="99218" points="216" reactiontime="+93" swimtime="00:02:49.79" resultid="101069" heatid="105298" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.66" />
                    <SPLIT distance="100" swimtime="00:01:20.54" />
                    <SPLIT distance="150" swimtime="00:02:06.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="283" reactiontime="+86" swimtime="00:01:11.43" resultid="105390" heatid="105218" lane="8" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-03" firstname="Ilona" gender="F" lastname="SZKUDLARZ" nation="POL" athleteid="101070">
              <RESULTS>
                <RESULT eventid="98777" points="274" swimtime="00:00:36.52" resultid="101071" heatid="105116" lane="1" entrytime="00:00:36.40" />
                <RESULT eventid="98907" points="283" reactiontime="+78" swimtime="00:00:41.21" resultid="101072" heatid="105175" lane="3" entrytime="00:00:41.30" />
                <RESULT eventid="98972" points="264" reactiontime="+85" swimtime="00:01:21.07" resultid="101073" heatid="105208" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="265" reactiontime="+91" swimtime="00:01:40.10" resultid="101074" heatid="105245" lane="4" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="221" reactiontime="+96" swimtime="00:01:36.04" resultid="101075" heatid="105278" lane="2" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="258" reactiontime="+102" swimtime="00:02:57.37" resultid="101076" heatid="105290" lane="3" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.05" />
                    <SPLIT distance="100" swimtime="00:01:26.96" />
                    <SPLIT distance="150" swimtime="00:02:14.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="213" reactiontime="+87" swimtime="00:03:27.62" resultid="101077" heatid="105333" lane="0" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.48" />
                    <SPLIT distance="100" swimtime="00:01:39.43" />
                    <SPLIT distance="150" swimtime="00:02:33.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" status="WDR" swimtime="00:00:00.00" resultid="101078" entrytime="00:06:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-06-04" firstname="Karol" gender="M" lastname="SOSNA" nation="POL" athleteid="101245">
              <RESULTS>
                <RESULT eventid="98798" points="252" reactiontime="+112" swimtime="00:00:33.10" resultid="101249" heatid="105133" lane="0" entrytime="00:00:30.33" />
                <RESULT eventid="99091" points="319" reactiontime="+98" swimtime="00:01:25.53" resultid="101250" heatid="105251" lane="1" entrytime="00:01:39.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="308" reactiontime="+100" swimtime="00:01:09.42" resultid="101251" heatid="105217" lane="3" entrytime="00:01:12.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="394" reactiontime="+93" swimtime="00:00:36.37" resultid="101252" heatid="105356" lane="1" entrytime="00:00:40.15" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-12-08" firstname="Paweł" gender="M" lastname="STAWIARZ" nation="POL" athleteid="101246">
              <RESULTS>
                <RESULT eventid="98798" points="387" reactiontime="+77" swimtime="00:00:28.68" resultid="101253" heatid="105133" lane="8" entrytime="00:00:30.24" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-02-18" firstname="Robert" gender="M" lastname="NOWICKI" nation="POL" swrid="4754751" athleteid="101247">
              <RESULTS>
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="101254" heatid="105296" lane="0" entrytime="00:03:30.00" />
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="101255" entrytime="00:07:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-03-04" firstname="Norbert" gender="M" lastname="TCHORZEWSKI" nation="POL" athleteid="101248">
              <RESULTS>
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="101256" entrytime="00:05:50.00" />
                <RESULT eventid="99361" points="210" reactiontime="+85" swimtime="00:01:23.76" resultid="101257" heatid="105327" lane="0" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="179" reactiontime="+110" swimtime="00:07:12.33" resultid="101258" heatid="106050" lane="0" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.11" />
                    <SPLIT distance="100" swimtime="00:01:28.01" />
                    <SPLIT distance="150" swimtime="00:02:24.92" />
                    <SPLIT distance="200" swimtime="00:03:24.01" />
                    <SPLIT distance="250" swimtime="00:04:31.22" />
                    <SPLIT distance="300" swimtime="00:05:37.35" />
                    <SPLIT distance="350" swimtime="00:06:25.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="297" reactiontime="+79" swimtime="00:01:10.30" resultid="101259" heatid="105219" lane="9" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="101260" heatid="105132" lane="0" entrytime="00:00:31.00" />
                <RESULT eventid="98830" points="199" reactiontime="+95" swimtime="00:03:15.14" resultid="101261" heatid="105153" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                    <SPLIT distance="100" swimtime="00:01:24.05" />
                    <SPLIT distance="150" swimtime="00:02:28.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="289" reactiontime="+87" swimtime="00:00:33.90" resultid="104382" heatid="105270" lane="2" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-11-02" firstname="Monika" gender="F" lastname="NOWAK" nation="POL" swrid="4311814" athleteid="102587">
              <RESULTS>
                <RESULT eventid="98777" status="DNS" swimtime="00:00:00.00" resultid="102954" heatid="105119" lane="3" entrytime="00:00:31.49" entrycourse="LCM" />
                <RESULT eventid="98814" status="DNS" swimtime="00:00:00.00" resultid="102955" heatid="105145" lane="4" entrytime="00:03:10.00" />
                <RESULT eventid="98907" status="DNS" swimtime="00:00:00.00" resultid="102956" heatid="105176" lane="9" entrytime="00:00:40.00" />
                <RESULT eventid="98972" status="DNS" swimtime="00:00:00.00" resultid="102957" heatid="105211" lane="1" entrytime="00:01:10.00" />
                <RESULT eventid="99314" status="DNS" swimtime="00:00:00.00" resultid="102958" heatid="105279" lane="9" entrytime="00:01:30.00" />
                <RESULT eventid="99266" status="DNS" swimtime="00:00:00.00" resultid="102959" heatid="106046" lane="7" entrytime="00:07:00.00" />
                <RESULT eventid="99377" status="DNS" swimtime="00:00:00.00" resultid="102960" heatid="105333" lane="6" entrytime="00:03:10.00" />
                <RESULT eventid="99409" status="DNS" swimtime="00:00:00.00" resultid="102961" heatid="105347" lane="5" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-03-04" firstname="Piotr" gender="M" lastname="DROGOSZ" nation="POL" athleteid="102912">
              <RESULTS>
                <RESULT comment="04" eventid="98798" reactiontime="+80" status="DSQ" swimtime="00:00:28.36" resultid="102913" heatid="105123" lane="6" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="102914" heatid="105213" lane="0" />
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="102915" heatid="105248" lane="3" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="102916" heatid="105351" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-11-29" firstname="Andrzej" gender="M" lastname="DASZYŃSKI" nation="POL" swrid="4361205" athleteid="102917">
              <RESULTS>
                <RESULT eventid="98798" points="137" reactiontime="+86" swimtime="00:00:40.47" resultid="102946" heatid="105124" lane="7" entrytime="00:00:44.00" />
                <RESULT eventid="98830" points="92" reactiontime="+84" swimtime="00:04:11.74" resultid="102947" heatid="105149" lane="6" entrytime="00:04:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.99" />
                    <SPLIT distance="100" swimtime="00:02:03.41" />
                    <SPLIT distance="150" swimtime="00:03:18.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="107" reactiontime="+92" swimtime="00:00:50.52" resultid="102948" heatid="105181" lane="1" entrytime="00:00:55.00" />
                <RESULT eventid="99020" points="65" reactiontime="+84" swimtime="00:04:36.99" resultid="102949" heatid="105232" lane="8" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.00" />
                    <SPLIT distance="100" swimtime="00:02:13.22" />
                    <SPLIT distance="150" swimtime="00:03:28.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="100" reactiontime="+100" swimtime="00:01:51.86" resultid="102950" heatid="105282" lane="0" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="100" reactiontime="+96" swimtime="00:08:44.77" resultid="102951" heatid="106048" lane="2" entrytime="00:08:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.84" />
                    <SPLIT distance="100" swimtime="00:02:07.97" />
                    <SPLIT distance="150" swimtime="00:03:16.57" />
                    <SPLIT distance="200" swimtime="00:04:21.33" />
                    <SPLIT distance="250" swimtime="00:05:35.72" />
                    <SPLIT distance="300" swimtime="00:06:49.65" />
                    <SPLIT distance="350" swimtime="00:07:49.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="62" reactiontime="+89" swimtime="00:02:05.42" resultid="102952" heatid="105325" lane="7" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="103" reactiontime="+87" swimtime="00:03:58.21" resultid="102953" heatid="105337" lane="7" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.22" />
                    <SPLIT distance="100" swimtime="00:01:56.89" />
                    <SPLIT distance="150" swimtime="00:02:59.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-04-26" firstname="Rafał" gender="M" lastname="NOWAK" nation="POL" swrid="4311815" athleteid="102918">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="102962" heatid="105130" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="102963" heatid="105151" lane="4" entrytime="00:03:10.00" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="102964" heatid="105219" lane="1" entrytime="00:01:10.00" />
                <RESULT eventid="99020" status="DNS" swimtime="00:00:00.00" resultid="102965" heatid="105234" lane="1" entrytime="00:03:20.00" />
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="102966" heatid="105327" lane="9" entrytime="00:01:30.00" />
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="102967" entrytime="00:06:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-12" firstname="Zbigniew" gender="M" lastname="SZOZDA" nation="POL" athleteid="102919">
              <RESULTS>
                <RESULT eventid="98830" points="233" reactiontime="+115" swimtime="00:03:05.24" resultid="103015" heatid="105152" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.78" />
                    <SPLIT distance="100" swimtime="00:01:23.79" />
                    <SPLIT distance="150" swimtime="00:02:19.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="252" reactiontime="+77" swimtime="00:00:38.05" resultid="103016" heatid="105184" lane="7" entrytime="00:00:41.00" />
                <RESULT eventid="98956" points="233" reactiontime="+122" swimtime="00:03:26.37" resultid="103017" heatid="105199" lane="3" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.27" />
                    <SPLIT distance="100" swimtime="00:01:39.02" />
                    <SPLIT distance="150" swimtime="00:02:33.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="227" reactiontime="+129" swimtime="00:02:47.12" resultid="103018" heatid="105298" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.49" />
                    <SPLIT distance="100" swimtime="00:01:20.01" />
                    <SPLIT distance="150" swimtime="00:02:03.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" status="DNS" swimtime="00:00:00.00" resultid="103019" heatid="106049" lane="1" entrytime="00:07:40.00" />
                <RESULT comment="04" eventid="99425" reactiontime="+81" status="DSQ" swimtime="00:00:00.00" resultid="103020" heatid="105354" lane="7" entrytime="00:00:43.00" />
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="103021" entrytime="00:06:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-04-08" firstname="Łukasz" gender="M" lastname="RYBOŁOWICZ" nation="POL" athleteid="102920">
              <RESULTS>
                <RESULT eventid="98798" points="484" reactiontime="+62" swimtime="00:00:26.63" resultid="102987" heatid="105140" lane="9" entrytime="00:00:27.20" />
                <RESULT eventid="98830" points="318" reactiontime="+66" swimtime="00:02:46.91" resultid="102988" heatid="105154" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.92" />
                    <SPLIT distance="100" swimtime="00:01:22.23" />
                    <SPLIT distance="150" swimtime="00:02:10.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="481" reactiontime="+56" swimtime="00:00:59.85" resultid="102989" heatid="105226" lane="8" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99020" points="198" reactiontime="+82" swimtime="00:03:11.09" resultid="102990" heatid="105235" lane="1" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.98" />
                    <SPLIT distance="100" swimtime="00:01:28.85" />
                    <SPLIT distance="150" swimtime="00:02:19.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="102991" heatid="105254" lane="5" entrytime="00:01:23.00" />
                <RESULT eventid="99218" points="292" reactiontime="+68" swimtime="00:02:33.60" resultid="102992" heatid="105301" lane="7" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.09" />
                    <SPLIT distance="100" swimtime="00:01:15.47" />
                    <SPLIT distance="150" swimtime="00:01:55.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="298" reactiontime="+72" swimtime="00:01:14.53" resultid="102993" heatid="105328" lane="4" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="382" reactiontime="+69" swimtime="00:00:36.75" resultid="102994" heatid="105358" lane="7" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-01" firstname="Grzegorz" gender="M" lastname="MONCZAK" nation="POL" athleteid="102921">
              <RESULTS>
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="102980" heatid="105154" lane="4" entrytime="00:02:45.00" />
                <RESULT eventid="98891" status="WDR" swimtime="00:00:00.00" resultid="102982" entrytime="00:19:30.00" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="102983" heatid="105225" lane="4" entrytime="00:00:59.90" />
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="102984" heatid="105305" lane="9" entrytime="00:02:10.00" />
                <RESULT eventid="99282" status="DNS" swimtime="00:00:00.00" resultid="102985" heatid="106052" lane="2" entrytime="00:05:45.00" />
                <RESULT eventid="99473" status="WDR" swimtime="00:00:00.00" resultid="102986" entrytime="00:04:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-11-29" firstname="Edward" gender="M" lastname="DZIEKOŃSKI" nation="POL" athleteid="102922">
              <RESULTS>
                <RESULT eventid="99473" points="118" reactiontime="+125" swimtime="00:07:27.63" resultid="102972" heatid="106066" lane="2" entrytime="00:07:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.13" />
                    <SPLIT distance="100" swimtime="00:01:42.47" />
                    <SPLIT distance="150" swimtime="00:02:39.19" />
                    <SPLIT distance="200" swimtime="00:03:38.14" />
                    <SPLIT distance="250" swimtime="00:04:36.79" />
                    <SPLIT distance="300" swimtime="00:05:35.62" />
                    <SPLIT distance="350" swimtime="00:06:33.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="104" reactiontime="+105" swimtime="00:00:51.06" resultid="102973" heatid="105182" lane="0" entrytime="00:00:50.00" />
                <RESULT eventid="98798" points="150" reactiontime="+106" swimtime="00:00:39.33" resultid="102974" heatid="105125" lane="6" entrytime="00:00:39.00" />
                <RESULT eventid="98891" points="123" swimtime="00:29:08.92" resultid="102975" heatid="105424" lane="9" entrytime="00:29:50.00" />
                <RESULT eventid="98988" points="123" reactiontime="+112" swimtime="00:01:34.30" resultid="102976" heatid="105214" lane="0" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.21" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="04" eventid="99170" status="DSQ" swimtime="00:00:00.00" resultid="102977" heatid="105266" lane="7" entrytime="00:00:42.50" />
                <RESULT eventid="99218" points="113" reactiontime="+100" swimtime="00:03:30.71" resultid="102978" heatid="105296" lane="8" entrytime="00:03:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.52" />
                    <SPLIT distance="100" swimtime="00:01:43.15" />
                    <SPLIT distance="150" swimtime="00:02:38.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="76" reactiontime="+98" swimtime="00:04:23.29" resultid="102979" heatid="105337" lane="9" entrytime="00:04:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.72" />
                    <SPLIT distance="100" swimtime="00:02:08.89" />
                    <SPLIT distance="150" swimtime="00:03:17.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-06-28" firstname="Bolesław" gender="M" lastname="CZYŻ" nation="POL" swrid="4992699" athleteid="102923">
              <RESULTS>
                <RESULT eventid="99020" status="WDR" swimtime="00:00:00.00" resultid="102969" heatid="105232" lane="4" entrytime="00:04:10.00" />
                <RESULT eventid="99218" status="WDR" swimtime="00:00:00.00" resultid="102970" heatid="105295" lane="4" entrytime="00:03:35.00" />
                <RESULT eventid="99282" status="WDR" swimtime="00:00:00.00" resultid="102971" entrytime="00:08:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-02-06" firstname="Piotr" gender="M" lastname="DĄMBSKI" nation="POL" athleteid="102924">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="103007" heatid="105128" lane="3" entrytime="00:00:34.00" />
                <RESULT eventid="98830" status="DNS" swimtime="00:00:00.00" resultid="103008" heatid="105148" lane="8" />
                <RESULT eventid="98956" status="DNS" swimtime="00:00:00.00" resultid="103009" heatid="105196" lane="1" />
                <RESULT eventid="99020" status="DNS" swimtime="00:00:00.00" resultid="103010" heatid="105231" lane="5" />
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="103011" heatid="105249" lane="8" />
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="103012" heatid="105265" lane="8" />
                <RESULT eventid="99361" status="DNS" swimtime="00:00:00.00" resultid="103013" heatid="105324" lane="3" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="103014" heatid="105350" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-07-01" firstname="Katarzyna" gender="F" lastname="KOBA" nation="POL" swrid="4992695" athleteid="102925">
              <RESULTS>
                <RESULT eventid="98777" points="388" reactiontime="+85" swimtime="00:00:32.51" resultid="103004" heatid="105119" lane="8" entrytime="00:00:31.87" entrycourse="SCM" />
                <RESULT eventid="98972" points="333" swimtime="00:01:15.10" resultid="103005" heatid="105209" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="261" reactiontime="+85" swimtime="00:02:56.78" resultid="103006" heatid="105293" lane="9" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.61" />
                    <SPLIT distance="100" swimtime="00:01:22.50" />
                    <SPLIT distance="150" swimtime="00:02:10.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-17" firstname="Bogusław" gender="M" lastname="WOŹNIAK" nation="POL" athleteid="102926">
              <RESULTS>
                <RESULT eventid="98891" status="WDR" swimtime="00:00:00.00" resultid="102995" entrytime="00:22:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-05-15" firstname="Magdalena" gender="F" lastname="CZAPLA" nation="POL" swrid="4072135" athleteid="102929">
              <RESULTS>
                <RESULT eventid="98777" status="DNS" swimtime="00:00:00.00" resultid="103057" heatid="105120" lane="5" entrytime="00:00:29.82" entrycourse="LCM" />
                <RESULT eventid="98814" status="DNS" swimtime="00:00:00.00" resultid="103058" heatid="105147" lane="2" entrytime="00:02:50.00" />
                <RESULT eventid="98907" points="431" reactiontime="+83" swimtime="00:00:35.81" resultid="103059" heatid="105178" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="98940" points="409" reactiontime="+77" swimtime="00:03:07.33" resultid="103060" heatid="105194" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.49" />
                    <SPLIT distance="100" swimtime="00:01:30.44" />
                    <SPLIT distance="150" swimtime="00:02:20.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="338" reactiontime="+78" swimtime="00:01:32.31" resultid="103061" heatid="105247" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" status="DNS" swimtime="00:00:00.00" resultid="103062" heatid="105264" lane="9" entrytime="00:00:33.00" />
                <RESULT eventid="99344" status="DNS" swimtime="00:00:00.00" resultid="103063" heatid="105323" lane="6" entrytime="00:01:15.00" />
                <RESULT eventid="99409" status="DNS" swimtime="00:00:00.00" resultid="103064" heatid="105349" lane="5" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Anna" gender="F" lastname="KOTUSIŃSKA" nation="POL" swrid="4992692" athleteid="102930">
              <RESULTS>
                <RESULT comment="04" eventid="98972" reactiontime="+83" status="DSQ" swimtime="00:00:00.00" resultid="103055" heatid="105208" lane="6" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="207" reactiontime="+112" swimtime="00:00:42.32" resultid="103056" heatid="105261" lane="0" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-27" firstname="Magdalena" gender="F" lastname="KUMIŃSKA" nation="POL" athleteid="102932">
              <RESULTS>
                <RESULT eventid="98777" points="302" reactiontime="+69" swimtime="00:00:35.36" resultid="103026" heatid="105120" lane="8" entrytime="00:00:30.35" />
                <RESULT eventid="98907" points="213" reactiontime="+71" swimtime="00:00:45.26" resultid="103027" heatid="105178" lane="6" entrytime="00:00:33.45" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-09-16" firstname="Monika" gender="F" lastname="WINOGRODZKA" nation="POL" athleteid="102942">
              <RESULTS>
                <RESULT eventid="99314" points="352" reactiontime="+73" swimtime="00:01:22.27" resultid="102943" heatid="105280" lane="4" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="399" reactiontime="+70" swimtime="00:00:36.73" resultid="102944" heatid="105178" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="99409" points="313" reactiontime="+87" swimtime="00:00:43.39" resultid="102945" heatid="105349" lane="4" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-02-20" firstname="Zofia" gender="F" lastname="BRUNKA" nation="POL" athleteid="104376">
              <RESULTS>
                <RESULT eventid="98907" points="306" reactiontime="+70" swimtime="00:00:40.15" resultid="104377" heatid="105176" lane="6" entrytime="00:00:39.00" />
                <RESULT eventid="98972" points="358" reactiontime="+85" swimtime="00:01:13.30" resultid="104378" heatid="105210" lane="4" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="290" swimtime="00:00:37.85" resultid="104379" heatid="105262" lane="7" entrytime="00:00:36.00" />
                <RESULT eventid="99314" status="DNS" swimtime="00:00:00.00" resultid="104380" heatid="105280" lane="1" entrytime="00:01:21.00" />
                <RESULT eventid="99377" points="278" reactiontime="+74" swimtime="00:03:09.86" resultid="104381" heatid="105333" lane="2" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.71" />
                    <SPLIT distance="100" swimtime="00:01:31.70" />
                    <SPLIT distance="150" swimtime="00:02:21.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-02-01" firstname="Mariusz" gender="M" lastname="WÓJCICKI" nation="POL" athleteid="104398">
              <RESULTS>
                <RESULT eventid="98830" points="252" reactiontime="+85" swimtime="00:03:00.46" resultid="104399" heatid="105153" lane="4" entrytime="00:02:54.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                    <SPLIT distance="100" swimtime="00:01:17.05" />
                    <SPLIT distance="150" swimtime="00:02:15.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" points="302" reactiontime="+83" swimtime="00:00:35.80" resultid="104400" heatid="105187" lane="3" entrytime="00:00:33.72" />
                <RESULT eventid="99020" points="187" reactiontime="+90" swimtime="00:03:14.96" resultid="104401" heatid="105231" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.10" />
                    <SPLIT distance="100" swimtime="00:01:27.40" />
                    <SPLIT distance="150" swimtime="00:02:21.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="306" reactiontime="+86" swimtime="00:00:33.26" resultid="104402" heatid="105271" lane="2" entrytime="00:00:31.80" />
                <RESULT eventid="99186" points="272" reactiontime="+73" swimtime="00:01:20.12" resultid="104403" heatid="105285" lane="2" entrytime="00:01:17.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="289" reactiontime="+79" swimtime="00:01:15.31" resultid="104404" heatid="105324" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" points="216" reactiontime="+81" swimtime="00:03:06.42" resultid="104405" heatid="105340" lane="0" entrytime="00:02:55.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                    <SPLIT distance="100" swimtime="00:01:26.65" />
                    <SPLIT distance="150" swimtime="00:02:16.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-14" firstname="Andrzej" gender="M" lastname="FAJDASZ" nation="POL" athleteid="105067">
              <RESULTS>
                <RESULT eventid="98798" points="362" reactiontime="+79" swimtime="00:00:29.33" resultid="105072" heatid="105133" lane="7" entrytime="00:00:30.15" />
                <RESULT eventid="98830" points="283" reactiontime="+81" swimtime="00:02:53.61" resultid="105073" heatid="105153" lane="7" entrytime="00:02:55.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                    <SPLIT distance="100" swimtime="00:01:21.46" />
                    <SPLIT distance="150" swimtime="00:02:13.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="263" reactiontime="+79" swimtime="00:00:34.99" resultid="105074" heatid="105270" lane="7" entrytime="00:00:34.30" />
                <RESULT eventid="99186" points="238" reactiontime="+84" swimtime="00:01:23.75" resultid="105075" heatid="105285" lane="7" entrytime="00:01:17.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.65" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="04" eventid="98988" reactiontime="+69" status="WDR" swimtime="00:00:00.00" resultid="105076" heatid="105223" lane="6" entrytime="00:01:03.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-05-20" firstname="Katarzyna" gender="F" lastname="MICHAŁOWSKA" nation="POL" athleteid="105068">
              <RESULTS>
                <RESULT eventid="98972" points="306" reactiontime="+113" swimtime="00:01:17.23" resultid="105069" heatid="105210" lane="2" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="272" reactiontime="+110" swimtime="00:02:54.26" resultid="105070" heatid="105292" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.30" />
                    <SPLIT distance="100" swimtime="00:01:20.95" />
                    <SPLIT distance="150" swimtime="00:02:07.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="263" reactiontime="+108" swimtime="00:06:13.12" resultid="105071" heatid="106055" lane="6" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.70" />
                    <SPLIT distance="100" swimtime="00:01:25.92" />
                    <SPLIT distance="150" swimtime="00:02:13.12" />
                    <SPLIT distance="200" swimtime="00:03:01.36" />
                    <SPLIT distance="250" swimtime="00:03:49.74" />
                    <SPLIT distance="300" swimtime="00:04:38.42" />
                    <SPLIT distance="350" swimtime="00:05:27.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="UKR" region="ZTM" clubid="100642" name="Zhytomyr Aqua Masters">
          <CONTACT city="ZHYTOMYR" email="reservation007@mail.ru" fax="+380412418911" internet="mastersswim.com.ua" name="IGOR KUKHARYEV" phone="+380674102880" state="UKR" street="MOSKOVSKA 35, APT 4" zip="10029" />
          <ATHLETES>
            <ATHLETE birthdate="1974-02-05" firstname="Volodymyr" gender="M" lastname="KRYUKOV" nation="UKR" swrid="4992747" athleteid="100654">
              <RESULTS>
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="100655" heatid="105256" lane="1" entrytime="00:01:20.06" entrycourse="LCM" />
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="100656" heatid="105273" lane="8" entrytime="00:00:30.03" entrycourse="LCM" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="100657" heatid="105360" lane="0" entrytime="00:00:35.02" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-11-02" firstname="Petro" gender="M" lastname="KHYMOVYCH" nation="UKR" swrid="4776780" athleteid="100658">
              <RESULTS>
                <RESULT eventid="98924" points="281" reactiontime="+87" swimtime="00:00:36.70" resultid="100659" heatid="105186" lane="8" entrytime="00:00:36.10" entrycourse="SCM" />
                <RESULT eventid="99186" points="263" reactiontime="+75" swimtime="00:01:20.99" resultid="100660" heatid="105285" lane="6" entrytime="00:01:17.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="100661" heatid="105340" lane="3" entrytime="00:02:50.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-06-06" firstname="Mykhaylo" gender="M" lastname="YURCHAK" nation="UKR" athleteid="100662">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="100663" heatid="105140" lane="8" entrytime="00:00:27.02" entrycourse="SCM" />
                <RESULT eventid="98988" points="347" reactiontime="+89" swimtime="00:01:06.74" resultid="100664" heatid="105225" lane="6" entrytime="00:01:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-12-09" firstname="Oleksiy" gender="M" lastname="YRCHAK" nation="UKR" athleteid="100665">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="100666" heatid="105134" lane="2" entrytime="00:00:30.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="RUS" clubid="103075" name="Zvezdy Rosii">
          <CONTACT email="a.tervinsky@gov39.ru" name="Trevinski Aleksandr" />
          <ATHLETES>
            <ATHLETE birthdate="1938-01-01" firstname="Luiza" gender="F" lastname="SHCHERBICH" nation="RUS" swrid="4382600" athleteid="103076">
              <RESULTS>
                <RESULT eventid="98777" points="47" reactiontime="+128" swimtime="00:01:05.38" resultid="103077" heatid="105113" lane="8" entrytime="00:00:58.16" entrycourse="SCM" />
                <RESULT eventid="98972" points="34" reactiontime="+125" swimtime="00:02:39.90" resultid="103078" heatid="105205" lane="4" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="60" reactiontime="+116" swimtime="00:02:43.78" resultid="103079" heatid="105243" lane="4" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="61" reactiontime="+113" swimtime="00:01:14.50" resultid="103080" heatid="105344" lane="8" entrytime="00:01:09.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Elena" gender="F" lastname="KOLYADINA" nation="RUS" swrid="4776662" athleteid="103081">
              <RESULTS>
                <RESULT eventid="98777" points="260" reactiontime="+95" swimtime="00:00:37.16" resultid="103082" heatid="105116" lane="4" entrytime="00:00:35.60" />
                <RESULT eventid="98940" points="264" reactiontime="+104" swimtime="00:03:36.61" resultid="103083" heatid="105193" lane="1" entrytime="00:03:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.72" />
                    <SPLIT distance="100" swimtime="00:01:45.57" />
                    <SPLIT distance="150" swimtime="00:02:40.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" points="269" reactiontime="+95" swimtime="00:01:39.61" resultid="103084" heatid="105246" lane="1" entrytime="00:01:38.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="285" reactiontime="+89" swimtime="00:00:44.78" resultid="103085" heatid="105347" lane="6" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Natalia" gender="F" lastname="ALESHCHENKO" nation="RUS" swrid="4269968" athleteid="103086">
              <RESULTS>
                <RESULT eventid="98777" points="335" reactiontime="+85" swimtime="00:00:34.16" resultid="103087" heatid="105117" lane="9" entrytime="00:00:35.20" />
                <RESULT eventid="98814" points="300" reactiontime="+84" swimtime="00:03:08.40" resultid="103088" heatid="105146" lane="9" entrytime="00:03:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.44" />
                    <SPLIT distance="100" swimtime="00:01:28.49" />
                    <SPLIT distance="150" swimtime="00:02:23.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="319" reactiontime="+98" swimtime="00:01:16.17" resultid="103089" heatid="105208" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="301" reactiontime="+103" swimtime="00:00:37.39" resultid="103090" heatid="105261" lane="3" entrytime="00:00:38.50" />
                <RESULT eventid="99409" points="257" reactiontime="+95" swimtime="00:00:46.31" resultid="103091" heatid="105347" lane="7" entrytime="00:00:44.50" />
                <RESULT eventid="99457" points="279" reactiontime="+91" swimtime="00:06:05.73" resultid="103092" heatid="106055" lane="9" entrytime="00:05:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.95" />
                    <SPLIT distance="100" swimtime="00:01:27.12" />
                    <SPLIT distance="150" swimtime="00:02:14.58" />
                    <SPLIT distance="200" swimtime="00:03:02.52" />
                    <SPLIT distance="250" swimtime="00:03:50.17" />
                    <SPLIT distance="300" swimtime="00:04:37.72" />
                    <SPLIT distance="350" swimtime="00:05:24.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-01-01" firstname="Irina" gender="F" lastname="TITOVA" nation="RUS" athleteid="103093">
              <RESULTS>
                <RESULT eventid="98777" points="287" reactiontime="+89" swimtime="00:00:35.95" resultid="103094" heatid="105116" lane="8" entrytime="00:00:36.50" />
                <RESULT eventid="98972" points="302" reactiontime="+113" swimtime="00:01:17.60" resultid="103095" heatid="105208" lane="2" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99202" points="306" swimtime="00:02:47.50" resultid="103096" heatid="105292" lane="8" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                    <SPLIT distance="100" swimtime="00:01:19.64" />
                    <SPLIT distance="150" swimtime="00:02:03.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" status="WDR" swimtime="00:00:00.00" resultid="103097" entrytime="00:06:03.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-01" firstname="Marina" gender="F" lastname="KILINA" nation="RUS" swrid="4302393" athleteid="103098">
              <RESULTS>
                <RESULT eventid="98777" points="341" reactiontime="+90" swimtime="00:00:33.95" resultid="103099" heatid="105118" lane="9" entrytime="00:00:34.01" entrycourse="LCM" />
                <RESULT eventid="98907" points="323" reactiontime="+79" swimtime="00:00:39.40" resultid="103100" heatid="105176" lane="8" entrytime="00:00:39.50" />
                <RESULT eventid="99154" status="DNS" swimtime="00:00:00.00" resultid="103101" heatid="105261" lane="4" entrytime="00:00:37.50" />
                <RESULT eventid="99314" status="DNS" swimtime="00:00:00.00" resultid="103102" heatid="105279" lane="8" entrytime="00:01:27.50" />
                <RESULT eventid="99409" status="DNS" swimtime="00:00:00.00" resultid="103103" heatid="105347" lane="3" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-01" firstname="Olga" gender="F" lastname="TIKHOMIROVA" nation="RUS" swrid="4792314" athleteid="103104">
              <RESULTS>
                <RESULT eventid="98814" status="DNS" swimtime="00:00:00.00" resultid="103105" heatid="105145" lane="9" entrytime="00:03:39.00" />
                <RESULT eventid="98907" status="DNS" swimtime="00:00:00.00" resultid="103106" heatid="105174" lane="6" entrytime="00:00:44.50" />
                <RESULT eventid="99154" status="DNS" swimtime="00:00:00.00" resultid="103107" heatid="105260" lane="8" entrytime="00:00:44.00" />
                <RESULT eventid="99314" status="DNS" swimtime="00:00:00.00" resultid="103108" heatid="105278" lane="0" entrytime="00:01:43.50" />
                <RESULT eventid="99344" status="DNS" swimtime="00:00:00.00" resultid="103109" heatid="105322" lane="8" entrytime="00:01:42.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-01-01" firstname="Tatiana" gender="F" lastname="LOGVINOVA" nation="RUS" swrid="4992865" athleteid="103110">
              <RESULTS>
                <RESULT eventid="98777" points="216" reactiontime="+88" swimtime="00:00:39.53" resultid="103111" heatid="105116" lane="9" entrytime="00:00:36.53" entrycourse="SCM" />
                <RESULT eventid="98814" points="221" reactiontime="+100" swimtime="00:03:28.37" resultid="103112" heatid="105144" lane="4" entrytime="00:03:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.76" />
                    <SPLIT distance="100" swimtime="00:01:43.03" />
                    <SPLIT distance="150" swimtime="00:02:41.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98907" points="198" reactiontime="+77" swimtime="00:00:46.42" resultid="103113" heatid="105174" lane="3" entrytime="00:00:44.50" />
                <RESULT eventid="98940" points="229" reactiontime="+116" swimtime="00:03:47.20" resultid="103114" heatid="105192" lane="5" entrytime="00:03:46.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.58" />
                    <SPLIT distance="100" swimtime="00:01:51.24" />
                    <SPLIT distance="150" swimtime="00:02:50.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99089" status="DNS" swimtime="00:00:00.00" resultid="103115" heatid="105246" lane="9" entrytime="00:01:41.50" />
                <RESULT eventid="99314" points="182" reactiontime="+82" swimtime="00:01:42.50" resultid="103116" heatid="105278" lane="1" entrytime="00:01:41.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99409" points="255" reactiontime="+91" swimtime="00:00:46.43" resultid="103117" heatid="105347" lane="1" entrytime="00:00:44.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-01" firstname="Olga" gender="F" lastname="BORISOVA" nation="RUS" swrid="4595550" athleteid="103118">
              <RESULTS>
                <RESULT eventid="98777" points="586" reactiontime="+81" swimtime="00:00:28.35" resultid="103119" heatid="105121" lane="5" entrytime="00:00:27.97" entrycourse="LCM" />
                <RESULT eventid="98972" points="560" reactiontime="+69" swimtime="00:01:03.17" resultid="103120" heatid="105212" lane="9" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="471" reactiontime="+83" swimtime="00:00:32.20" resultid="103121" heatid="105263" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="99202" points="490" reactiontime="+67" swimtime="00:02:23.22" resultid="103122" heatid="105294" lane="8" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                    <SPLIT distance="100" swimtime="00:01:12.10" />
                    <SPLIT distance="150" swimtime="00:01:48.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-01" firstname="Elena" gender="F" lastname="DAUTOVA" nation="RUS" swrid="4754732" athleteid="103123">
              <RESULTS>
                <RESULT eventid="98777" points="373" reactiontime="+82" swimtime="00:00:32.96" resultid="103124" heatid="105119" lane="9" entrytime="00:00:32.13" entrycourse="SCM" />
                <RESULT eventid="98907" points="333" reactiontime="+79" swimtime="00:00:39.04" resultid="103125" heatid="105176" lane="2" entrytime="00:00:39.00" />
                <RESULT eventid="98972" points="348" reactiontime="+82" swimtime="00:01:13.96" resultid="103126" heatid="105210" lane="9" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="268" reactiontime="+67" swimtime="00:01:30.08" resultid="103127" heatid="105279" lane="4" entrytime="00:01:24.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99377" points="235" reactiontime="+60" swimtime="00:03:21.00" resultid="103128" heatid="105333" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.22" />
                    <SPLIT distance="100" swimtime="00:01:37.89" />
                    <SPLIT distance="150" swimtime="00:02:31.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-01" firstname="Olga" gender="F" lastname="VERYUKINA" nation="RUS" swrid="4754733" athleteid="103129">
              <RESULTS>
                <RESULT eventid="98777" points="389" reactiontime="+89" swimtime="00:00:32.49" resultid="103130" heatid="105119" lane="6" entrytime="00:00:31.50" entrycourse="SCM" />
                <RESULT eventid="98814" points="345" reactiontime="+88" swimtime="00:02:59.76" resultid="103131" heatid="105146" lane="6" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.05" />
                    <SPLIT distance="100" swimtime="00:01:25.93" />
                    <SPLIT distance="150" swimtime="00:02:17.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98972" points="370" reactiontime="+99" swimtime="00:01:12.48" resultid="103132" heatid="105211" lane="0" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="357" reactiontime="+98" swimtime="00:00:35.31" resultid="103133" heatid="105263" lane="0" entrytime="00:00:34.50" />
                <RESULT eventid="99202" points="362" reactiontime="+93" swimtime="00:02:38.49" resultid="103134" heatid="105293" lane="7" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                    <SPLIT distance="100" swimtime="00:01:16.70" />
                    <SPLIT distance="150" swimtime="00:01:57.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" points="365" reactiontime="+95" swimtime="00:05:34.37" resultid="103135" heatid="106055" lane="4" entrytime="00:05:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.27" />
                    <SPLIT distance="100" swimtime="00:01:19.73" />
                    <SPLIT distance="150" swimtime="00:02:01.71" />
                    <SPLIT distance="200" swimtime="00:02:44.84" />
                    <SPLIT distance="250" swimtime="00:03:27.76" />
                    <SPLIT distance="300" swimtime="00:04:11.24" />
                    <SPLIT distance="350" swimtime="00:04:53.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-01" firstname="Alla" gender="F" lastname="FEOKTISTOVA" nation="RUS" swrid="4875570" athleteid="103136">
              <RESULTS>
                <RESULT eventid="98777" points="501" reactiontime="+97" swimtime="00:00:29.86" resultid="103137" heatid="105121" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="98814" points="453" reactiontime="+103" swimtime="00:02:44.18" resultid="103138" heatid="105147" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="100" swimtime="00:01:19.43" />
                    <SPLIT distance="150" swimtime="00:02:06.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="547" reactiontime="+98" swimtime="00:00:30.64" resultid="103139" heatid="105264" lane="3" entrytime="00:00:30.50" />
                <RESULT eventid="99344" points="495" reactiontime="+87" swimtime="00:01:10.73" resultid="103140" heatid="105323" lane="5" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-01-01" firstname="Regina" gender="F" lastname="SYCH" nation="RUS" swrid="4042762" athleteid="103141">
              <RESULTS>
                <RESULT eventid="98777" points="633" reactiontime="+92" swimtime="00:00:27.63" resultid="103142" heatid="105121" lane="3" entrytime="00:00:28.56" entrycourse="LCM" />
                <RESULT eventid="98972" points="625" reactiontime="+95" swimtime="00:01:00.88" resultid="103143" heatid="105212" lane="1" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99154" points="553" reactiontime="+84" swimtime="00:00:30.53" resultid="103144" heatid="105264" lane="6" entrytime="00:00:30.50" />
                <RESULT eventid="99202" points="598" reactiontime="+84" swimtime="00:02:14.06" resultid="103145" heatid="105294" lane="6" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.88" />
                    <SPLIT distance="100" swimtime="00:01:05.14" />
                    <SPLIT distance="150" swimtime="00:01:39.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99457" status="WDR" swimtime="00:00:00.00" resultid="103146" entrytime="00:05:04.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-01-01" firstname="Vyacheslav" gender="M" lastname="TIKHONOV" nation="RUS" athleteid="103147">
              <RESULTS>
                <RESULT eventid="98798" points="213" reactiontime="+95" swimtime="00:00:35.00" resultid="103148" heatid="105127" lane="8" entrytime="00:00:35.80" />
                <RESULT eventid="98924" points="147" reactiontime="+117" swimtime="00:00:45.45" resultid="103149" heatid="105183" lane="0" entrytime="00:00:45.00" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="103150" heatid="105215" lane="2" entrytime="00:01:22.50" />
                <RESULT eventid="99170" points="122" reactiontime="+119" swimtime="00:00:45.16" resultid="103151" heatid="105266" lane="1" entrytime="00:00:43.00" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="103152" heatid="105353" lane="8" entrytime="00:00:45.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-01-01" firstname="Boris" gender="M" lastname="KOZYNCHENKO" nation="RUS" athleteid="103153">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="103154" heatid="105125" lane="2" entrytime="00:00:39.00" />
                <RESULT comment="Rekord Litwy 800 dow" eventid="98891" status="DNS" swimtime="00:00:00.00" resultid="103155" heatid="105424" lane="7" entrytime="00:27:19.00">
                  <SPLITS>
                    <SPLIT distance="800" swimtime="00:15:51.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98924" status="DNS" swimtime="00:00:00.00" resultid="103156" heatid="105182" lane="8" entrytime="00:00:49.50" />
                <RESULT eventid="98956" status="DNS" swimtime="00:00:00.00" resultid="103157" heatid="105196" lane="5" entrytime="00:04:19.00" />
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="103158" heatid="105249" lane="6" entrytime="00:01:56.00" />
                <RESULT eventid="99218" status="DNS" swimtime="00:00:00.00" resultid="103159" heatid="105296" lane="6" entrytime="00:03:19.00" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="103160" heatid="105351" lane="4" entrytime="00:00:49.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-01" firstname="Vitaliy" gender="M" lastname="AVDEEV" nation="RUS" swrid="4754734" athleteid="103161">
              <RESULTS>
                <RESULT eventid="98798" points="205" reactiontime="+108" swimtime="00:00:35.42" resultid="103162" heatid="105126" lane="6" entrytime="00:00:36.20" />
                <RESULT eventid="98830" points="158" reactiontime="+110" swimtime="00:03:30.87" resultid="103163" heatid="105150" lane="2" entrytime="00:03:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.94" />
                    <SPLIT distance="100" swimtime="00:01:47.29" />
                    <SPLIT distance="150" swimtime="00:02:47.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="98988" points="218" reactiontime="+107" swimtime="00:01:17.94" resultid="103164" heatid="105215" lane="6" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="194" reactiontime="+118" swimtime="00:00:38.68" resultid="103165" heatid="105267" lane="2" entrytime="00:00:39.00" />
                <RESULT eventid="99218" points="192" reactiontime="+115" swimtime="00:02:56.80" resultid="103166" heatid="105297" lane="1" entrytime="00:03:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.99" />
                    <SPLIT distance="100" swimtime="00:01:25.32" />
                    <SPLIT distance="150" swimtime="00:02:11.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="182" reactiontime="+108" swimtime="00:00:47.05" resultid="103167" heatid="105352" lane="3" entrytime="00:00:47.50" />
                <RESULT eventid="99473" points="202" reactiontime="+120" swimtime="00:06:15.06" resultid="103168" heatid="106065" lane="3" entrytime="00:06:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.32" />
                    <SPLIT distance="100" swimtime="00:01:25.50" />
                    <SPLIT distance="150" swimtime="00:02:12.74" />
                    <SPLIT distance="200" swimtime="00:03:02.09" />
                    <SPLIT distance="250" swimtime="00:03:51.60" />
                    <SPLIT distance="300" swimtime="00:04:41.51" />
                    <SPLIT distance="350" swimtime="00:05:29.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-01" firstname="Yuriy" gender="M" lastname="YAKOVENKO" nation="RUS" swrid="4223539" athleteid="103169">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="103170" heatid="105129" lane="6" entrytime="00:00:32.90" />
                <RESULT eventid="98924" status="DNS" swimtime="00:00:00.00" resultid="103171" heatid="105182" lane="4" entrytime="00:00:46.50" />
                <RESULT eventid="98956" status="DNS" swimtime="00:00:00.00" resultid="103172" heatid="105197" lane="5" entrytime="00:03:54.00" />
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="103173" heatid="105250" lane="3" entrytime="00:01:46.00" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="103174" heatid="105354" lane="0" entrytime="00:00:43.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Akim" gender="M" lastname="DENISENKO" nation="RUS" swrid="4223536" athleteid="103175">
              <RESULTS>
                <RESULT eventid="98798" points="188" reactiontime="+100" swimtime="00:00:36.46" resultid="103176" heatid="105128" lane="1" entrytime="00:00:34.40" />
                <RESULT eventid="98988" points="140" swimtime="00:01:30.17" resultid="103177" heatid="105215" lane="7" entrytime="00:01:23.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="132" reactiontime="+107" swimtime="00:00:44.03" resultid="103178" heatid="105266" lane="2" entrytime="00:00:42.50" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="103179" heatid="105353" lane="9" entrytime="00:00:46.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Viktor" gender="M" lastname="POPOV" nation="RUS" athleteid="103180">
              <RESULTS>
                <RESULT eventid="98798" points="237" reactiontime="+102" swimtime="00:00:33.75" resultid="103181" heatid="105128" lane="4" entrytime="00:00:33.40" />
                <RESULT eventid="98924" points="170" reactiontime="+133" swimtime="00:00:43.32" resultid="103182" heatid="105183" lane="3" entrytime="00:00:42.80" />
                <RESULT eventid="98988" points="192" reactiontime="+107" swimtime="00:01:21.26" resultid="103183" heatid="105216" lane="0" entrytime="00:01:19.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99186" points="160" reactiontime="+81" swimtime="00:01:35.67" resultid="103184" heatid="105283" lane="9" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="103185" heatid="105353" lane="4" entrytime="00:00:44.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-02-01" firstname="Aleksandr" gender="M" lastname="TERVINSKI" nation="RUS" athleteid="103186">
              <RESULTS>
                <RESULT comment="04" eventid="98798" status="DSQ" swimtime="00:00:00.00" resultid="103187" heatid="105128" lane="7" entrytime="00:00:34.40" />
                <RESULT eventid="98924" points="190" reactiontime="+88" swimtime="00:00:41.77" resultid="103188" heatid="105183" lane="6" entrytime="00:00:42.90" />
                <RESULT eventid="98956" points="192" reactiontime="+101" swimtime="00:03:40.02" resultid="103189" heatid="105198" lane="6" entrytime="00:03:43.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.76" />
                    <SPLIT distance="100" swimtime="00:01:47.58" />
                    <SPLIT distance="150" swimtime="00:02:46.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="217" reactiontime="+89" swimtime="00:01:37.22" resultid="103190" heatid="105251" lane="9" entrytime="00:01:40.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="283" reactiontime="+94" swimtime="00:00:40.58" resultid="103191" heatid="105354" lane="5" entrytime="00:00:42.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-02-01" firstname="Sergey" gender="M" lastname="MIKHAYLOV" nation="RUS" athleteid="103192">
              <RESULTS>
                <RESULT eventid="98798" points="127" reactiontime="+106" swimtime="00:00:41.58" resultid="103193" heatid="105125" lane="7" entrytime="00:00:39.50" />
                <RESULT eventid="98891" points="147" swimtime="00:27:27.83" resultid="103194" heatid="105424" lane="3" entrytime="00:26:59.00" />
                <RESULT eventid="98988" points="135" reactiontime="+117" swimtime="00:01:31.42" resultid="103195" heatid="105215" lane="1" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="140" reactiontime="+99" swimtime="00:03:16.42" resultid="103196" heatid="105296" lane="4" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.02" />
                    <SPLIT distance="100" swimtime="00:01:34.40" />
                    <SPLIT distance="150" swimtime="00:02:26.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="156" reactiontime="+122" swimtime="00:06:48.65" resultid="103197" heatid="106065" lane="0" entrytime="00:06:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.29" />
                    <SPLIT distance="100" swimtime="00:01:37.00" />
                    <SPLIT distance="150" swimtime="00:02:30.29" />
                    <SPLIT distance="200" swimtime="00:03:23.85" />
                    <SPLIT distance="250" swimtime="00:04:16.82" />
                    <SPLIT distance="300" swimtime="00:05:08.79" />
                    <SPLIT distance="350" swimtime="00:06:00.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-02-01" firstname="Vladlen" gender="M" lastname="NESVETAEV" nation="RUS" swrid="4776740" athleteid="103198">
              <RESULTS>
                <RESULT eventid="99020" points="299" reactiontime="+88" swimtime="00:02:46.67" resultid="103199" heatid="105236" lane="8" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.87" />
                    <SPLIT distance="100" swimtime="00:01:17.82" />
                    <SPLIT distance="150" swimtime="00:02:02.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99282" points="367" reactiontime="+86" swimtime="00:05:40.39" resultid="103200" heatid="106053" lane="8" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                    <SPLIT distance="100" swimtime="00:01:13.70" />
                    <SPLIT distance="150" swimtime="00:02:00.59" />
                    <SPLIT distance="200" swimtime="00:02:45.66" />
                    <SPLIT distance="250" swimtime="00:03:36.35" />
                    <SPLIT distance="300" swimtime="00:04:25.63" />
                    <SPLIT distance="350" swimtime="00:05:04.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99361" points="363" reactiontime="+88" swimtime="00:01:09.83" resultid="103201" heatid="105330" lane="2" entrytime="00:01:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="409" reactiontime="+92" swimtime="00:04:56.34" resultid="103202" heatid="106060" lane="2" entrytime="00:04:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                    <SPLIT distance="100" swimtime="00:01:10.59" />
                    <SPLIT distance="150" swimtime="00:01:48.20" />
                    <SPLIT distance="200" swimtime="00:02:26.58" />
                    <SPLIT distance="250" swimtime="00:03:04.56" />
                    <SPLIT distance="300" swimtime="00:03:43.24" />
                    <SPLIT distance="350" swimtime="00:04:20.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-01" firstname="Grigoriy" gender="M" lastname="LOPIN" nation="RUS" swrid="4992861" athleteid="103203">
              <RESULTS>
                <RESULT eventid="98798" points="274" reactiontime="+107" swimtime="00:00:32.17" resultid="103204" heatid="105131" lane="0" entrytime="00:00:31.80" />
                <RESULT eventid="98891" points="161" swimtime="00:26:37.84" resultid="103205" heatid="105423" lane="5" entrytime="00:23:39.00" />
                <RESULT eventid="98956" points="219" reactiontime="+99" swimtime="00:03:30.45" resultid="103206" heatid="105200" lane="9" entrytime="00:03:26.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.40" />
                    <SPLIT distance="100" swimtime="00:01:38.29" />
                    <SPLIT distance="150" swimtime="00:02:32.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99091" points="243" reactiontime="+107" swimtime="00:01:33.62" resultid="103207" heatid="105252" lane="1" entrytime="00:01:31.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99425" points="287" reactiontime="+91" swimtime="00:00:40.39" resultid="103208" heatid="105356" lane="8" entrytime="00:00:40.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-01" firstname="Sergey" gender="M" lastname="DIRINDYAEV" nation="RUS" swrid="4992862" athleteid="103209">
              <RESULTS>
                <RESULT eventid="98798" points="333" reactiontime="+83" swimtime="00:00:30.14" resultid="103210" heatid="105132" lane="6" entrytime="00:00:30.80" />
                <RESULT eventid="98891" points="191" swimtime="00:25:11.87" resultid="103211" heatid="105423" lane="3" entrytime="00:23:39.00" />
                <RESULT eventid="98924" status="DNS" swimtime="00:00:00.00" resultid="103212" heatid="105184" lane="8" entrytime="00:00:41.80" />
                <RESULT eventid="98988" points="334" reactiontime="+85" swimtime="00:01:07.58" resultid="103213" heatid="105220" lane="9" entrytime="00:01:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="239" reactiontime="+77" swimtime="00:00:36.11" resultid="103214" heatid="105269" lane="8" entrytime="00:00:35.50" />
                <RESULT eventid="99425" points="275" reactiontime="+78" swimtime="00:00:40.97" resultid="103215" heatid="105355" lane="3" entrytime="00:00:41.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-01" firstname="Aleksandr" gender="M" lastname="SINILNIKOV" nation="RUS" athleteid="103216">
              <RESULTS>
                <RESULT eventid="98798" points="277" reactiontime="+95" swimtime="00:00:32.06" resultid="103217" heatid="105131" lane="1" entrytime="00:00:31.50" />
                <RESULT eventid="98924" points="131" reactiontime="+88" swimtime="00:00:47.22" resultid="103218" heatid="105184" lane="0" entrytime="00:00:41.80" />
                <RESULT eventid="98988" points="230" reactiontime="+110" swimtime="00:01:16.47" resultid="103219" heatid="105217" lane="2" entrytime="00:01:13.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="248" reactiontime="+103" swimtime="00:00:35.68" resultid="103220" heatid="105269" lane="0" entrytime="00:00:35.50" />
                <RESULT eventid="99425" points="204" reactiontime="+101" swimtime="00:00:45.30" resultid="103221" heatid="105355" lane="6" entrytime="00:00:41.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-01-01" firstname="Andrey" gender="M" lastname="MAKAROV" nation="RUS" athleteid="103222">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="103223" heatid="105132" lane="3" entrytime="00:00:30.80" />
                <RESULT eventid="98956" status="DNS" swimtime="00:00:00.00" resultid="103224" heatid="105201" lane="5" entrytime="00:03:09.00" />
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="103225" heatid="105255" lane="0" entrytime="00:01:22.50" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="103226" heatid="105359" lane="0" entrytime="00:00:36.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-01-01" firstname="Vadim" gender="M" lastname="EZHKOV" nation="RUS" swrid="4754735" athleteid="103227">
              <RESULTS>
                <RESULT eventid="98798" points="304" reactiontime="+78" swimtime="00:00:31.08" resultid="103228" heatid="105131" lane="2" entrytime="00:00:31.20" />
                <RESULT eventid="98956" status="DNS" swimtime="00:00:00.00" resultid="103229" heatid="105202" lane="7" entrytime="00:03:04.00" />
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="103230" heatid="105254" lane="4" entrytime="00:01:23.00" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="103231" heatid="105359" lane="8" entrytime="00:00:36.50" />
                <RESULT eventid="99170" points="279" reactiontime="+75" swimtime="00:00:34.32" resultid="105095" heatid="105270" lane="3" entrytime="00:00:33.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Viktor" gender="M" lastname="LYUBAVIN" nation="RUS" swrid="4754736" athleteid="103232">
              <RESULTS>
                <RESULT eventid="98798" points="380" reactiontime="+75" swimtime="00:00:28.85" resultid="103233" heatid="105138" lane="9" entrytime="00:00:28.40" />
                <RESULT eventid="98891" status="DNF" swimtime="00:00:00.00" resultid="103234" heatid="105421" lane="7" entrytime="00:21:09.00" />
                <RESULT eventid="98988" points="408" reactiontime="+87" swimtime="00:01:03.22" resultid="103235" heatid="105223" lane="2" entrytime="00:01:03.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99170" points="344" reactiontime="+75" swimtime="00:00:31.99" resultid="103236" heatid="105271" lane="9" entrytime="00:00:32.50" />
                <RESULT eventid="99218" points="313" reactiontime="+85" swimtime="00:02:30.21" resultid="103237" heatid="105301" lane="3" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                    <SPLIT distance="100" swimtime="00:01:12.55" />
                    <SPLIT distance="150" swimtime="00:01:52.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="290" reactiontime="+91" swimtime="00:05:32.24" resultid="103238" heatid="106062" lane="2" entrytime="00:05:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.49" />
                    <SPLIT distance="100" swimtime="00:01:20.65" />
                    <SPLIT distance="150" swimtime="00:02:03.49" />
                    <SPLIT distance="200" swimtime="00:02:46.12" />
                    <SPLIT distance="250" swimtime="00:03:28.54" />
                    <SPLIT distance="300" swimtime="00:04:12.19" />
                    <SPLIT distance="350" swimtime="00:04:53.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-01" firstname="Vladimir" gender="M" lastname="CHEKUTOV" nation="RUS" swrid="4754737" athleteid="103239">
              <RESULTS>
                <RESULT eventid="98798" points="387" reactiontime="+87" swimtime="00:00:28.67" resultid="103240" heatid="105138" lane="0" entrytime="00:00:28.30" />
                <RESULT eventid="98924" points="353" reactiontime="+82" swimtime="00:00:33.99" resultid="103241" heatid="105186" lane="5" entrytime="00:00:35.50" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="103242" heatid="105223" lane="7" entrytime="00:01:03.40" />
                <RESULT eventid="99186" status="DNS" swimtime="00:00:00.00" resultid="103243" heatid="105286" lane="1" entrytime="00:01:14.15" />
                <RESULT eventid="99393" status="DNS" swimtime="00:00:00.00" resultid="103244" heatid="105341" lane="0" entrytime="00:02:45.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Aleksandr" gender="M" lastname="SMIRNOV" nation="RUS" athleteid="103245">
              <RESULTS>
                <RESULT eventid="98891" points="366" swimtime="00:20:17.22" resultid="103246" heatid="105421" lane="3" entrytime="00:20:29.00" />
                <RESULT eventid="98988" points="419" reactiontime="+81" swimtime="00:01:02.68" resultid="103247" heatid="105223" lane="8" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="386" reactiontime="+86" swimtime="00:02:20.05" resultid="103248" heatid="105302" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                    <SPLIT distance="100" swimtime="00:01:07.82" />
                    <SPLIT distance="150" swimtime="00:01:44.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="383" reactiontime="+91" swimtime="00:05:02.90" resultid="103249" heatid="106062" lane="4" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.71" />
                    <SPLIT distance="100" swimtime="00:01:13.55" />
                    <SPLIT distance="150" swimtime="00:01:52.36" />
                    <SPLIT distance="200" swimtime="00:02:31.87" />
                    <SPLIT distance="250" swimtime="00:03:10.09" />
                    <SPLIT distance="300" swimtime="00:03:48.79" />
                    <SPLIT distance="350" swimtime="00:04:26.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-01" firstname="Boris" gender="M" lastname="KONKIN" nation="RUS" swrid="4776798" athleteid="103250">
              <RESULTS>
                <RESULT eventid="98798" points="449" reactiontime="+88" swimtime="00:00:27.30" resultid="103251" heatid="105141" lane="3" entrytime="00:00:26.50" />
                <RESULT eventid="98988" points="512" reactiontime="+91" swimtime="00:00:58.60" resultid="103252" heatid="105227" lane="3" entrytime="00:00:57.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99218" points="456" reactiontime="+85" swimtime="00:02:12.50" resultid="103253" heatid="105305" lane="6" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.20" />
                    <SPLIT distance="100" swimtime="00:01:02.75" />
                    <SPLIT distance="150" swimtime="00:01:36.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99473" points="421" reactiontime="+96" swimtime="00:04:53.46" resultid="103254" heatid="106060" lane="4" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                    <SPLIT distance="100" swimtime="00:01:12.64" />
                    <SPLIT distance="150" swimtime="00:01:50.90" />
                    <SPLIT distance="200" swimtime="00:02:29.94" />
                    <SPLIT distance="250" swimtime="00:03:07.38" />
                    <SPLIT distance="300" swimtime="00:03:44.24" />
                    <SPLIT distance="350" swimtime="00:04:19.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-01" firstname="Aleksandr" gender="M" lastname="MASLAKOV" nation="RUS" athleteid="103255">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="103256" heatid="105137" lane="4" entrytime="00:00:28.40" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="103257" heatid="105223" lane="1" entrytime="00:01:03.50" />
                <RESULT eventid="99091" status="DNS" swimtime="00:00:00.00" resultid="103258" heatid="105256" lane="3" entrytime="00:01:19.50" />
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="103259" heatid="105272" lane="5" entrytime="00:00:30.90" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="103260" heatid="105360" lane="3" entrytime="00:00:34.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-01" firstname="Sergey" gender="M" lastname="BOLGOV" nation="RUS" swrid="4754739" athleteid="103261">
              <RESULTS>
                <RESULT eventid="98798" status="DNS" swimtime="00:00:00.00" resultid="103262" heatid="105139" lane="0" entrytime="00:00:27.60" />
                <RESULT eventid="98988" status="DNS" swimtime="00:00:00.00" resultid="103263" heatid="105224" lane="3" entrytime="00:01:01.80" />
                <RESULT eventid="99170" status="DNS" swimtime="00:00:00.00" resultid="103264" heatid="105271" lane="8" entrytime="00:00:32.40" />
                <RESULT eventid="99425" status="DNS" swimtime="00:00:00.00" resultid="103265" heatid="105359" lane="1" entrytime="00:00:36.40" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Zvezdy Rossii C" number="1">
              <RESULTS>
                <RESULT eventid="99059" points="324" reactiontime="+83" swimtime="00:02:15.90" resultid="103278" heatid="105241" lane="5" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                    <SPLIT distance="100" swimtime="00:01:13.22" />
                    <SPLIT distance="150" swimtime="00:01:45.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103245" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="103255" number="2" reactiontime="+33" />
                    <RELAYPOSITION athleteid="103232" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="103261" number="4" reactiontime="+52" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" points="342" reactiontime="+90" swimtime="00:02:01.29" resultid="103283" heatid="105310" lane="5" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.36" />
                    <SPLIT distance="100" swimtime="00:00:59.66" />
                    <SPLIT distance="150" swimtime="00:01:31.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103245" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="103255" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="103232" number="3" reactiontime="+76" />
                    <RELAYPOSITION athleteid="103261" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="Zvezdy Rossii D" number="1">
              <RESULTS>
                <RESULT eventid="99059" points="360" reactiontime="+92" swimtime="00:02:11.31" resultid="103275" heatid="105241" lane="2" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                    <SPLIT distance="100" swimtime="00:01:13.59" />
                    <SPLIT distance="150" swimtime="00:01:44.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103239" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="103186" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="103198" number="3" reactiontime="+15" />
                    <RELAYPOSITION athleteid="103250" number="4" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" points="384" reactiontime="+84" swimtime="00:01:56.64" resultid="103276" heatid="105310" lane="1" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.70" />
                    <SPLIT distance="100" swimtime="00:01:01.23" />
                    <SPLIT distance="150" swimtime="00:01:29.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103239" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="103186" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="103198" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="103250" number="4" reactiontime="+51" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" name="Zvezdy Rossii E" number="1">
              <RESULTS>
                <RESULT eventid="99059" points="226" reactiontime="+75" swimtime="00:02:33.29" resultid="103273" heatid="105240" lane="7" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.15" />
                    <SPLIT distance="100" swimtime="00:01:23.89" />
                    <SPLIT distance="150" swimtime="00:02:03.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103180" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="103227" number="2" reactiontime="+85" />
                    <RELAYPOSITION athleteid="103161" number="3" />
                    <RELAYPOSITION athleteid="103147" number="4" reactiontime="+68" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99250" points="257" reactiontime="+98" swimtime="00:02:13.45" resultid="103274" heatid="105309" lane="7" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.67" />
                    <SPLIT distance="100" swimtime="00:01:03.21" />
                    <SPLIT distance="150" swimtime="00:01:39.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103180" number="1" reactiontime="+98" />
                    <RELAYPOSITION athleteid="103227" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="103161" number="3" reactiontime="+65" />
                    <RELAYPOSITION athleteid="103147" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" name="Zvezdy Rossii C" number="1">
              <RESULTS>
                <RESULT eventid="99036" points="426" reactiontime="+90" swimtime="00:02:20.85" resultid="103270" heatid="105238" lane="3" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.05" />
                    <SPLIT distance="100" swimtime="00:01:22.22" />
                    <SPLIT distance="150" swimtime="00:01:52.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103136" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="103086" number="2" reactiontime="+43" />
                    <RELAYPOSITION athleteid="103141" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="103118" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99234" points="528" reactiontime="+91" swimtime="00:01:59.69" resultid="103271" heatid="105307" lane="4" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.56" />
                    <SPLIT distance="100" swimtime="00:01:02.98" />
                    <SPLIT distance="150" swimtime="00:01:31.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103136" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="103086" number="2" reactiontime="+45" />
                    <RELAYPOSITION athleteid="103141" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="103118" number="4" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="Zvezdy Rossii D" number="1">
              <RESULTS>
                <RESULT eventid="99036" points="306" reactiontime="+72" swimtime="00:02:37.34" resultid="103272" heatid="105238" lane="1" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.67" />
                    <SPLIT distance="100" swimtime="00:01:24.92" />
                    <SPLIT distance="150" swimtime="00:02:01.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103098" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="103081" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="103129" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="103093" number="4" reactiontime="+72" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99234" points="335" reactiontime="+75" swimtime="00:02:19.26" resultid="103277" heatid="105307" lane="8" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                    <SPLIT distance="100" swimtime="00:01:10.73" />
                    <SPLIT distance="150" swimtime="00:01:43.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103098" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="103081" number="2" reactiontime="+67" />
                    <RELAYPOSITION athleteid="103129" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="103093" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="Zvezdy Rossii B" number="1">
              <RESULTS>
                <RESULT eventid="98846" status="DNS" swimtime="00:00:00.00" resultid="103281" heatid="105161" lane="3" entrytime="00:01:57.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103239" number="1" />
                    <RELAYPOSITION athleteid="103255" number="2" />
                    <RELAYPOSITION athleteid="103136" number="3" />
                    <RELAYPOSITION athleteid="103141" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" status="DNS" swimtime="00:00:00.00" resultid="103282" heatid="105365" lane="6" entrytime="00:02:12.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103239" number="1" />
                    <RELAYPOSITION athleteid="103255" number="2" />
                    <RELAYPOSITION athleteid="103136" number="3" />
                    <RELAYPOSITION athleteid="103141" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Zvezdy Rossii C" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="384" reactiontime="+99" swimtime="00:01:56.73" resultid="103266" heatid="105161" lane="0" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.66" />
                    <SPLIT distance="100" swimtime="00:00:57.56" />
                    <SPLIT distance="150" swimtime="00:01:30.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103123" number="1" reactiontime="+99" />
                    <RELAYPOSITION athleteid="103245" number="2" reactiontime="+43" />
                    <RELAYPOSITION athleteid="103129" number="3" reactiontime="+64" />
                    <RELAYPOSITION athleteid="103250" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" points="323" reactiontime="+88" swimtime="00:02:16.05" resultid="103267" heatid="105364" lane="4" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.99" />
                    <SPLIT distance="100" swimtime="00:01:14.82" />
                    <SPLIT distance="150" swimtime="00:01:49.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103123" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="103245" number="2" reactiontime="+75" />
                    <RELAYPOSITION athleteid="103129" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="103250" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Zvezdy Rossii D" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="350" reactiontime="+94" swimtime="00:02:00.37" resultid="103279" heatid="105161" lane="9" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                    <SPLIT distance="100" swimtime="00:01:01.99" />
                    <SPLIT distance="150" swimtime="00:01:32.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103098" number="1" reactiontime="+94" />
                    <RELAYPOSITION athleteid="103232" number="2" />
                    <RELAYPOSITION athleteid="103198" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="103118" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" points="333" reactiontime="+67" swimtime="00:02:14.73" resultid="103280" heatid="105364" lane="5" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.16" />
                    <SPLIT distance="100" swimtime="00:01:16.22" />
                    <SPLIT distance="150" swimtime="00:01:47.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103098" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="103232" number="2" reactiontime="-1" />
                    <RELAYPOSITION athleteid="103198" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="103118" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" name="Zvezdy Rossii E" number="1">
              <RESULTS>
                <RESULT eventid="98846" points="230" reactiontime="+89" swimtime="00:02:18.45" resultid="103268" heatid="105160" lane="9" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                    <SPLIT distance="100" swimtime="00:01:10.66" />
                    <SPLIT distance="150" swimtime="00:01:44.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103186" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="103081" number="2" />
                    <RELAYPOSITION athleteid="103086" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="103147" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="99441" points="190" reactiontime="+100" swimtime="00:02:42.48" resultid="103269" heatid="105364" lane="0" entrytime="00:02:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.45" />
                    <SPLIT distance="100" swimtime="00:01:29.83" />
                    <SPLIT distance="150" swimtime="00:02:08.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="103186" number="1" reactiontime="+100" />
                    <RELAYPOSITION athleteid="103081" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="103086" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="103147" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="04114" nation="POL" clubid="101565" name="Śródmiejski UKS Polna Warszawa" shortname="Śródmiejski U.K.S.Polna Warsza">
          <CONTACT city="Warszawa" name="Piotr Przybylski" phone="501704665" street="ul Polna 7a" zip="00-625" />
          <ATHLETES>
            <ATHLETE birthdate="1947-05-18" firstname="Barbara" gender="F" lastname="ŁOWKIS" nation="POL" swrid="4992752" athleteid="101566">
              <RESULTS>
                <RESULT eventid="98777" points="206" reactiontime="+134" swimtime="00:00:40.16" resultid="101567" heatid="105114" lane="0" entrytime="00:00:43.26" entrycourse="SCM" />
                <RESULT eventid="98907" points="165" reactiontime="+89" swimtime="00:00:49.27" resultid="101568" heatid="105174" lane="0" entrytime="00:00:47.28" />
                <RESULT eventid="98972" points="131" reactiontime="+124" swimtime="00:01:42.43" resultid="101569" heatid="105205" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="99314" points="140" reactiontime="+81" swimtime="00:01:51.87" resultid="101570" heatid="105277" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
  <TIMESTANDARDLISTS>
    <TIMESTANDARDLIST timestandardlistid="1077" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="29" agemin="25" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:32.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:30.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:13:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:38.75">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:43.75">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:37.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:22.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:36.75">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:22.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:20.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1103" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="29" agemin="25" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:28.25">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:07.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:22.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:15.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:11:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:21:30.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:34.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:42.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:36.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:22.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:57.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:32.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:50.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1075" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="34" agemin="30" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:33.75">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:22.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:52.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:45.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:13:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:40.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:10.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:38.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:22.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1101" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="34" agemin="30" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:29.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:25.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:22.50">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:11:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:22:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:35.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:17.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:37.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:05.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:33.75">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:17.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:52.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1073" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="39" agemin="35" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:35.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:14:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:42.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:35.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:20.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:47.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:40.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:40.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:40.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1099" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="39" agemin="35" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:30.75">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:12.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:30.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:12:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:22:30.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:37.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:52.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:38.75">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:27.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:12.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:35.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:10.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1071" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="44" agemin="40" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:37.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:27.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:07.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:15.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:15:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:50.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:42.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:35.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:40.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:50.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1097" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="44" agemin="40" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:32.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:17.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:37.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:45.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:12:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:38.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:40.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:20.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:37.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:22.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:10.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:20.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1069" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="49" agemin="45" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:40.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:30.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:15:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:52.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:55.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:50.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1095" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="49" agemin="45" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:33.75">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:13:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:40.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:10.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:42.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:35.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:40.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:20.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1067" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="54" agemin="50" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:42.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:37.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:45.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:16:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:55.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:10.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:55.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1093" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="54" agemin="50" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:35.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:52.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:15.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:13:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:42.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:35.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:20.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:42.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1065" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="59" agemin="55" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:08:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:16:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:10.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:57.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:10.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:55.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1091" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="59" agemin="55" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:37.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:30.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:14:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1063" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="64" agemin="60" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:52.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:08:30.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:20.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:20.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:10.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1089" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="64" agemin="60" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:40.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:35.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:45.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:15:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:55.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1059" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="74" agemin="70" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:00.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:21.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:30.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:20:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1085" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="74" agemin="70" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:08:15.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:20.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:02.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1057" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="79" agemin="75" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:05.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:20.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:21:15.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:27.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:17.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1083" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="79" agemin="75" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:08:45.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:18:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:22.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1615" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="84" agemin="80" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:55.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:57.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:30.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:19:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:17.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:17.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1617" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="84" agemin="80" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:10.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:45.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:23:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:05.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1619" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="89" agemin="85" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:00.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:05.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:15.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:20:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1621" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="89" agemin="85" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:15.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:12:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:24:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:35.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1623" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="94" agemin="90" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:10.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:11:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:23:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:37.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1625" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="94" agemin="90" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:20.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:13:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:26:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:08:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:08:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:08:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:08:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1627" course="LCM" gender="M" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="-1" agemin="95" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:22.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:13:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:27:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:08:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1629" course="LCM" gender="F" name="Time standard 1" type="MAXIMUM">
      <AGEGROUP agemax="-1" agemin="95" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:14:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:29:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:15.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:55.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1061" course="LCM" gender="F" type="DEFAULT">
      <AGEGROUP agemax="69" agemin="65" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:55.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:15:45.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:12.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:17.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1087" course="LCM" gender="M" type="DEFAULT">
      <AGEGROUP agemax="69" agemin="65" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:42.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:30.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:16:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:55.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:10.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:55.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
  </TIMESTANDARDLISTS>
</LENEX>

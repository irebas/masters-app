<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Tomasz Bachórz" version="11.72268">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Łódź" name="Puchar Polski Masters Łódź 2022" course="LCM" deadline="2022-03-25" organizer="MUKS Zgierz" reservecount="2" startmethod="1" timing="AUTOMATIC" nation="POL">
      <AGEDATE value="2022-04-10" type="YEAR" />
      <POOL lanemax="9" />
      <FACILITY city="Łódź" nation="POL" />
      <POINTTABLE pointtableid="3015" name="FINA Point Scoring" version="2022" />
      <QUALIFY from="2021-01-01" until="2022-04-08" />
      <SESSIONS>
        <SESSION date="2022-04-09" daytime="14:00" endtime="17:57" name="BLOK I" number="1" warmupfrom="13:00" warmupuntil="13:45">
          <EVENTS>
            <EVENT eventid="1059" gender="F" number="1" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1060" agemax="24" agemin="20" name="&quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2110" />
                    <RANKING order="2" place="2" resultid="2474" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1062" agemax="29" agemin="25" name="&quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1719" />
                    <RANKING order="2" place="2" resultid="2715" />
                    <RANKING order="3" place="3" resultid="1714" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1063" agemax="34" agemin="30" name="&quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2639" />
                    <RANKING order="2" place="2" resultid="2783" />
                    <RANKING order="3" place="3" resultid="2278" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1064" agemax="39" agemin="35" name="&quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2710" />
                    <RANKING order="2" place="2" resultid="1568" />
                    <RANKING order="3" place="3" resultid="1825" />
                    <RANKING order="4" place="4" resultid="1830" />
                    <RANKING order="5" place="5" resultid="2262" />
                    <RANKING order="6" place="-1" resultid="2094" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="44" agemin="40" name="&quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1860" />
                    <RANKING order="2" place="2" resultid="2091" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2507" />
                    <RANKING order="2" place="2" resultid="2512" />
                    <RANKING order="3" place="3" resultid="2764" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2503" />
                    <RANKING order="2" place="2" resultid="1576" />
                    <RANKING order="3" place="3" resultid="1546" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1068" agemax="59" agemin="55" name="&quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2273" />
                    <RANKING order="2" place="2" resultid="2006" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2498" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="69" agemin="65" name="&quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1941" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="74" agemin="70" name="&quot;J&quot; 70-74" />
                <AGEGROUP agegroupid="1072" agemax="79" agemin="75" name="&quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="1073" agemax="84" agemin="80" name="&quot;L&quot; 80-84" />
                <AGEGROUP agegroupid="1074" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="1075" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
                <AGEGROUP agegroupid="3984" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2503" />
                    <RANKING order="2" place="2" resultid="2273" />
                    <RANKING order="3" place="3" resultid="1719" />
                    <RANKING order="4" place="4" resultid="2639" />
                    <RANKING order="5" place="5" resultid="2507" />
                    <RANKING order="6" place="6" resultid="2498" />
                    <RANKING order="7" place="7" resultid="2710" />
                    <RANKING order="8" place="8" resultid="2715" />
                    <RANKING order="9" place="9" resultid="2783" />
                    <RANKING order="10" place="10" resultid="2278" />
                    <RANKING order="11" place="11" resultid="1568" />
                    <RANKING order="12" place="12" resultid="1714" />
                    <RANKING order="13" place="13" resultid="1825" />
                    <RANKING order="14" place="14" resultid="2512" />
                    <RANKING order="15" place="15" resultid="1576" />
                    <RANKING order="16" place="16" resultid="2764" />
                    <RANKING order="17" place="17" resultid="1830" />
                    <RANKING order="18" place="18" resultid="1860" />
                    <RANKING order="19" place="19" resultid="2262" />
                    <RANKING order="20" place="20" resultid="2006" />
                    <RANKING order="21" place="21" resultid="2091" />
                    <RANKING order="22" place="22" resultid="1941" />
                    <RANKING order="23" place="23" resultid="1546" />
                    <RANKING order="24" place="24" resultid="2110" />
                    <RANKING order="25" place="24" resultid="2474" />
                    <RANKING order="26" place="-1" resultid="2094" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2836" daytime="14:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2837" daytime="14:12" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2838" daytime="14:13" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1076" gender="M" number="2" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3810" agemax="24" agemin="20" name="&quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1788" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3811" agemax="29" agemin="25" name="&quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2052" />
                    <RANKING order="2" place="2" resultid="1573" />
                    <RANKING order="3" place="3" resultid="1704" />
                    <RANKING order="4" place="4" resultid="2435" />
                    <RANKING order="5" place="5" resultid="1868" />
                    <RANKING order="6" place="6" resultid="1709" />
                    <RANKING order="7" place="-1" resultid="2013" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3812" agemax="34" agemin="30" name="&quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2018" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3813" agemax="39" agemin="35" name="&quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2078" />
                    <RANKING order="2" place="2" resultid="2530" />
                    <RANKING order="3" place="3" resultid="2425" />
                    <RANKING order="4" place="4" resultid="2649" />
                    <RANKING order="5" place="5" resultid="2521" />
                    <RANKING order="6" place="-1" resultid="1893" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3814" agemax="44" agemin="40" name="&quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2176" />
                    <RANKING order="2" place="2" resultid="2621" />
                    <RANKING order="3" place="3" resultid="1592" />
                    <RANKING order="4" place="4" resultid="1820" />
                    <RANKING order="5" place="5" resultid="1842" />
                    <RANKING order="6" place="6" resultid="1851" />
                    <RANKING order="7" place="7" resultid="1883" />
                    <RANKING order="8" place="8" resultid="2041" />
                    <RANKING order="9" place="9" resultid="2074" />
                    <RANKING order="10" place="10" resultid="2045" />
                    <RANKING order="11" place="11" resultid="2037" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3815" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2725" />
                    <RANKING order="2" place="2" resultid="1743" />
                    <RANKING order="3" place="3" resultid="2180" />
                    <RANKING order="4" place="4" resultid="2730" />
                    <RANKING order="5" place="5" resultid="2654" />
                    <RANKING order="6" place="6" resultid="2720" />
                    <RANKING order="7" place="7" resultid="2454" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3816" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2283" />
                    <RANKING order="2" place="2" resultid="2525" />
                    <RANKING order="3" place="3" resultid="2430" />
                    <RANKING order="4" place="4" resultid="2449" />
                    <RANKING order="5" place="5" resultid="1749" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3817" agemax="59" agemin="55" name="&quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1971" />
                    <RANKING order="2" place="2" resultid="2419" />
                    <RANKING order="3" place="3" resultid="1612" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3818" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2288" />
                    <RANKING order="2" place="2" resultid="1551" />
                    <RANKING order="3" place="3" resultid="2267" />
                    <RANKING order="4" place="4" resultid="2293" />
                    <RANKING order="5" place="5" resultid="2644" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3819" agemax="69" agemin="65" name="&quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2517" />
                    <RANKING order="2" place="2" resultid="1655" />
                    <RANKING order="3" place="3" resultid="1557" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3820" agemax="74" agemin="70" name="&quot;J&quot; 70-74" />
                <AGEGROUP agegroupid="3821" agemax="79" agemin="75" name="&quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2298" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3822" agemax="84" agemin="80" name="&quot;L&quot; 80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1645" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3823" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="3824" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
                <AGEGROUP agegroupid="3985" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2725" />
                    <RANKING order="2" place="2" resultid="2052" />
                    <RANKING order="3" place="3" resultid="2078" />
                    <RANKING order="4" place="4" resultid="1573" />
                    <RANKING order="5" place="5" resultid="1704" />
                    <RANKING order="6" place="6" resultid="2176" />
                    <RANKING order="7" place="7" resultid="2530" />
                    <RANKING order="8" place="8" resultid="2283" />
                    <RANKING order="9" place="9" resultid="1743" />
                    <RANKING order="10" place="10" resultid="2288" />
                    <RANKING order="11" place="11" resultid="2621" />
                    <RANKING order="12" place="12" resultid="2435" />
                    <RANKING order="13" place="13" resultid="2180" />
                    <RANKING order="14" place="14" resultid="2425" />
                    <RANKING order="15" place="15" resultid="1592" />
                    <RANKING order="16" place="16" resultid="2517" />
                    <RANKING order="17" place="17" resultid="1820" />
                    <RANKING order="18" place="18" resultid="2730" />
                    <RANKING order="19" place="19" resultid="1868" />
                    <RANKING order="20" place="20" resultid="1842" />
                    <RANKING order="21" place="21" resultid="1851" />
                    <RANKING order="22" place="22" resultid="2649" />
                    <RANKING order="23" place="23" resultid="2018" />
                    <RANKING order="24" place="24" resultid="2654" />
                    <RANKING order="25" place="25" resultid="2525" />
                    <RANKING order="26" place="26" resultid="1883" />
                    <RANKING order="27" place="27" resultid="2720" />
                    <RANKING order="28" place="28" resultid="2430" />
                    <RANKING order="29" place="29" resultid="1709" />
                    <RANKING order="30" place="30" resultid="2041" />
                    <RANKING order="31" place="31" resultid="1971" />
                    <RANKING order="32" place="32" resultid="1551" />
                    <RANKING order="33" place="33" resultid="2419" />
                    <RANKING order="34" place="34" resultid="2449" />
                    <RANKING order="35" place="35" resultid="2298" />
                    <RANKING order="36" place="36" resultid="2074" />
                    <RANKING order="37" place="37" resultid="2267" />
                    <RANKING order="38" place="38" resultid="1655" />
                    <RANKING order="39" place="39" resultid="2293" />
                    <RANKING order="40" place="40" resultid="1612" />
                    <RANKING order="41" place="41" resultid="2454" />
                    <RANKING order="42" place="42" resultid="1749" />
                    <RANKING order="43" place="43" resultid="2045" />
                    <RANKING order="44" place="44" resultid="1557" />
                    <RANKING order="45" place="45" resultid="2037" />
                    <RANKING order="46" place="46" resultid="2644" />
                    <RANKING order="47" place="47" resultid="1645" />
                    <RANKING order="48" place="48" resultid="2521" />
                    <RANKING order="49" place="49" resultid="1788" />
                    <RANKING order="50" place="-1" resultid="1893" />
                    <RANKING order="51" place="-1" resultid="2013" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2839" daytime="14:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2840" daytime="14:17" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2841" daytime="14:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2842" daytime="14:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2843" daytime="14:21" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2844" daytime="14:22" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1092" gender="F" number="3" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3825" agemax="24" agemin="20" name="&quot;0&quot; 20-24" />
                <AGEGROUP agegroupid="3826" agemax="29" agemin="25" name="&quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2479" />
                    <RANKING order="2" place="2" resultid="2825" />
                    <RANKING order="3" place="3" resultid="2659" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3827" agemax="34" agemin="30" name="&quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2625" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3828" agemax="39" agemin="35" name="&quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1569" />
                    <RANKING order="2" place="2" resultid="2064" />
                    <RANKING order="3" place="3" resultid="2210" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3829" agemax="44" agemin="40" name="&quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2303" />
                    <RANKING order="2" place="2" resultid="2788" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3830" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2459" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3831" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2831" />
                    <RANKING order="2" place="2" resultid="1878" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3832" agemax="59" agemin="55" name="&quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2361" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3833" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2366" />
                    <RANKING order="2" place="-1" resultid="2613" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3834" agemax="69" agemin="65" name="&quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1873" />
                    <RANKING order="2" place="2" resultid="1755" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3835" agemax="74" agemin="70" name="&quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1650" />
                    <RANKING order="2" place="2" resultid="1932" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3836" agemax="79" agemin="75" name="&quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="3837" agemax="84" agemin="80" name="&quot;L&quot; 80-84" />
                <AGEGROUP agegroupid="3838" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="3839" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2845" daytime="14:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2846" daytime="14:27" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1108" gender="M" number="4" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3840" agemax="24" agemin="20" name="&quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1983" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3841" agemax="29" agemin="25" name="&quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2484" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3842" agemax="34" agemin="30" name="&quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2308" />
                    <RANKING order="2" place="2" resultid="2465" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3843" agemax="39" agemin="35" name="&quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="2663" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3844" agemax="44" agemin="40" name="&quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1811" />
                    <RANKING order="2" place="2" resultid="1888" />
                    <RANKING order="3" place="3" resultid="2380" />
                    <RANKING order="4" place="4" resultid="2733" />
                    <RANKING order="5" place="5" resultid="2793" />
                    <RANKING order="6" place="6" resultid="1761" />
                    <RANKING order="7" place="-1" resultid="2672" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3845" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2440" />
                    <RANKING order="2" place="2" resultid="1921" />
                    <RANKING order="3" place="3" resultid="2069" />
                    <RANKING order="4" place="4" resultid="1798" />
                    <RANKING order="5" place="-1" resultid="2462" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3846" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2317" />
                    <RANKING order="2" place="2" resultid="1805" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3847" agemax="59" agemin="55" name="&quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2667" />
                    <RANKING order="2" place="2" resultid="2376" />
                    <RANKING order="3" place="3" resultid="2214" />
                    <RANKING order="4" place="4" resultid="1783" />
                    <RANKING order="5" place="5" resultid="1562" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3848" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2628" />
                    <RANKING order="2" place="2" resultid="1966" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3849" agemax="69" agemin="65" name="&quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2677" />
                    <RANKING order="2" place="2" resultid="1958" />
                    <RANKING order="3" place="3" resultid="2312" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3850" agemax="74" agemin="70" name="&quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1951" />
                    <RANKING order="2" place="2" resultid="1955" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3851" agemax="79" agemin="75" name="&quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2371" />
                    <RANKING order="2" place="2" resultid="1737" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3852" agemax="84" agemin="80" name="&quot;L&quot; 80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1774" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3853" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="3854" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2847" daytime="14:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2848" daytime="14:33" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2849" daytime="14:37" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2850" daytime="14:40" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1124" gender="F" number="5" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3855" agemax="24" agemin="20" name="&quot;0&quot; 20-24" />
                <AGEGROUP agegroupid="3856" agemax="29" agemin="25" name="&quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2716" />
                    <RANKING order="2" place="2" resultid="2780" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3857" agemax="34" agemin="30" name="&quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2640" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3858" agemax="39" agemin="35" name="&quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2633" />
                    <RANKING order="2" place="2" resultid="2774" />
                    <RANKING order="3" place="3" resultid="2322" />
                    <RANKING order="4" place="-1" resultid="2096" />
                    <RANKING order="5" place="-1" resultid="2684" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3859" agemax="44" agemin="40" name="&quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2538" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3860" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2508" />
                    <RANKING order="2" place="2" resultid="2533" />
                    <RANKING order="3" place="3" resultid="2234" />
                    <RANKING order="4" place="4" resultid="2760" />
                    <RANKING order="5" place="5" resultid="2390" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3861" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2194" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3862" agemax="59" agemin="55" name="&quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2274" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3863" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2499" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3864" agemax="69" agemin="65" name="&quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2395" />
                    <RANKING order="2" place="2" resultid="1769" />
                    <RANKING order="3" place="3" resultid="2385" />
                    <RANKING order="4" place="4" resultid="1942" />
                    <RANKING order="5" place="5" resultid="1946" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3865" agemax="74" agemin="70" name="&quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1665" />
                    <RANKING order="2" place="2" resultid="1933" />
                    <RANKING order="3" place="-1" resultid="2681" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3866" agemax="79" agemin="75" name="&quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="3867" agemax="84" agemin="80" name="&quot;L&quot; 80-84" />
                <AGEGROUP agegroupid="3868" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="3869" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2851" daytime="14:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2852" daytime="14:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2853" daytime="14:45" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1140" gender="M" number="6" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3870" agemax="24" agemin="20" name="&quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1608" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3871" agemax="29" agemin="25" name="&quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2127" />
                    <RANKING order="2" place="2" resultid="1699" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3872" agemax="34" agemin="30" name="&quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2030" />
                    <RANKING order="2" place="2" resultid="2019" />
                    <RANKING order="3" place="3" resultid="2309" />
                    <RANKING order="4" place="-1" resultid="2022" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3873" agemax="39" agemin="35" name="&quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2531" />
                    <RANKING order="2" place="2" resultid="1846" />
                    <RANKING order="3" place="3" resultid="1536" />
                    <RANKING order="4" place="4" resultid="1598" />
                    <RANKING order="5" place="5" resultid="1584" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3874" agemax="44" agemin="40" name="&quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2404" />
                    <RANKING order="2" place="2" resultid="2561" />
                    <RANKING order="3" place="3" resultid="2239" />
                    <RANKING order="4" place="4" resultid="1852" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3875" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2689" />
                    <RANKING order="2" place="2" resultid="2181" />
                    <RANKING order="3" place="3" resultid="2327" />
                    <RANKING order="4" place="4" resultid="2551" />
                    <RANKING order="5" place="5" resultid="2470" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3876" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1604" />
                    <RANKING order="2" place="2" resultid="2244" />
                    <RANKING order="3" place="3" resultid="2798" />
                    <RANKING order="4" place="4" resultid="2489" />
                    <RANKING order="5" place="-1" resultid="2101" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3877" agemax="59" agemin="55" name="&quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2742" />
                    <RANKING order="2" place="2" resultid="1972" />
                    <RANKING order="3" place="3" resultid="2337" />
                    <RANKING order="4" place="4" resultid="2222" />
                    <RANKING order="5" place="5" resultid="1864" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3878" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2289" />
                    <RANKING order="2" place="2" resultid="2400" />
                    <RANKING order="3" place="3" resultid="2543" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3879" agemax="69" agemin="65" name="&quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1587" />
                    <RANKING order="2" place="2" resultid="2556" />
                    <RANKING order="3" place="-1" resultid="2249" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3880" agemax="74" agemin="70" name="&quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2758" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3881" agemax="79" agemin="75" name="&quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1738" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3882" agemax="84" agemin="80" name="&quot;L&quot; 80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1901" />
                    <RANKING order="2" place="2" resultid="2332" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3883" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="3884" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2854" daytime="14:47" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2855" daytime="14:49" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2856" daytime="14:51" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2857" daytime="14:53" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2858" daytime="14:55" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1156" gender="F" number="7" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3885" agemax="24" agemin="20" name="&quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2111" />
                    <RANKING order="2" place="2" resultid="2475" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3886" agemax="29" agemin="25" name="&quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1720" />
                    <RANKING order="2" place="2" resultid="2480" />
                    <RANKING order="3" place="3" resultid="1715" />
                    <RANKING order="4" place="4" resultid="2055" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3887" agemax="34" agemin="30" name="&quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2769" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3888" agemax="39" agemin="35" name="&quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2711" />
                    <RANKING order="2" place="2" resultid="2254" />
                    <RANKING order="3" place="3" resultid="1826" />
                    <RANKING order="4" place="4" resultid="1831" />
                    <RANKING order="5" place="5" resultid="2566" />
                    <RANKING order="6" place="6" resultid="2185" />
                    <RANKING order="7" place="7" resultid="2775" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3889" agemax="44" agemin="40" name="&quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2495" />
                    <RANKING order="2" place="2" resultid="1835" />
                    <RANKING order="3" place="3" resultid="2304" />
                    <RANKING order="4" place="4" resultid="1861" />
                    <RANKING order="5" place="5" resultid="2789" />
                    <RANKING order="6" place="6" resultid="2092" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3890" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2765" />
                    <RANKING order="2" place="2" resultid="2445" />
                    <RANKING order="3" place="3" resultid="2571" />
                    <RANKING order="4" place="-1" resultid="1766" />
                    <RANKING order="5" place="-1" resultid="2235" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3891" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2830" />
                    <RANKING order="2" place="2" resultid="1577" />
                    <RANKING order="3" place="3" resultid="1547" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3892" agemax="59" agemin="55" name="&quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2362" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3893" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2342" />
                    <RANKING order="2" place="-1" resultid="2614" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3894" agemax="69" agemin="65" name="&quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2396" />
                    <RANKING order="2" place="2" resultid="1756" />
                    <RANKING order="3" place="3" resultid="1874" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3895" agemax="74" agemin="70" name="&quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1937" />
                    <RANKING order="2" place="2" resultid="1651" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3896" agemax="79" agemin="75" name="&quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="3897" agemax="84" agemin="80" name="&quot;L&quot; 80-84" />
                <AGEGROUP agegroupid="3898" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="3899" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2859" daytime="14:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2860" daytime="14:59" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2861" daytime="15:02" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2862" daytime="15:04" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1172" gender="M" number="8" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3900" agemax="24" agemin="20" name="&quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1790" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3901" agemax="29" agemin="25" name="&quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2436" />
                    <RANKING order="2" place="2" resultid="1705" />
                    <RANKING order="3" place="3" resultid="1574" />
                    <RANKING order="4" place="4" resultid="2485" />
                    <RANKING order="5" place="5" resultid="1702" />
                    <RANKING order="6" place="6" resultid="1869" />
                    <RANKING order="7" place="7" resultid="1710" />
                    <RANKING order="8" place="8" resultid="2014" />
                    <RANKING order="9" place="9" resultid="2347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3902" agemax="34" agemin="30" name="&quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2751" />
                    <RANKING order="2" place="2" resultid="2048" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3903" agemax="39" agemin="35" name="&quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2079" />
                    <RANKING order="2" place="2" resultid="2426" />
                    <RANKING order="3" place="3" resultid="1731" />
                    <RANKING order="4" place="4" resultid="2522" />
                    <RANKING order="5" place="5" resultid="2590" />
                    <RANKING order="6" place="-1" resultid="1894" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3904" agemax="44" agemin="40" name="&quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2617" />
                    <RANKING order="2" place="2" resultid="2562" />
                    <RANKING order="3" place="3" resultid="2405" />
                    <RANKING order="4" place="4" resultid="1821" />
                    <RANKING order="5" place="5" resultid="2794" />
                    <RANKING order="6" place="6" resultid="2703" />
                    <RANKING order="7" place="7" resultid="1593" />
                    <RANKING order="8" place="8" resultid="1843" />
                    <RANKING order="9" place="9" resultid="1760" />
                    <RANKING order="10" place="10" resultid="1884" />
                    <RANKING order="11" place="11" resultid="2026" />
                    <RANKING order="12" place="12" resultid="2042" />
                    <RANKING order="13" place="13" resultid="2834" />
                    <RANKING order="14" place="14" resultid="2046" />
                    <RANKING order="15" place="15" resultid="2038" />
                    <RANKING order="16" place="16" resultid="2083" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3905" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2726" />
                    <RANKING order="2" place="2" resultid="1922" />
                    <RANKING order="3" place="3" resultid="2721" />
                    <RANKING order="4" place="4" resultid="2070" />
                    <RANKING order="5" place="5" resultid="1799" />
                    <RANKING order="6" place="6" resultid="2455" />
                    <RANKING order="7" place="7" resultid="2803" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3906" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2284" />
                    <RANKING order="2" place="2" resultid="2526" />
                    <RANKING order="3" place="3" resultid="1975" />
                    <RANKING order="4" place="4" resultid="1750" />
                    <RANKING order="5" place="5" resultid="2033" />
                    <RANKING order="6" place="6" resultid="2450" />
                    <RANKING order="7" place="7" resultid="2087" />
                    <RANKING order="8" place="-1" resultid="1988" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3907" agemax="59" agemin="55" name="&quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1779" />
                    <RANKING order="2" place="2" resultid="1613" />
                    <RANKING order="3" place="3" resultid="2215" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3908" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2694" />
                    <RANKING order="2" place="2" resultid="2580" />
                    <RANKING order="3" place="3" resultid="2746" />
                    <RANKING order="4" place="4" resultid="2645" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3909" agemax="69" agemin="65" name="&quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1588" />
                    <RANKING order="2" place="2" resultid="1656" />
                    <RANKING order="3" place="3" resultid="1924" />
                    <RANKING order="4" place="4" resultid="2585" />
                    <RANKING order="5" place="-1" resultid="1963" />
                    <RANKING order="6" place="-1" resultid="2250" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3910" agemax="74" agemin="70" name="&quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2575" />
                    <RANKING order="2" place="-1" resultid="2699" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3911" agemax="79" agemin="75" name="&quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2299" />
                    <RANKING order="2" place="2" resultid="2372" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3912" agemax="84" agemin="80" name="&quot;L&quot; 80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1646" />
                    <RANKING order="2" place="2" resultid="2333" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3913" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="3914" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2863" daytime="15:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2864" daytime="15:09" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2865" daytime="15:12" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2866" daytime="15:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2867" daytime="15:17" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2868" daytime="15:19" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="2869" daytime="15:21" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1188" gender="F" number="9" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3041" agemax="24" agemin="20" name="&quot;0&quot; 20-24" />
                <AGEGROUP agegroupid="3042" agemax="29" agemin="25" name="&quot;A&quot; 25-29" />
                <AGEGROUP agegroupid="3043" agemax="34" agemin="30" name="&quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2784" />
                    <RANKING order="2" place="-1" resultid="2279" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3044" agemax="39" agemin="35" name="&quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2066" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3045" agemax="44" agemin="40" name="&quot;D&quot; 40-44" />
                <AGEGROUP agegroupid="3046" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2513" />
                    <RANKING order="2" place="2" resultid="1815" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3047" agemax="54" agemin="50" name="&quot;F&quot; 50-54" />
                <AGEGROUP agegroupid="3048" agemax="59" agemin="55" name="&quot;G&quot; 55-59" />
                <AGEGROUP agegroupid="3049" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2351" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3050" agemax="69" agemin="65" name="&quot;I&quot; 65-69" />
                <AGEGROUP agegroupid="3051" agemax="74" agemin="70" name="&quot;J&quot; 70-74" />
                <AGEGROUP agegroupid="3052" agemax="79" agemin="75" name="&quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="3053" agemax="84" agemin="80" name="&quot;L&quot; 80-84" />
                <AGEGROUP agegroupid="3054" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="3055" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2870" daytime="15:23" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1204" gender="M" number="10" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3056" agemax="24" agemin="20" name="&quot;0&quot; 20-24" />
                <AGEGROUP agegroupid="3057" agemax="29" agemin="25" name="&quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2808" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3058" agemax="34" agemin="30" name="&quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1793" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3059" agemax="39" agemin="35" name="&quot;C&quot; 35-39" />
                <AGEGROUP agegroupid="3060" agemax="44" agemin="40" name="&quot;D&quot; 40-44" />
                <AGEGROUP agegroupid="3061" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2813" />
                    <RANKING order="2" place="2" resultid="1918" />
                    <RANKING order="3" place="3" resultid="2731" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3062" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1806" />
                    <RANKING order="2" place="2" resultid="1541" />
                    <RANKING order="3" place="-1" resultid="2431" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3063" agemax="59" agemin="55" name="&quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2420" />
                    <RANKING order="2" place="2" resultid="2226" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3064" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2268" />
                    <RANKING order="2" place="2" resultid="2294" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3065" agemax="69" agemin="65" name="&quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2518" />
                    <RANKING order="2" place="2" resultid="2593" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3066" agemax="74" agemin="70" name="&quot;J&quot; 70-74" />
                <AGEGROUP agegroupid="3067" agemax="79" agemin="75" name="&quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="3068" agemax="84" agemin="80" name="&quot;L&quot; 80-84" />
                <AGEGROUP agegroupid="3069" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="3070" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2871" daytime="15:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2872" daytime="15:32" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1220" gender="F" number="11" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3071" agemax="24" agemin="20" name="&quot;0&quot; 20-24" />
                <AGEGROUP agegroupid="3072" agemax="29" agemin="25" name="&quot;A&quot; 25-29" />
                <AGEGROUP agegroupid="3073" agemax="34" agemin="30" name="&quot;B&quot; 30-34" />
                <AGEGROUP agegroupid="3074" agemax="39" agemin="35" name="&quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2634" />
                    <RANKING order="2" place="2" resultid="2567" />
                    <RANKING order="3" place="3" resultid="2323" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3075" agemax="44" agemin="40" name="&quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2539" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3076" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2534" />
                    <RANKING order="2" place="2" resultid="1816" />
                    <RANKING order="3" place="3" resultid="2391" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3077" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2219" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3078" agemax="59" agemin="55" name="&quot;G&quot; 55-59" />
                <AGEGROUP agegroupid="3079" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2409" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3080" agemax="69" agemin="65" name="&quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1770" />
                    <RANKING order="2" place="2" resultid="2386" />
                    <RANKING order="3" place="3" resultid="1947" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3081" agemax="74" agemin="70" name="&quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1666" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3082" agemax="79" agemin="75" name="&quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="3083" agemax="84" agemin="80" name="&quot;L&quot; 80-84" />
                <AGEGROUP agegroupid="3084" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="3085" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2873" daytime="15:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2874" daytime="15:43" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1236" gender="M" number="12" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3086" agemax="24" agemin="20" name="&quot;0&quot; 20-24" />
                <AGEGROUP agegroupid="3087" agemax="29" agemin="25" name="&quot;A&quot; 25-29" />
                <AGEGROUP agegroupid="3088" agemax="34" agemin="30" name="&quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2466" />
                    <RANKING order="2" place="2" resultid="1794" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3089" agemax="39" agemin="35" name="&quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2650" />
                    <RANKING order="2" place="2" resultid="1847" />
                    <RANKING order="3" place="3" resultid="1537" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3090" agemax="44" agemin="40" name="&quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2240" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3091" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2690" />
                    <RANKING order="2" place="2" resultid="2328" />
                    <RANKING order="3" place="3" resultid="2804" />
                    <RANKING order="4" place="4" resultid="2552" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3092" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1605" />
                    <RANKING order="2" place="2" resultid="2318" />
                    <RANKING order="3" place="3" resultid="2245" />
                    <RANKING order="4" place="4" resultid="1976" />
                    <RANKING order="5" place="5" resultid="2490" />
                    <RANKING order="6" place="-1" resultid="1989" />
                    <RANKING order="7" place="-1" resultid="2103" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3093" agemax="59" agemin="55" name="&quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2754" />
                    <RANKING order="2" place="2" resultid="2227" />
                    <RANKING order="3" place="3" resultid="2223" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3094" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2401" />
                    <RANKING order="2" place="2" resultid="2581" />
                    <RANKING order="3" place="3" resultid="2544" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3095" agemax="69" agemin="65" name="&quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2313" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3096" agemax="74" agemin="70" name="&quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2598" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3097" agemax="79" agemin="75" name="&quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="3098" agemax="84" agemin="80" name="&quot;L&quot; 80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1775" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3099" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="3100" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2875" daytime="15:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2876" daytime="15:57" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2877" daytime="16:04" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1252" gender="F" number="13" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3101" agemax="24" agemin="20" name="&quot;0&quot; 20-24" />
                <AGEGROUP agegroupid="3102" agemax="29" agemin="25" name="&quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2056" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3103" agemax="34" agemin="30" name="&quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2770" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3104" agemax="39" agemin="35" name="&quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2255" />
                    <RANKING order="2" place="2" resultid="2263" />
                    <RANKING order="3" place="-1" resultid="2685" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3105" agemax="44" agemin="40" name="&quot;D&quot; 40-44" />
                <AGEGROUP agegroupid="3106" agemax="49" agemin="45" name="&quot;E&quot; 45-49" />
                <AGEGROUP agegroupid="3107" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2504" />
                    <RANKING order="2" place="2" resultid="1879" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3108" agemax="59" agemin="55" name="&quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2007" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3109" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2367" />
                    <RANKING order="2" place="2" resultid="2343" />
                    <RANKING order="3" place="3" resultid="2410" />
                    <RANKING order="4" place="-1" resultid="2352" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3110" agemax="69" agemin="65" name="&quot;I&quot; 65-69" />
                <AGEGROUP agegroupid="3111" agemax="74" agemin="70" name="&quot;J&quot; 70-74" />
                <AGEGROUP agegroupid="3112" agemax="79" agemin="75" name="&quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="3113" agemax="84" agemin="80" name="&quot;L&quot; 80-84" />
                <AGEGROUP agegroupid="3114" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="3115" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2878" daytime="16:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2879" daytime="16:14" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1268" gender="M" number="14" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3116" agemax="24" agemin="20" name="&quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1984" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3117" agemax="29" agemin="25" name="&quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2809" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3118" agemax="34" agemin="30" name="&quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2752" />
                    <RANKING order="2" place="-1" resultid="2023" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3119" agemax="39" agemin="35" name="&quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1733" />
                    <RANKING order="2" place="2" resultid="1599" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3120" agemax="44" agemin="40" name="&quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2622" />
                    <RANKING order="2" place="2" resultid="2734" />
                    <RANKING order="3" place="3" resultid="2075" />
                    <RANKING order="4" place="-1" resultid="1889" />
                    <RANKING order="5" place="-1" resultid="2381" />
                    <RANKING order="6" place="-1" resultid="2673" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3121" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2814" />
                    <RANKING order="2" place="2" resultid="1744" />
                    <RANKING order="3" place="3" resultid="2655" />
                    <RANKING order="4" place="4" resultid="1919" />
                    <RANKING order="5" place="5" resultid="2441" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3122" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2799" />
                    <RANKING order="2" place="2" resultid="1542" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3123" agemax="59" agemin="55" name="&quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2668" />
                    <RANKING order="2" place="2" resultid="2338" />
                    <RANKING order="3" place="3" resultid="1563" />
                    <RANKING order="4" place="4" resultid="1784" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3124" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2695" />
                    <RANKING order="2" place="2" resultid="2747" />
                    <RANKING order="3" place="3" resultid="1552" />
                    <RANKING order="4" place="4" resultid="1967" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3125" agemax="69" agemin="65" name="&quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1959" />
                    <RANKING order="2" place="2" resultid="2557" />
                    <RANKING order="3" place="3" resultid="1925" />
                    <RANKING order="4" place="4" resultid="1558" />
                    <RANKING order="5" place="5" resultid="2586" />
                    <RANKING order="6" place="6" resultid="2594" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3126" agemax="74" agemin="70" name="&quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2576" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3127" agemax="79" agemin="75" name="&quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="3128" agemax="84" agemin="80" name="&quot;L&quot; 80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1902" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3129" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="3130" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2880" daytime="16:19" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2881" daytime="16:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2882" daytime="16:31" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2883" daytime="16:36" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1284" gender="X" number="15" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1285" agemax="96" agemin="80" name="&quot;0&quot; 80-96" calculate="TOTAL" />
                <AGEGROUP agegroupid="1286" agemax="119" agemin="100" name="&quot;A&quot; 100-119" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1697" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1287" agemax="159" agemin="120" name="&quot;B&quot; 120-159" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2705" />
                    <RANKING order="2" place="2" resultid="2166" />
                    <RANKING order="3" place="-1" resultid="3319" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1288" agemax="199" agemin="160" name="&quot;C&quot; 160-199" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2756" />
                    <RANKING order="2" place="2" resultid="2081" />
                    <RANKING order="3" place="3" resultid="2356" />
                    <RANKING order="4" place="4" resultid="2258" />
                    <RANKING order="5" place="5" resultid="2603" />
                    <RANKING order="6" place="6" resultid="1856" />
                    <RANKING order="7" place="7" resultid="1897" />
                    <RANKING order="8" place="8" resultid="2230" />
                    <RANKING order="9" place="9" resultid="2604" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1289" agemax="239" agemin="200" name="&quot;D&quot; 200-239" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2605" />
                    <RANKING order="2" place="2" resultid="2413" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1290" agemax="279" agemin="240" name="&quot;E&quot; 240-279" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2355" />
                    <RANKING order="2" place="2" resultid="2606" />
                    <RANKING order="3" place="3" resultid="2414" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1291" agemax="9999" agemin="280" name="&quot;F&quot; 280 +" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1979" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3969" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3970" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2022-04-10" daytime="10:00" endtime="13:36" name="BLOK II" number="2" warmupfrom="09:00" warmupuntil="09:50">
          <EVENTS>
            <EVENT eventid="1301" daytime="10:00" gender="F" number="16" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3131" agemax="24" agemin="20" name="&quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2112" />
                    <RANKING order="2" place="2" resultid="2476" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3132" agemax="29" agemin="25" name="&quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1721" />
                    <RANKING order="2" place="2" resultid="2717" />
                    <RANKING order="3" place="3" resultid="2004" />
                    <RANKING order="4" place="4" resultid="1716" />
                    <RANKING order="5" place="5" resultid="2779" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3133" agemax="34" agemin="30" name="&quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2641" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3134" agemax="39" agemin="35" name="&quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2635" />
                    <RANKING order="2" place="2" resultid="2712" />
                    <RANKING order="3" place="3" resultid="2256" />
                    <RANKING order="4" place="4" resultid="1827" />
                    <RANKING order="5" place="5" resultid="2324" />
                    <RANKING order="6" place="-1" resultid="2095" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3135" agemax="44" agemin="40" name="&quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1836" />
                    <RANKING order="2" place="2" resultid="2305" />
                    <RANKING order="3" place="3" resultid="2790" />
                    <RANKING order="4" place="4" resultid="2540" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3136" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2509" />
                    <RANKING order="2" place="2" resultid="1992" />
                    <RANKING order="3" place="3" resultid="2236" />
                    <RANKING order="4" place="4" resultid="2446" />
                    <RANKING order="5" place="5" resultid="2572" />
                    <RANKING order="6" place="6" resultid="2392" />
                    <RANKING order="7" place="-1" resultid="1767" />
                    <RANKING order="8" place="-1" resultid="2761" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3137" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2828" />
                    <RANKING order="2" place="2" resultid="1578" />
                    <RANKING order="3" place="3" resultid="1548" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3138" agemax="59" agemin="55" name="&quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2275" />
                    <RANKING order="2" place="2" resultid="2008" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3139" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2500" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3140" agemax="69" agemin="65" name="&quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2397" />
                    <RANKING order="2" place="2" resultid="1771" />
                    <RANKING order="3" place="3" resultid="2387" />
                    <RANKING order="4" place="4" resultid="1948" />
                    <RANKING order="5" place="5" resultid="1943" />
                    <RANKING order="6" place="6" resultid="1875" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3141" agemax="74" agemin="70" name="&quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1938" />
                    <RANKING order="2" place="2" resultid="1652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3142" agemax="79" agemin="75" name="&quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="3143" agemax="84" agemin="80" name="&quot;L&quot; 80-84" />
                <AGEGROUP agegroupid="3144" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="3145" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2886" daytime="10:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2887" daytime="10:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2888" daytime="10:03" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2889" daytime="10:05" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1318" gender="M" number="17" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3146" agemax="24" agemin="20" name="&quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1789" />
                    <RANKING order="2" place="2" resultid="1610" />
                    <RANKING order="3" place="3" resultid="1985" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3147" agemax="29" agemin="25" name="&quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1706" />
                    <RANKING order="2" place="2" resultid="2437" />
                    <RANKING order="3" place="3" resultid="2128" />
                    <RANKING order="4" place="4" resultid="2486" />
                    <RANKING order="5" place="5" resultid="1700" />
                    <RANKING order="6" place="6" resultid="1870" />
                    <RANKING order="7" place="7" resultid="1711" />
                    <RANKING order="8" place="8" resultid="2348" />
                    <RANKING order="9" place="9" resultid="2015" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3148" agemax="34" agemin="30" name="&quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2031" />
                    <RANKING order="2" place="2" resultid="1995" />
                    <RANKING order="3" place="3" resultid="2020" />
                    <RANKING order="4" place="4" resultid="2049" />
                    <RANKING order="5" place="-1" resultid="2011" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3149" agemax="39" agemin="35" name="&quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2427" />
                    <RANKING order="2" place="2" resultid="1848" />
                    <RANKING order="3" place="3" resultid="2651" />
                    <RANKING order="4" place="4" resultid="1732" />
                    <RANKING order="5" place="5" resultid="2060" />
                    <RANKING order="6" place="6" resultid="2523" />
                    <RANKING order="7" place="7" resultid="2591" />
                    <RANKING order="8" place="8" resultid="1600" />
                    <RANKING order="9" place="-1" resultid="1895" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3150" agemax="44" agemin="40" name="&quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2674" />
                    <RANKING order="2" place="2" resultid="2618" />
                    <RANKING order="3" place="3" resultid="2177" />
                    <RANKING order="4" place="4" resultid="2563" />
                    <RANKING order="5" place="5" resultid="1822" />
                    <RANKING order="6" place="6" resultid="2406" />
                    <RANKING order="7" place="7" resultid="2382" />
                    <RANKING order="8" place="8" resultid="1594" />
                    <RANKING order="9" place="9" resultid="1844" />
                    <RANKING order="10" place="10" resultid="1853" />
                    <RANKING order="11" place="11" resultid="1885" />
                    <RANKING order="12" place="12" resultid="2818" />
                    <RANKING order="13" place="13" resultid="2027" />
                    <RANKING order="14" place="14" resultid="2043" />
                    <RANKING order="15" place="15" resultid="2076" />
                    <RANKING order="16" place="16" resultid="2084" />
                    <RANKING order="17" place="17" resultid="2833" />
                    <RANKING order="18" place="18" resultid="2039" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3151" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2691" />
                    <RANKING order="2" place="2" resultid="2463" />
                    <RANKING order="3" place="3" resultid="1839" />
                    <RANKING order="4" place="4" resultid="2722" />
                    <RANKING order="5" place="5" resultid="2329" />
                    <RANKING order="6" place="6" resultid="1800" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3152" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2285" />
                    <RANKING order="2" place="2" resultid="2432" />
                    <RANKING order="3" place="3" resultid="2527" />
                    <RANKING order="4" place="4" resultid="1977" />
                    <RANKING order="5" place="5" resultid="2034" />
                    <RANKING order="6" place="6" resultid="2246" />
                    <RANKING order="7" place="7" resultid="2451" />
                    <RANKING order="8" place="8" resultid="1751" />
                    <RANKING order="9" place="9" resultid="1543" />
                    <RANKING order="10" place="-1" resultid="2088" />
                    <RANKING order="11" place="-1" resultid="2102" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3153" agemax="59" agemin="55" name="&quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2743" />
                    <RANKING order="2" place="2" resultid="1780" />
                    <RANKING order="3" place="3" resultid="2339" />
                    <RANKING order="4" place="4" resultid="2201" />
                    <RANKING order="5" place="5" resultid="2228" />
                    <RANKING order="6" place="-1" resultid="1614" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3154" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2696" />
                    <RANKING order="2" place="2" resultid="2582" />
                    <RANKING order="3" place="3" resultid="2748" />
                    <RANKING order="4" place="4" resultid="1553" />
                    <RANKING order="5" place="5" resultid="2646" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3155" agemax="69" agemin="65" name="&quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1589" />
                    <RANKING order="2" place="2" resultid="2678" />
                    <RANKING order="3" place="3" resultid="1926" />
                    <RANKING order="4" place="4" resultid="1559" />
                    <RANKING order="5" place="5" resultid="2587" />
                    <RANKING order="6" place="6" resultid="2314" />
                    <RANKING order="7" place="-1" resultid="1964" />
                    <RANKING order="8" place="-1" resultid="2251" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3156" agemax="74" agemin="70" name="&quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2577" />
                    <RANKING order="2" place="2" resultid="2700" />
                    <RANKING order="3" place="3" resultid="1581" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3157" agemax="79" agemin="75" name="&quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2300" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3158" agemax="84" agemin="80" name="&quot;L&quot; 80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1647" />
                    <RANKING order="2" place="2" resultid="2334" />
                    <RANKING order="3" place="3" resultid="1903" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3159" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="3160" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2890" daytime="10:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2891" daytime="10:08" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2892" daytime="10:09" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2893" daytime="10:11" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2894" daytime="10:13" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2895" daytime="10:14" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="2896" daytime="10:15" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="2897" daytime="10:16" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="2898" daytime="10:18" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1334" gender="F" number="18" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3161" agemax="24" agemin="20" name="&quot;0&quot; 20-24" />
                <AGEGROUP agegroupid="3162" agemax="29" agemin="25" name="&quot;A&quot; 25-29" />
                <AGEGROUP agegroupid="3163" agemax="34" agemin="30" name="&quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2785" />
                    <RANKING order="2" place="2" resultid="2280" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3164" agemax="39" agemin="35" name="&quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2065" />
                    <RANKING order="2" place="2" resultid="1832" />
                    <RANKING order="3" place="3" resultid="2264" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3165" agemax="44" agemin="40" name="&quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1862" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3166" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2514" />
                    <RANKING order="2" place="2" resultid="2766" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3167" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2505" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3168" agemax="59" agemin="55" name="&quot;G&quot; 55-59" />
                <AGEGROUP agegroupid="3169" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2344" />
                    <RANKING order="2" place="2" resultid="2411" />
                    <RANKING order="3" place="3" resultid="2353" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3170" agemax="69" agemin="65" name="&quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1757" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3171" agemax="74" agemin="70" name="&quot;J&quot; 70-74" />
                <AGEGROUP agegroupid="3172" agemax="79" agemin="75" name="&quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="3173" agemax="84" agemin="80" name="&quot;L&quot; 80-84" />
                <AGEGROUP agegroupid="3174" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="3175" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2899" daytime="10:19" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2900" daytime="10:24" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1350" gender="M" number="19" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3176" agemax="24" agemin="20" name="&quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1791" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3177" agemax="29" agemin="25" name="&quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1707" />
                    <RANKING order="2" place="2" resultid="2810" />
                    <RANKING order="3" place="3" resultid="2438" />
                    <RANKING order="4" place="4" resultid="1871" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3178" agemax="34" agemin="30" name="&quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1795" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3179" agemax="39" agemin="35" name="&quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2080" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3180" agemax="44" agemin="40" name="&quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2178" />
                    <RANKING order="2" place="2" resultid="1823" />
                    <RANKING order="3" place="3" resultid="2623" />
                    <RANKING order="4" place="4" resultid="1595" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3181" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2815" />
                    <RANKING order="2" place="2" resultid="1745" />
                    <RANKING order="3" place="3" resultid="2656" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3182" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1807" />
                    <RANKING order="2" place="2" resultid="2800" />
                    <RANKING order="3" place="3" resultid="1544" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3183" agemax="59" agemin="55" name="&quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2421" />
                    <RANKING order="2" place="2" resultid="1564" />
                    <RANKING order="3" place="-1" resultid="1615" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3184" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2290" />
                    <RANKING order="2" place="2" resultid="2269" />
                    <RANKING order="3" place="3" resultid="2295" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3185" agemax="69" agemin="65" name="&quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2519" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3186" agemax="74" agemin="70" name="&quot;J&quot; 70-74" />
                <AGEGROUP agegroupid="3187" agemax="79" agemin="75" name="&quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="3188" agemax="84" agemin="80" name="&quot;L&quot; 80-84" />
                <AGEGROUP agegroupid="3189" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="3190" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2901" daytime="10:29" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2902" daytime="10:31" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2903" daytime="10:34" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1366" gender="F" number="20" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3191" agemax="24" agemin="20" name="&quot;0&quot; 20-24" />
                <AGEGROUP agegroupid="3192" agemax="29" agemin="25" name="&quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2660" />
                    <RANKING order="2" place="-1" resultid="2824" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3193" agemax="34" agemin="30" name="&quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2626" />
                    <RANKING order="2" place="2" resultid="2771" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3194" agemax="39" agemin="35" name="&quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2713" />
                    <RANKING order="2" place="2" resultid="1570" />
                    <RANKING order="3" place="3" resultid="2686" />
                    <RANKING order="4" place="4" resultid="2212" />
                    <RANKING order="5" place="5" resultid="2325" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3195" agemax="44" agemin="40" name="&quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2306" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3196" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2510" />
                    <RANKING order="2" place="2" resultid="2460" />
                    <RANKING order="3" place="3" resultid="1993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3197" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2829" />
                    <RANKING order="2" place="2" resultid="1880" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3198" agemax="59" agemin="55" name="&quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2009" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3199" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2501" />
                    <RANKING order="2" place="2" resultid="2368" />
                    <RANKING order="3" place="3" resultid="2354" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3200" agemax="69" agemin="65" name="&quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2398" />
                    <RANKING order="2" place="2" resultid="1944" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3201" agemax="74" agemin="70" name="&quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1939" />
                    <RANKING order="2" place="2" resultid="1653" />
                    <RANKING order="3" place="3" resultid="1667" />
                    <RANKING order="4" place="4" resultid="1934" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3202" agemax="79" agemin="75" name="&quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="3203" agemax="84" agemin="80" name="&quot;L&quot; 80-84" />
                <AGEGROUP agegroupid="3204" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="3205" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2904" daytime="10:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2905" daytime="10:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2906" daytime="10:40" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1382" gender="M" number="21" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3206" agemax="24" agemin="20" name="&quot;0&quot; 20-24" />
                <AGEGROUP agegroupid="3207" agemax="29" agemin="25" name="&quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2129" />
                    <RANKING order="2" place="2" resultid="2349" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3208" agemax="34" agemin="30" name="&quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2310" />
                    <RANKING order="2" place="2" resultid="2467" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3209" agemax="39" agemin="35" name="&quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2664" />
                    <RANKING order="2" place="2" resultid="2601" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3210" agemax="44" agemin="40" name="&quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2675" />
                    <RANKING order="2" place="2" resultid="1812" />
                    <RANKING order="3" place="3" resultid="1890" />
                    <RANKING order="4" place="4" resultid="2383" />
                    <RANKING order="5" place="5" resultid="2735" />
                    <RANKING order="6" place="6" resultid="1762" />
                    <RANKING order="7" place="7" resultid="1854" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3211" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2727" />
                    <RANKING order="2" place="2" resultid="2442" />
                    <RANKING order="3" place="3" resultid="2182" />
                    <RANKING order="4" place="4" resultid="1840" />
                    <RANKING order="5" place="5" resultid="2071" />
                    <RANKING order="6" place="6" resultid="2456" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3212" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2801" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3213" agemax="59" agemin="55" name="&quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2669" />
                    <RANKING order="2" place="2" resultid="2377" />
                    <RANKING order="3" place="3" resultid="1865" />
                    <RANKING order="4" place="4" resultid="2216" />
                    <RANKING order="5" place="5" resultid="1785" />
                    <RANKING order="6" place="6" resultid="2207" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3214" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2629" />
                    <RANKING order="2" place="2" resultid="1554" />
                    <RANKING order="3" place="3" resultid="1968" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3215" agemax="69" agemin="65" name="&quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2558" />
                    <RANKING order="2" place="2" resultid="1657" />
                    <RANKING order="3" place="3" resultid="1927" />
                    <RANKING order="4" place="4" resultid="1960" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3216" agemax="74" agemin="70" name="&quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1952" />
                    <RANKING order="2" place="2" resultid="1956" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3217" agemax="79" agemin="75" name="&quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2373" />
                    <RANKING order="2" place="2" resultid="1740" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3218" agemax="84" agemin="80" name="&quot;L&quot; 80-84" />
                <AGEGROUP agegroupid="3219" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="3220" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2907" daytime="10:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2908" daytime="10:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2909" daytime="10:46" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2910" daytime="10:47" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1398" gender="F" number="22" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3221" agemax="24" agemin="20" name="&quot;0&quot; 20-24" />
                <AGEGROUP agegroupid="3222" agemax="29" agemin="25" name="&quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2718" />
                    <RANKING order="2" place="2" resultid="2058" />
                    <RANKING order="3" place="3" resultid="2781" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3223" agemax="34" agemin="30" name="&quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2642" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3224" agemax="39" agemin="35" name="&quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2636" />
                    <RANKING order="2" place="2" resultid="2257" />
                    <RANKING order="3" place="3" resultid="2568" />
                    <RANKING order="4" place="4" resultid="2776" />
                    <RANKING order="5" place="-1" resultid="2097" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3225" agemax="44" agemin="40" name="&quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2541" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3226" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2535" />
                    <RANKING order="2" place="2" resultid="2393" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3227" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2220" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3228" agemax="59" agemin="55" name="&quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2276" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3229" agemax="64" agemin="60" name="&quot;H&quot; 60-64" />
                <AGEGROUP agegroupid="3230" agemax="69" agemin="65" name="&quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1772" />
                    <RANKING order="2" place="2" resultid="2388" />
                    <RANKING order="3" place="3" resultid="1949" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3231" agemax="74" agemin="70" name="&quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1935" />
                    <RANKING order="2" place="2" resultid="1668" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3232" agemax="79" agemin="75" name="&quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="3233" agemax="84" agemin="80" name="&quot;L&quot; 80-84" />
                <AGEGROUP agegroupid="3234" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="3235" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2911" daytime="10:49" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2912" daytime="10:52" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1414" gender="M" number="23" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3236" agemax="24" agemin="20" name="&quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1609" />
                    <RANKING order="2" place="2" resultid="1986" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3237" agemax="29" agemin="25" name="&quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1701" />
                    <RANKING order="2" place="-1" resultid="2016" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3238" agemax="34" agemin="30" name="&quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2021" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3239" agemax="39" agemin="35" name="&quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2652" />
                    <RANKING order="2" place="2" resultid="1849" />
                    <RANKING order="3" place="3" resultid="1538" />
                    <RANKING order="4" place="4" resultid="1601" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3240" agemax="44" agemin="40" name="&quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2407" />
                    <RANKING order="2" place="2" resultid="2564" />
                    <RANKING order="3" place="3" resultid="2241" />
                    <RANKING order="4" place="4" resultid="2819" />
                    <RANKING order="5" place="5" resultid="2085" />
                    <RANKING order="6" place="-1" resultid="1891" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3241" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2692" />
                    <RANKING order="2" place="2" resultid="2330" />
                    <RANKING order="3" place="3" resultid="2457" />
                    <RANKING order="4" place="4" resultid="2553" />
                    <RANKING order="5" place="5" resultid="2471" />
                    <RANKING order="6" place="6" resultid="2723" />
                    <RANKING order="7" place="7" resultid="2805" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3242" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1606" />
                    <RANKING order="2" place="2" resultid="2286" />
                    <RANKING order="3" place="3" resultid="2319" />
                    <RANKING order="4" place="4" resultid="2247" />
                    <RANKING order="5" place="5" resultid="2491" />
                    <RANKING order="6" place="-1" resultid="2104" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3243" agemax="59" agemin="55" name="&quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2744" />
                    <RANKING order="2" place="2" resultid="1973" />
                    <RANKING order="3" place="3" resultid="2340" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3244" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2402" />
                    <RANKING order="2" place="2" resultid="2296" />
                    <RANKING order="3" place="3" resultid="2545" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3245" agemax="69" agemin="65" name="&quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1590" />
                    <RANKING order="2" place="2" resultid="2559" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3246" agemax="74" agemin="70" name="&quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2599" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3247" agemax="79" agemin="75" name="&quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1739" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3248" agemax="84" agemin="80" name="&quot;L&quot; 80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1904" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3249" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="3250" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2913" daytime="10:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2914" daytime="10:58" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2915" daytime="11:01" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2916" daytime="11:03" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1430" gender="F" number="24" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3251" agemax="24" agemin="20" name="&quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2477" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3252" agemax="29" agemin="25" name="&quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1722" />
                    <RANKING order="2" place="2" resultid="2481" />
                    <RANKING order="3" place="3" resultid="1717" />
                    <RANKING order="4" place="4" resultid="2057" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3253" agemax="34" agemin="30" name="&quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2281" />
                    <RANKING order="2" place="2" resultid="2786" />
                    <RANKING order="3" place="3" resultid="2772" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3254" agemax="39" agemin="35" name="&quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1828" />
                    <RANKING order="2" place="2" resultid="2265" />
                    <RANKING order="3" place="3" resultid="1833" />
                    <RANKING order="4" place="4" resultid="2569" />
                    <RANKING order="5" place="5" resultid="2687" />
                    <RANKING order="6" place="6" resultid="2777" />
                    <RANKING order="7" place="7" resultid="2187" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3255" agemax="44" agemin="40" name="&quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2496" />
                    <RANKING order="2" place="2" resultid="1837" />
                    <RANKING order="3" place="3" resultid="2791" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3256" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2767" />
                    <RANKING order="2" place="2" resultid="2515" />
                    <RANKING order="3" place="3" resultid="2237" />
                    <RANKING order="4" place="4" resultid="1817" />
                    <RANKING order="5" place="5" resultid="2573" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3257" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2221" />
                    <RANKING order="2" place="2" resultid="1549" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3258" agemax="59" agemin="55" name="&quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2363" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3259" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2345" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3260" agemax="69" agemin="65" name="&quot;I&quot; 65-69" />
                <AGEGROUP agegroupid="3261" agemax="74" agemin="70" name="&quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2682" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3262" agemax="79" agemin="75" name="&quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="3263" agemax="84" agemin="80" name="&quot;L&quot; 80-84" />
                <AGEGROUP agegroupid="3264" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="3265" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
                <AGEGROUP agegroupid="3995" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1722" />
                    <RANKING order="2" place="2" resultid="2481" />
                    <RANKING order="3" place="3" resultid="2496" />
                    <RANKING order="4" place="4" resultid="1837" />
                    <RANKING order="5" place="5" resultid="1717" />
                    <RANKING order="6" place="6" resultid="2767" />
                    <RANKING order="7" place="7" resultid="2057" />
                    <RANKING order="8" place="8" resultid="2221" />
                    <RANKING order="9" place="9" resultid="2281" />
                    <RANKING order="10" place="10" resultid="2345" />
                    <RANKING order="11" place="11" resultid="2515" />
                    <RANKING order="12" place="12" resultid="2786" />
                    <RANKING order="13" place="13" resultid="1828" />
                    <RANKING order="14" place="14" resultid="2237" />
                    <RANKING order="15" place="15" resultid="2363" />
                    <RANKING order="16" place="16" resultid="2265" />
                    <RANKING order="17" place="17" resultid="1833" />
                    <RANKING order="18" place="18" resultid="2569" />
                    <RANKING order="19" place="19" resultid="2772" />
                    <RANKING order="20" place="20" resultid="1817" />
                    <RANKING order="21" place="21" resultid="2791" />
                    <RANKING order="22" place="22" resultid="2687" />
                    <RANKING order="23" place="23" resultid="2777" />
                    <RANKING order="24" place="24" resultid="2187" />
                    <RANKING order="25" place="25" resultid="2573" />
                    <RANKING order="26" place="26" resultid="2682" />
                    <RANKING order="27" place="27" resultid="1549" />
                    <RANKING order="28" place="28" resultid="2477" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2917" daytime="11:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2918" daytime="11:11" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2919" daytime="11:16" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1446" gender="M" number="25" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3996" agemax="24" agemin="20" name="&quot;0&quot; 20-24" />
                <AGEGROUP agegroupid="3997" agemax="29" agemin="25" name="&quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2053" />
                    <RANKING order="2" place="2" resultid="2811" />
                    <RANKING order="3" place="3" resultid="1712" />
                    <RANKING order="4" place="4" resultid="2826" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3998" agemax="34" agemin="30" name="&quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1996" />
                    <RANKING order="2" place="2" resultid="2050" />
                    <RANKING order="3" place="3" resultid="2468" />
                    <RANKING order="4" place="-1" resultid="2024" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3999" agemax="39" agemin="35" name="&quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2428" />
                    <RANKING order="2" place="2" resultid="2665" />
                    <RANKING order="3" place="3" resultid="1734" />
                    <RANKING order="4" place="4" resultid="2602" />
                    <RANKING order="5" place="5" resultid="1539" />
                    <RANKING order="6" place="6" resultid="2934" />
                    <RANKING order="7" place="-1" resultid="1896" />
                    <RANKING order="8" place="-1" resultid="2061" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4000" agemax="44" agemin="40" name="&quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2795" />
                    <RANKING order="2" place="2" resultid="2704" />
                    <RANKING order="3" place="3" resultid="2242" />
                    <RANKING order="4" place="4" resultid="2835" />
                    <RANKING order="5" place="5" resultid="2028" />
                    <RANKING order="6" place="-1" resultid="1886" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4001" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2816" />
                    <RANKING order="2" place="2" resultid="1746" />
                    <RANKING order="3" place="3" resultid="2657" />
                    <RANKING order="4" place="4" resultid="2554" />
                    <RANKING order="5" place="5" resultid="2806" />
                    <RANKING order="6" place="-1" resultid="2728" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4002" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2433" />
                    <RANKING order="2" place="2" resultid="2528" />
                    <RANKING order="3" place="3" resultid="1978" />
                    <RANKING order="4" place="4" resultid="1752" />
                    <RANKING order="5" place="5" resultid="2452" />
                    <RANKING order="6" place="6" resultid="2035" />
                    <RANKING order="7" place="-1" resultid="2089" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4003" agemax="59" agemin="55" name="&quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2670" />
                    <RANKING order="2" place="2" resultid="2378" />
                    <RANKING order="3" place="3" resultid="2755" />
                    <RANKING order="4" place="4" resultid="1781" />
                    <RANKING order="5" place="5" resultid="2422" />
                    <RANKING order="6" place="6" resultid="1565" />
                    <RANKING order="7" place="7" resultid="2225" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4004" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2697" />
                    <RANKING order="2" place="2" resultid="2749" />
                    <RANKING order="3" place="3" resultid="2647" />
                    <RANKING order="4" place="4" resultid="2270" />
                    <RANKING order="5" place="5" resultid="2583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4005" agemax="69" agemin="65" name="&quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1658" />
                    <RANKING order="2" place="2" resultid="1560" />
                    <RANKING order="3" place="3" resultid="2588" />
                    <RANKING order="4" place="4" resultid="2595" />
                    <RANKING order="5" place="-1" resultid="2252" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4006" agemax="74" agemin="70" name="&quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2701" />
                    <RANKING order="2" place="2" resultid="2578" />
                    <RANKING order="3" place="3" resultid="1582" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4007" agemax="79" agemin="75" name="&quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2301" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4008" agemax="84" agemin="80" name="&quot;L&quot; 80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1648" />
                    <RANKING order="2" place="2" resultid="2335" />
                    <RANKING order="3" place="3" resultid="1776" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4009" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="4010" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
                <AGEGROUP agegroupid="4011" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2053" />
                    <RANKING order="2" place="2" resultid="2697" />
                    <RANKING order="3" place="3" resultid="2816" />
                    <RANKING order="4" place="4" resultid="2670" />
                    <RANKING order="5" place="5" resultid="1746" />
                    <RANKING order="6" place="6" resultid="2428" />
                    <RANKING order="7" place="7" resultid="1996" />
                    <RANKING order="8" place="8" resultid="2811" />
                    <RANKING order="9" place="9" resultid="2378" />
                    <RANKING order="10" place="10" resultid="2795" />
                    <RANKING order="11" place="11" resultid="2755" />
                    <RANKING order="12" place="12" resultid="1781" />
                    <RANKING order="13" place="13" resultid="2704" />
                    <RANKING order="14" place="14" resultid="2665" />
                    <RANKING order="15" place="15" resultid="2433" />
                    <RANKING order="16" place="16" resultid="2657" />
                    <RANKING order="17" place="17" resultid="2242" />
                    <RANKING order="18" place="17" resultid="2701" />
                    <RANKING order="19" place="19" resultid="1712" />
                    <RANKING order="20" place="20" resultid="1734" />
                    <RANKING order="21" place="21" resultid="2050" />
                    <RANKING order="22" place="22" resultid="2826" />
                    <RANKING order="23" place="23" resultid="2578" />
                    <RANKING order="24" place="24" resultid="2528" />
                    <RANKING order="25" place="25" resultid="2749" />
                    <RANKING order="26" place="26" resultid="1658" />
                    <RANKING order="27" place="27" resultid="2602" />
                    <RANKING order="28" place="28" resultid="1978" />
                    <RANKING order="29" place="28" resultid="2301" />
                    <RANKING order="30" place="30" resultid="1752" />
                    <RANKING order="31" place="31" resultid="2647" />
                    <RANKING order="32" place="32" resultid="2468" />
                    <RANKING order="33" place="33" resultid="2270" />
                    <RANKING order="34" place="34" resultid="2554" />
                    <RANKING order="35" place="35" resultid="2422" />
                    <RANKING order="36" place="36" resultid="1648" />
                    <RANKING order="37" place="37" resultid="2452" />
                    <RANKING order="38" place="38" resultid="2035" />
                    <RANKING order="39" place="39" resultid="2806" />
                    <RANKING order="40" place="40" resultid="2835" />
                    <RANKING order="41" place="41" resultid="2583" />
                    <RANKING order="42" place="42" resultid="1582" />
                    <RANKING order="43" place="43" resultid="2028" />
                    <RANKING order="44" place="44" resultid="2335" />
                    <RANKING order="45" place="45" resultid="1565" />
                    <RANKING order="46" place="46" resultid="1560" />
                    <RANKING order="47" place="47" resultid="2588" />
                    <RANKING order="48" place="48" resultid="2225" />
                    <RANKING order="49" place="49" resultid="1539" />
                    <RANKING order="50" place="50" resultid="2595" />
                    <RANKING order="51" place="51" resultid="2934" />
                    <RANKING order="52" place="52" resultid="1776" />
                    <RANKING order="53" place="-1" resultid="1886" />
                    <RANKING order="54" place="-1" resultid="1896" />
                    <RANKING order="55" place="-1" resultid="2024" />
                    <RANKING order="56" place="-1" resultid="2061" />
                    <RANKING order="57" place="-1" resultid="2089" />
                    <RANKING order="58" place="-1" resultid="2252" />
                    <RANKING order="59" place="-1" resultid="2728" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2920" daytime="11:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2921" daytime="11:27" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2922" daytime="11:33" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2923" daytime="11:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2924" daytime="11:44" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2925" daytime="11:48" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1462" gender="F" number="26" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3281" agemax="24" agemin="20" name="&quot;0&quot; 20-24" />
                <AGEGROUP agegroupid="3282" agemax="29" agemin="25" name="&quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2482" />
                    <RANKING order="2" place="2" resultid="2661" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3283" agemax="34" agemin="30" name="&quot;B&quot; 30-34" />
                <AGEGROUP agegroupid="3284" agemax="39" agemin="35" name="&quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1571" />
                    <RANKING order="2" place="2" resultid="2067" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3285" agemax="44" agemin="40" name="&quot;D&quot; 40-44" />
                <AGEGROUP agegroupid="3286" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2536" />
                    <RANKING order="2" place="2" resultid="1818" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3287" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1881" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3288" agemax="59" agemin="55" name="&quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2364" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3289" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2369" />
                    <RANKING order="2" place="2" resultid="2412" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3290" agemax="69" agemin="65" name="&quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1758" />
                    <RANKING order="2" place="2" resultid="1876" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3291" agemax="74" agemin="70" name="&quot;J&quot; 70-74" />
                <AGEGROUP agegroupid="3292" agemax="79" agemin="75" name="&quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="3293" agemax="84" agemin="80" name="&quot;L&quot; 80-84" />
                <AGEGROUP agegroupid="3294" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="3295" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2926" daytime="11:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2927" daytime="11:57" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1478" gender="M" number="27" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3296" agemax="24" agemin="20" name="&quot;0&quot; 20-24" />
                <AGEGROUP agegroupid="3297" agemax="29" agemin="25" name="&quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2487" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3298" agemax="34" agemin="30" name="&quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1796" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3299" agemax="39" agemin="35" name="&quot;C&quot; 35-39" />
                <AGEGROUP agegroupid="3300" agemax="44" agemin="40" name="&quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1813" />
                    <RANKING order="2" place="2" resultid="2796" />
                    <RANKING order="3" place="3" resultid="2736" />
                    <RANKING order="4" place="4" resultid="1763" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3301" agemax="49" agemin="45" name="&quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2443" />
                    <RANKING order="2" place="2" resultid="2072" />
                    <RANKING order="3" place="3" resultid="1801" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3302" agemax="54" agemin="50" name="&quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2320" />
                    <RANKING order="2" place="2" resultid="1808" />
                    <RANKING order="3" place="3" resultid="2492" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3303" agemax="59" agemin="55" name="&quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2217" />
                    <RANKING order="2" place="2" resultid="1786" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3304" agemax="64" agemin="60" name="&quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2630" />
                    <RANKING order="2" place="2" resultid="1969" />
                    <RANKING order="3" place="-1" resultid="2291" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3305" agemax="69" agemin="65" name="&quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2679" />
                    <RANKING order="2" place="2" resultid="1961" />
                    <RANKING order="3" place="3" resultid="2315" />
                    <RANKING order="4" place="-1" resultid="2596" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3306" agemax="74" agemin="70" name="&quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1953" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3307" agemax="79" agemin="75" name="&quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3308" agemax="84" agemin="80" name="&quot;L&quot; 80-84">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1777" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3309" agemax="89" agemin="85" name="&quot;M&quot; 85-89" />
                <AGEGROUP agegroupid="3310" agemax="94" agemin="90" name="&quot;N&quot; 90-94" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2928" daytime="12:03" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2929" daytime="12:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2930" daytime="12:17" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1494" gender="X" number="28" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3955" agemax="96" agemin="80" name="&quot;0&quot; 80-96" calculate="TOTAL" />
                <AGEGROUP agegroupid="3956" agemax="119" agemin="100" name="&quot;A&quot; 100-119" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1729" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3957" agemax="159" agemin="120" name="&quot;B&quot; 120-159" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2706" />
                    <RANKING order="2" place="2" resultid="2167" />
                    <RANKING order="3" place="3" resultid="1858" />
                    <RANKING order="4" place="4" resultid="3318" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3958" agemax="199" agemin="160" name="&quot;C&quot; 160-199" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2757" />
                    <RANKING order="2" place="2" resultid="2357" />
                    <RANKING order="3" place="3" resultid="1857" />
                    <RANKING order="4" place="4" resultid="2607" />
                    <RANKING order="5" place="5" resultid="2259" />
                    <RANKING order="6" place="6" resultid="2209" />
                    <RANKING order="7" place="7" resultid="2608" />
                    <RANKING order="8" place="-1" resultid="1898" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3959" agemax="239" agemin="200" name="&quot;D&quot; 200-239" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2609" />
                    <RANKING order="2" place="2" resultid="2415" />
                    <RANKING order="3" place="3" resultid="2707" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3960" agemax="279" agemin="240" name="&quot;E&quot; 240-279" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2358" />
                    <RANKING order="2" place="2" resultid="2610" />
                    <RANKING order="3" place="3" resultid="2416" />
                    <RANKING order="4" place="4" resultid="1980" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3961" agemax="9999" agemin="280" name="&quot;F&quot; 280 +" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1670" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3987" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3988" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3989" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" nation="POL" clubid="1616" name="Weteran Zabrze">
          <ATHLETES>
            <ATHLETE firstname="Stanisław" lastname="Twardysko" birthdate="1956-01-16" gender="M" nation="POL" license="502611700035" swrid="5464152" athleteid="1654">
              <RESULTS>
                <RESULT eventid="1076" points="123" reactiontime="+96" swimtime="00:00:44.67" resultid="1655" heatid="2842" lane="7" entrytime="00:00:45.29" entrycourse="LCM" />
                <RESULT eventid="1172" points="204" reactiontime="+93" swimtime="00:01:19.58" resultid="1656" heatid="2867" lane="8" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1382" points="173" reactiontime="+80" swimtime="00:00:42.65" resultid="1657" heatid="2909" lane="6" entrytime="00:00:42.50" />
                <RESULT eventid="1446" points="185" swimtime="00:02:58.89" resultid="1658" heatid="2924" lane="0" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.97" />
                    <SPLIT distance="100" swimtime="00:01:23.14" />
                    <SPLIT distance="150" swimtime="00:02:09.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Genowefa" lastname="Drużyńska" birthdate="1951-02-18" gender="F" nation="POL" license="102611600033" swrid="4655173" athleteid="1664">
              <RESULTS>
                <RESULT eventid="1124" points="85" swimtime="00:01:06.57" resultid="1665" heatid="2852" lane="0" entrytime="00:01:05.00" />
                <RESULT eventid="1220" points="59" swimtime="00:05:55.62" resultid="1666" heatid="2874" lane="0" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.79" />
                    <SPLIT distance="100" swimtime="00:02:51.96" />
                    <SPLIT distance="150" swimtime="00:04:24.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="72" reactiontime="+78" swimtime="00:01:04.78" resultid="1667" heatid="2905" lane="0" entrytime="00:01:05.00" />
                <RESULT eventid="1398" points="61" swimtime="00:02:42.88" resultid="1668" heatid="2911" lane="8" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Teresa" lastname="Żylińska" birthdate="1950-10-13" gender="F" nation="POL" license="102611600029" swrid="5464154" athleteid="1649">
              <RESULTS>
                <RESULT eventid="1092" points="69" reactiontime="+72" swimtime="00:02:19.65" resultid="1650" heatid="2845" lane="3" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="65" swimtime="00:02:08.30" resultid="1651" heatid="2860" lane="8" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="92" swimtime="00:00:52.36" resultid="1652" heatid="2886" lane="3" entrytime="00:00:58.00" />
                <RESULT eventid="1366" points="83" reactiontime="+76" swimtime="00:01:01.77" resultid="1653" heatid="2905" lane="2" entrytime="00:01:01.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Kosiak" birthdate="1940-04-20" gender="M" nation="POL" license="102611700027" swrid="5484411" athleteid="1644">
              <RESULTS>
                <RESULT eventid="1076" points="36" reactiontime="+112" swimtime="00:01:07.03" resultid="1645" heatid="2839" lane="5" />
                <RESULT eventid="1172" points="89" reactiontime="+113" swimtime="00:01:44.96" resultid="1646" heatid="2865" lane="4" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="103" reactiontime="+117" swimtime="00:00:44.47" resultid="1647" heatid="2893" lane="3" entrytime="00:00:44.00" />
                <RESULT eventid="1446" points="72" reactiontime="+101" swimtime="00:04:04.25" resultid="1648" heatid="2922" lane="3" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.16" />
                    <SPLIT distance="100" swimtime="00:02:04.75" />
                    <SPLIT distance="150" swimtime="00:03:08.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="9999" agetotalmin="280" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1494" reactiontime="+77" swimtime="00:03:39.06" resultid="1670" heatid="3988" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.43" />
                    <SPLIT distance="100" swimtime="00:02:08.33" />
                    <SPLIT distance="150" swimtime="00:02:53.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1649" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="1654" number="2" />
                    <RELAYPOSITION athleteid="1664" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="1644" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SIKRA" nation="POL" clubid="1566" name="Stow. Siemacha Kraków">
          <ATHLETES>
            <ATHLETE firstname="Paulina" lastname="Palmowska - Latuszek" birthdate="1985-08-01" gender="F" nation="POL" swrid="4992815" athleteid="1567">
              <RESULTS>
                <RESULT eventid="1059" points="335" reactiontime="+73" swimtime="00:00:35.16" resultid="1568" heatid="2836" lane="6" />
                <RESULT eventid="1092" points="397" reactiontime="+69" swimtime="00:01:18.11" resultid="1569" heatid="2846" lane="2" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="415" reactiontime="+72" swimtime="00:00:36.17" resultid="1570" heatid="2906" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1462" points="387" reactiontime="+72" swimtime="00:02:49.14" resultid="1571" heatid="2927" lane="3" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.03" />
                    <SPLIT distance="100" swimtime="00:01:23.18" />
                    <SPLIT distance="150" swimtime="00:02:06.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="05201" nation="POL" region="01" clubid="2260" name="KS JUST SWIM Jelenia Góra">
          <ATHLETES>
            <ATHLETE firstname="Marek" lastname="Lipka" birthdate="1958-06-05" gender="M" nation="POL" license="505201700087" swrid="5435204" athleteid="2266">
              <RESULTS>
                <RESULT eventid="1076" points="137" reactiontime="+101" swimtime="00:00:43.12" resultid="2267" heatid="2842" lane="9" />
                <RESULT eventid="1204" points="99" reactiontime="+85" swimtime="00:03:58.76" resultid="2268" heatid="2872" lane="2" entrytime="00:03:56.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.74" />
                    <SPLIT distance="100" swimtime="00:01:52.41" />
                    <SPLIT distance="150" swimtime="00:02:56.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="102" reactiontime="+82" swimtime="00:01:45.74" resultid="2269" heatid="2902" lane="3" entrytime="00:01:42.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="148" swimtime="00:03:12.72" resultid="2270" heatid="2923" lane="6" entrytime="00:03:10.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.96" />
                    <SPLIT distance="100" swimtime="00:01:35.20" />
                    <SPLIT distance="150" swimtime="00:02:27.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Lara" birthdate="1985-06-16" gender="F" nation="POL" license="505201600088" swrid="5435203" athleteid="2261">
              <RESULTS>
                <RESULT eventid="1059" points="183" reactiontime="+104" swimtime="00:00:42.97" resultid="2262" heatid="2836" lane="5" />
                <RESULT eventid="1252" points="206" reactiontime="+91" swimtime="00:03:33.33" resultid="2263" heatid="2879" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.08" />
                    <SPLIT distance="100" swimtime="00:01:48.35" />
                    <SPLIT distance="150" swimtime="00:02:46.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="155" reactiontime="+93" swimtime="00:01:43.13" resultid="2264" heatid="2899" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1430" points="257" reactiontime="+90" swimtime="00:02:57.52" resultid="2265" heatid="2918" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.10" />
                    <SPLIT distance="100" swimtime="00:01:24.81" />
                    <SPLIT distance="150" swimtime="00:02:11.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PIGUB" nation="POL" clubid="1596" name="K.S. Pionier Gubin">
          <ATHLETES>
            <ATHLETE firstname="Paweł" lastname="Krupiński" birthdate="1987-02-05" gender="M" nation="POL" athleteid="1597">
              <RESULTS>
                <RESULT eventid="1140" points="167" reactiontime="+103" swimtime="00:00:47.06" resultid="1598" heatid="2857" lane="0" entrytime="00:00:46.55" />
                <RESULT eventid="1268" points="140" swimtime="00:03:39.19" resultid="1599" heatid="2883" lane="8" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.84" />
                    <SPLIT distance="100" swimtime="00:01:44.55" />
                    <SPLIT distance="150" swimtime="00:02:40.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="135" reactiontime="+106" swimtime="00:00:40.75" resultid="1600" heatid="2893" lane="2" entrytime="00:00:46.50" />
                <RESULT eventid="1414" points="169" reactiontime="+107" swimtime="00:01:42.71" resultid="1601" heatid="2914" lane="3" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="104002" nation="POL" region="14" clubid="2822" name="Stow. AZS WSG">
          <ATHLETES>
            <ATHLETE firstname="Adrianna" lastname="Rzewuska" birthdate="1997-05-30" gender="F" nation="POL" license="504002600005" swrid="4261695" athleteid="2823">
              <RESULTS>
                <RESULT eventid="1366" status="DNS" swimtime="00:00:00.00" resultid="2824" heatid="2906" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1092" points="441" reactiontime="+73" swimtime="00:01:15.42" resultid="2825" heatid="2846" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04214" nation="POL" region="14" clubid="2637" name="Warsaw Masters Team">
          <ATHLETES>
            <ATHLETE firstname="Marcin" lastname="Giejsztowt" birthdate="1978-06-13" gender="M" nation="POL" license="504214700027" swrid="5241012" athleteid="2702">
              <RESULTS>
                <RESULT eventid="1172" points="435" reactiontime="+78" swimtime="00:01:01.88" resultid="2703" heatid="2864" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="391" reactiontime="+78" swimtime="00:02:19.41" resultid="2704" heatid="2922" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                    <SPLIT distance="100" swimtime="00:01:04.95" />
                    <SPLIT distance="150" swimtime="00:01:41.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mirosław" lastname="Warchoł" birthdate="1953-08-30" gender="M" nation="POL" license="504214700035" swrid="4222718" athleteid="2676">
              <RESULTS>
                <RESULT eventid="1108" points="230" reactiontime="+78" swimtime="00:01:24.53" resultid="2677" heatid="2847" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="285" reactiontime="+90" swimtime="00:00:31.76" resultid="2678" heatid="2896" lane="0" entrytime="00:00:31.53" entrycourse="LCM" />
                <RESULT eventid="1478" points="260" reactiontime="+110" swimtime="00:02:55.14" resultid="2679" heatid="2930" lane="1" entrytime="00:02:50.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Pfitzner" birthdate="1986-05-24" gender="M" nation="POL" license="104214700022" swrid="4992671" athleteid="2662">
              <RESULTS>
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="2663" heatid="2848" lane="0" />
                <RESULT eventid="1382" points="416" reactiontime="+84" swimtime="00:00:31.87" resultid="2664" heatid="2908" lane="3" />
                <RESULT eventid="1446" points="394" reactiontime="+80" swimtime="00:02:19.10" resultid="2665" heatid="2922" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                    <SPLIT distance="100" swimtime="00:01:08.39" />
                    <SPLIT distance="150" swimtime="00:01:45.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Rogosz" birthdate="1976-04-28" gender="M" nation="POL" license="504214700003" swrid="4270348" athleteid="2653">
              <RESULTS>
                <RESULT eventid="1076" points="313" reactiontime="+89" swimtime="00:00:32.78" resultid="2654" heatid="2841" lane="8" />
                <RESULT eventid="1268" points="355" reactiontime="+88" swimtime="00:02:40.99" resultid="2655" heatid="2881" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.53" />
                    <SPLIT distance="100" swimtime="00:01:20.44" />
                    <SPLIT distance="150" swimtime="00:02:04.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="264" reactiontime="+94" swimtime="00:01:17.04" resultid="2656" heatid="2903" lane="9" entrytime="00:01:16.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="312" reactiontime="+86" swimtime="00:02:30.24" resultid="2657" heatid="2921" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.10" />
                    <SPLIT distance="100" swimtime="00:01:15.58" />
                    <SPLIT distance="150" swimtime="00:01:54.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leszek" lastname="Madej" birthdate="1960-06-17" gender="M" nation="POL" license="504214700005" swrid="4183799" athleteid="2693">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1172" points="411" reactiontime="+83" swimtime="00:01:03.09" resultid="2694" heatid="2865" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="340" reactiontime="+86" swimtime="00:02:43.33" resultid="2695" heatid="2880" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                    <SPLIT distance="100" swimtime="00:01:17.36" />
                    <SPLIT distance="150" swimtime="00:02:06.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="379" reactiontime="+80" swimtime="00:00:28.89" resultid="2696" heatid="2890" lane="1" />
                <RESULT comment="Rekord Polski Masters" eventid="1446" points="384" reactiontime="+84" swimtime="00:02:20.26" resultid="2697" heatid="2920" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                    <SPLIT distance="100" swimtime="00:01:09.30" />
                    <SPLIT distance="150" swimtime="00:01:44.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Ostrowski" birthdate="1977-05-14" gender="M" nation="POL" license="504214700091" swrid="5506635" athleteid="2688">
              <RESULTS>
                <RESULT eventid="1140" points="517" reactiontime="+75" swimtime="00:00:32.32" resultid="2689" heatid="2855" lane="3" />
                <RESULT eventid="1236" points="403" reactiontime="+79" swimtime="00:02:50.61" resultid="2690" heatid="2876" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                    <SPLIT distance="100" swimtime="00:01:21.31" />
                    <SPLIT distance="150" swimtime="00:02:06.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="484" reactiontime="+75" swimtime="00:00:26.62" resultid="2691" heatid="2892" lane="8" />
                <RESULT eventid="1414" points="464" reactiontime="+78" swimtime="00:01:13.46" resultid="2692" heatid="2913" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robert" lastname="Sutowski" birthdate="1959-12-03" gender="M" nation="POL" license="104214700079" swrid="4992657" athleteid="2643">
              <RESULTS>
                <RESULT eventid="1076" points="75" reactiontime="+100" swimtime="00:00:52.80" resultid="2644" heatid="2840" lane="3" />
                <RESULT eventid="1172" points="147" reactiontime="+104" swimtime="00:01:28.78" resultid="2645" heatid="2863" lane="6" />
                <RESULT eventid="1318" points="139" reactiontime="+101" swimtime="00:00:40.27" resultid="2646" heatid="2890" lane="6" />
                <RESULT eventid="1446" points="152" reactiontime="+106" swimtime="00:03:10.95" resultid="2647" heatid="2920" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.98" />
                    <SPLIT distance="100" swimtime="00:01:32.41" />
                    <SPLIT distance="150" swimtime="00:02:23.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Kośla" birthdate="1993-01-05" gender="F" nation="POL" license="104214600085" swrid="4086961" athleteid="2658">
              <RESULTS>
                <RESULT eventid="1092" points="421" reactiontime="+78" swimtime="00:01:16.64" resultid="2659" heatid="2846" lane="4" entrytime="00:01:09.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="497" reactiontime="+82" swimtime="00:00:34.05" resultid="2660" heatid="2906" lane="5" entrytime="00:00:32.52" entrycourse="LCM" />
                <RESULT eventid="1462" points="365" reactiontime="+83" swimtime="00:02:52.47" resultid="2661" heatid="2927" lane="4" entrytime="00:02:38.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                    <SPLIT distance="100" swimtime="00:01:24.68" />
                    <SPLIT distance="150" swimtime="00:02:09.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Szemberg" birthdate="1949-07-26" gender="F" nation="POL" license="504214600017" swrid="4302692" athleteid="2680">
              <RESULTS>
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="2681" heatid="2851" lane="6" />
                <RESULT eventid="1430" points="69" swimtime="00:04:34.36" resultid="2682" heatid="2918" lane="7" entrytime="00:04:39.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.27" />
                    <SPLIT distance="100" swimtime="00:02:13.01" />
                    <SPLIT distance="150" swimtime="00:03:24.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Skośkiewicz" birthdate="1966-05-05" gender="M" nation="POL" license="504214700002" swrid="4183802" athleteid="2666">
              <RESULTS>
                <RESULT eventid="1108" points="355" reactiontime="+78" swimtime="00:01:13.18" resultid="2667" heatid="2850" lane="7" entrytime="00:01:12.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="368" reactiontime="+80" swimtime="00:02:38.96" resultid="2668" heatid="2881" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                    <SPLIT distance="100" swimtime="00:01:15.90" />
                    <SPLIT distance="150" swimtime="00:02:02.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1382" points="360" reactiontime="+80" swimtime="00:00:33.45" resultid="2669" heatid="2910" lane="7" entrytime="00:00:33.54" entrycourse="LCM" />
                <RESULT eventid="1446" points="392" reactiontime="+87" swimtime="00:02:19.30" resultid="2670" heatid="2920" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                    <SPLIT distance="100" swimtime="00:01:08.29" />
                    <SPLIT distance="150" swimtime="00:01:43.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katharina" lastname="Szymańska" birthdate="1985-05-31" gender="F" nation="POL" license="504214600036" swrid="5312493" athleteid="2683">
              <RESULTS>
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="2684" heatid="2851" lane="3" />
                <RESULT eventid="1252" status="DNS" swimtime="00:00:00.00" resultid="2685" heatid="2879" lane="0" />
                <RESULT eventid="1366" points="159" reactiontime="+81" swimtime="00:00:49.80" resultid="2686" heatid="2904" lane="4" />
                <RESULT eventid="1430" points="174" reactiontime="+100" swimtime="00:03:22.35" resultid="2687" heatid="2918" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.05" />
                    <SPLIT distance="100" swimtime="00:01:37.24" />
                    <SPLIT distance="150" swimtime="00:02:31.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Porada" birthdate="1983-06-10" gender="M" nation="POL" license="104214700058" swrid="5506638" athleteid="2648">
              <RESULTS>
                <RESULT eventid="1076" points="411" reactiontime="+74" swimtime="00:00:29.95" resultid="2649" heatid="2841" lane="7" />
                <RESULT eventid="1236" points="428" reactiontime="+78" swimtime="00:02:47.27" resultid="2650" heatid="2876" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                    <SPLIT distance="100" swimtime="00:01:19.47" />
                    <SPLIT distance="150" swimtime="00:02:02.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="408" reactiontime="+70" swimtime="00:00:28.18" resultid="2651" heatid="2891" lane="0" />
                <RESULT eventid="1414" points="418" reactiontime="+73" swimtime="00:01:16.04" resultid="2652" heatid="2913" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Burdelak" birthdate="1991-07-06" gender="F" nation="POL" license="504214600100" swrid="4072596" athleteid="2638">
              <RESULTS>
                <RESULT eventid="1059" points="453" reactiontime="+68" swimtime="00:00:31.80" resultid="2639" heatid="2838" lane="7" entrytime="00:00:32.37" entrycourse="LCM" />
                <RESULT eventid="1124" points="476" reactiontime="+79" swimtime="00:00:37.52" resultid="2640" heatid="2853" lane="5" entrytime="00:00:36.48" entrycourse="LCM" />
                <RESULT eventid="1301" points="507" reactiontime="+71" swimtime="00:00:29.67" resultid="2641" heatid="2889" lane="7" entrytime="00:00:29.18" entrycourse="LCM" />
                <RESULT eventid="1398" points="416" reactiontime="+71" swimtime="00:01:25.87" resultid="2642" heatid="2912" lane="3" entrytime="00:01:24.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Szymański" birthdate="1980-10-04" gender="M" nation="POL" license="504214700028" swrid="4542528" athleteid="2671">
              <RESULTS>
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="2672" heatid="2848" lane="8" />
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="2673" heatid="2881" lane="8" />
                <RESULT eventid="1318" points="514" reactiontime="+70" swimtime="00:00:26.09" resultid="2674" heatid="2891" lane="2" />
                <RESULT eventid="1382" points="527" reactiontime="+69" swimtime="00:00:29.46" resultid="2675" heatid="2907" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Waldemar" lastname="De Makay" birthdate="1950-10-17" gender="M" nation="POL" license="504214700148" athleteid="2698">
              <RESULTS>
                <RESULT eventid="1172" status="DNS" swimtime="00:00:00.00" resultid="2699" heatid="2863" lane="2" />
                <RESULT eventid="1318" points="162" reactiontime="+111" swimtime="00:00:38.34" resultid="2700" heatid="2890" lane="2" />
                <RESULT eventid="1446" points="164" reactiontime="+129" swimtime="00:03:06.00" resultid="2701" heatid="2920" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.14" />
                    <SPLIT distance="100" swimtime="00:01:30.29" />
                    <SPLIT distance="150" swimtime="00:02:18.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1284" reactiontime="+73" swimtime="00:01:52.10" resultid="2705" heatid="3970" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.16" />
                    <SPLIT distance="100" swimtime="00:00:52.94" />
                    <SPLIT distance="150" swimtime="00:01:23.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2671" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="2688" number="2" />
                    <RELAYPOSITION athleteid="2658" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="2638" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1494" reactiontime="+89" swimtime="00:02:06.77" resultid="2706" heatid="3989" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                    <SPLIT distance="100" swimtime="00:01:07.90" />
                    <SPLIT distance="150" swimtime="00:01:40.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2658" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="2648" number="2" />
                    <RELAYPOSITION athleteid="2638" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="2662" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1494" reactiontime="+77" swimtime="00:03:09.79" resultid="2707" heatid="3987" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                    <SPLIT distance="100" swimtime="00:01:24.73" />
                    <SPLIT distance="150" swimtime="00:02:11.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2666" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="2676" number="2" />
                    <RELAYPOSITION athleteid="2683" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="2680" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="1991" name="3Waters">
          <ATHLETES>
            <ATHLETE firstname="Sonia" lastname="Borkowska" birthdate="1975-08-09" gender="F" nation="POL" athleteid="1990">
              <RESULTS>
                <RESULT eventid="1301" points="361" reactiontime="+79" swimtime="00:00:33.22" resultid="1992" heatid="2888" lane="0" entrytime="00:00:36.00" />
                <RESULT eventid="1366" points="210" reactiontime="+103" swimtime="00:00:45.39" resultid="1993" heatid="2906" lane="9" entrytime="00:00:46.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="100111" nation="POL" clubid="1671" name="UKS TRÓJKA Częstochowa">
          <ATHLETES>
            <ATHLETE firstname="Mateusz" lastname="Kurek" birthdate="1994-07-11" gender="M" nation="POL" license="100111700097" swrid="5502059" athleteid="1708">
              <RESULTS>
                <RESULT eventid="1076" points="323" reactiontime="+68" swimtime="00:00:32.44" resultid="1709" heatid="2843" lane="4" entrytime="00:00:29.97" />
                <RESULT eventid="1172" points="415" reactiontime="+70" swimtime="00:01:02.87" resultid="1710" heatid="2868" lane="6" entrytime="00:01:03.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="405" reactiontime="+67" swimtime="00:00:28.25" resultid="1711" heatid="2897" lane="9" entrytime="00:00:28.34" />
                <RESULT eventid="1446" points="329" reactiontime="+67" swimtime="00:02:27.68" resultid="1712" heatid="2925" lane="0" entrytime="00:02:29.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.19" />
                    <SPLIT distance="100" swimtime="00:01:08.59" />
                    <SPLIT distance="150" swimtime="00:01:48.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Gajda" birthdate="1995-04-23" gender="M" nation="POL" license="100111700062" swrid="4762175" athleteid="1703">
              <RESULTS>
                <RESULT eventid="1076" points="591" reactiontime="+76" swimtime="00:00:26.53" resultid="1704" heatid="2844" lane="5" entrytime="00:00:26.92" />
                <RESULT eventid="1172" points="587" reactiontime="+73" swimtime="00:00:56.01" resultid="1705" heatid="2869" lane="3" entrytime="00:00:55.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="586" reactiontime="+71" swimtime="00:00:24.98" resultid="1706" heatid="2898" lane="5" entrytime="00:00:25.04" />
                <RESULT eventid="1350" points="530" reactiontime="+71" swimtime="00:01:01.09" resultid="1707" heatid="2903" lane="5" entrytime="00:01:00.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sonia" lastname="Nowak" birthdate="1996-05-23" gender="F" nation="POL" license="100111600092" swrid="4289072" athleteid="1713">
              <RESULTS>
                <RESULT eventid="1059" points="379" reactiontime="+88" swimtime="00:00:33.73" resultid="1714" heatid="2838" lane="1" entrytime="00:00:33.80" />
                <RESULT eventid="1156" points="447" reactiontime="+89" swimtime="00:01:07.59" resultid="1715" heatid="2862" lane="7" entrytime="00:01:08.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="397" reactiontime="+93" swimtime="00:00:32.20" resultid="1716" heatid="2889" lane="8" entrytime="00:00:32.00" />
                <RESULT eventid="1430" points="411" reactiontime="+87" swimtime="00:02:31.91" resultid="1717" heatid="2919" lane="2" entrytime="00:02:31.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.87" />
                    <SPLIT distance="100" swimtime="00:01:12.87" />
                    <SPLIT distance="150" swimtime="00:01:52.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Musik" birthdate="1997-08-04" gender="F" nation="POL" license="100111600053" swrid="4602697" athleteid="1718">
              <RESULTS>
                <RESULT eventid="1059" points="530" reactiontime="+79" swimtime="00:00:30.17" resultid="1719" heatid="2838" lane="5" entrytime="00:00:30.83" />
                <RESULT eventid="1156" points="622" reactiontime="+80" swimtime="00:01:00.55" resultid="1720" heatid="2862" lane="4" entrytime="00:01:00.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="639" reactiontime="+78" swimtime="00:00:27.48" resultid="1721" heatid="2889" lane="4" entrytime="00:00:27.29" />
                <RESULT eventid="1430" points="546" reactiontime="+80" swimtime="00:02:18.20" resultid="1722" heatid="2919" lane="4" entrytime="00:02:12.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.92" />
                    <SPLIT distance="100" swimtime="00:01:04.85" />
                    <SPLIT distance="150" swimtime="00:01:42.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1284" reactiontime="+67" swimtime="00:01:49.94" resultid="1697" heatid="3970" lane="4" entrytime="00:02:07.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.71" />
                    <SPLIT distance="100" swimtime="00:00:58.86" />
                    <SPLIT distance="150" swimtime="00:01:25.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1708" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="1713" number="2" />
                    <RELAYPOSITION athleteid="1718" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="1703" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1494" reactiontime="+78" swimtime="00:02:07.23" resultid="1729" heatid="3989" lane="4" entrytime="00:02:07.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                    <SPLIT distance="100" swimtime="00:01:10.20" />
                    <SPLIT distance="150" swimtime="00:00:50.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1718" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="1708" number="2" />
                    <RELAYPOSITION athleteid="1703" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="1713" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00501" nation="POL" clubid="1910" name="UKS Energetyk Zgorzelec" />
        <CLUB type="CLUB" code="03415" nation="POL" clubid="1930" name="UKS Cityzen">
          <ATHLETES>
            <ATHLETE firstname="Teresa" lastname="Barełkowska" birthdate="1948-01-01" gender="F" nation="POL" swrid="4920301" athleteid="1931">
              <RESULTS>
                <RESULT eventid="1092" points="33" reactiontime="+94" swimtime="00:02:57.71" resultid="1932" heatid="2845" lane="5" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="70" swimtime="00:01:10.76" resultid="1933" heatid="2852" lane="8" entrytime="00:01:00.00" />
                <RESULT eventid="1366" points="45" swimtime="00:01:15.52" resultid="1934" heatid="2905" lane="6" entrytime="00:01:00.00" />
                <RESULT eventid="1398" points="65" swimtime="00:02:39.22" resultid="1935" heatid="2911" lane="2" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sławomir" lastname="Cybertowicz" birthdate="1966-01-01" gender="M" nation="POL" swrid="4269915" athleteid="1970">
              <RESULTS>
                <RESULT eventid="1076" points="214" reactiontime="+87" swimtime="00:00:37.23" resultid="1971" heatid="2842" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="1140" points="300" reactiontime="+84" swimtime="00:00:38.75" resultid="1972" heatid="2857" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="1414" points="265" reactiontime="+85" swimtime="00:01:28.52" resultid="1973" heatid="2915" lane="7" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Boryski" birthdate="1951-01-01" gender="M" nation="POL" swrid="4754708" athleteid="1950">
              <RESULTS>
                <RESULT eventid="1108" points="116" reactiontime="+93" swimtime="00:01:46.05" resultid="1951" heatid="2849" lane="1" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1382" points="137" reactiontime="+82" swimtime="00:00:46.08" resultid="1952" heatid="2909" lane="1" entrytime="00:00:45.00" />
                <RESULT eventid="1478" points="103" reactiontime="+98" swimtime="00:03:58.32" resultid="1953" heatid="2929" lane="2" entrytime="00:03:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.95" />
                    <SPLIT distance="100" swimtime="00:02:00.59" />
                    <SPLIT distance="150" swimtime="00:03:01.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Łutowicz" birthdate="1950-01-01" gender="F" nation="POL" swrid="4188428" athleteid="1936">
              <RESULTS>
                <RESULT eventid="1156" points="95" swimtime="00:01:53.27" resultid="1937" heatid="2860" lane="7" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="104" swimtime="00:00:50.24" resultid="1938" heatid="2887" lane="9" entrytime="00:00:53.00" />
                <RESULT eventid="1366" points="96" swimtime="00:00:58.92" resultid="1939" heatid="2905" lane="8" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Łasińska" birthdate="1954-01-01" gender="F" nation="POL" athleteid="1940">
              <RESULTS>
                <RESULT eventid="1059" points="69" reactiontime="+117" swimtime="00:00:59.44" resultid="1941" heatid="2837" lane="9" entrytime="00:01:00.00" />
                <RESULT eventid="1124" points="123" reactiontime="+108" swimtime="00:00:58.85" resultid="1942" heatid="2852" lane="1" entrytime="00:01:00.00" />
                <RESULT eventid="1301" points="97" reactiontime="+90" swimtime="00:00:51.36" resultid="1943" heatid="2887" lane="0" entrytime="00:00:50.00" />
                <RESULT eventid="1366" points="93" reactiontime="+90" swimtime="00:00:59.51" resultid="1944" heatid="2905" lane="3" entrytime="00:00:56.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Matyszczak" birthdate="1970-01-01" gender="M" nation="POL" swrid="5471729" athleteid="1974">
              <RESULTS>
                <RESULT eventid="1172" points="249" reactiontime="+89" swimtime="00:01:14.49" resultid="1975" heatid="2867" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="160" reactiontime="+101" swimtime="00:03:51.99" resultid="1976" heatid="2877" lane="0" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.97" />
                    <SPLIT distance="100" swimtime="00:01:47.79" />
                    <SPLIT distance="150" swimtime="00:02:48.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="299" reactiontime="+112" swimtime="00:00:31.25" resultid="1977" heatid="2896" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="1446" points="198" reactiontime="+105" swimtime="00:02:54.80" resultid="1978" heatid="2924" lane="1" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:08.10" />
                    <SPLIT distance="100" swimtime="00:01:21.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zbigniew" lastname="Pietraszewski" birthdate="1955-01-01" gender="M" nation="POL" swrid="4187282" athleteid="1957">
              <RESULTS>
                <RESULT eventid="1108" points="150" reactiontime="+94" swimtime="00:01:37.58" resultid="1958" heatid="2849" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="168" reactiontime="+96" swimtime="00:03:26.58" resultid="1959" heatid="2883" lane="1" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.80" />
                    <SPLIT distance="100" swimtime="00:01:44.01" />
                    <SPLIT distance="150" swimtime="00:02:40.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1382" points="140" reactiontime="+89" swimtime="00:00:45.73" resultid="1960" heatid="2909" lane="7" entrytime="00:00:44.00" />
                <RESULT eventid="1478" points="160" reactiontime="+88" swimtime="00:03:25.77" resultid="1961" heatid="2929" lane="4" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.47" />
                    <SPLIT distance="100" swimtime="00:01:41.84" />
                    <SPLIT distance="150" swimtime="00:02:34.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Nochowicz" birthdate="1951-01-01" gender="M" nation="POL" swrid="5471731" athleteid="1954">
              <RESULTS>
                <RESULT eventid="1108" points="69" reactiontime="+97" swimtime="00:02:06.08" resultid="1955" heatid="2848" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1382" points="68" reactiontime="+87" swimtime="00:00:58.13" resultid="1956" heatid="2908" lane="5" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Szczesiak" birthdate="1955-01-01" gender="M" nation="POL" athleteid="1962">
              <RESULTS>
                <RESULT eventid="1172" status="DNS" swimtime="00:00:00.00" resultid="1963" heatid="2867" lane="0" entrytime="00:01:20.00" />
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="1964" heatid="2894" lane="5" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jarosław" lastname="Miśkiewicz" birthdate="1959-01-01" gender="M" nation="POL" swrid="4920302" athleteid="1965">
              <RESULTS>
                <RESULT eventid="1108" points="109" reactiontime="+96" swimtime="00:01:48.53" resultid="1966" heatid="2849" lane="8" entrytime="00:01:46.00" />
                <RESULT eventid="1268" points="73" reactiontime="+112" swimtime="00:04:31.70" resultid="1967" heatid="2882" lane="5" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.86" />
                    <SPLIT distance="100" swimtime="00:02:05.96" />
                    <SPLIT distance="150" swimtime="00:03:26.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1382" points="124" reactiontime="+101" swimtime="00:00:47.67" resultid="1968" heatid="2909" lane="8" entrytime="00:00:50.00" />
                <RESULT eventid="1478" points="99" reactiontime="+101" swimtime="00:04:01.88" resultid="1969" heatid="2929" lane="6" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.49" />
                    <SPLIT distance="100" swimtime="00:01:56.90" />
                    <SPLIT distance="150" swimtime="00:03:00.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dorota" lastname="Masłek" birthdate="1953-01-01" gender="F" nation="POL" athleteid="1945">
              <RESULTS>
                <RESULT eventid="1124" points="122" reactiontime="+104" swimtime="00:00:58.99" resultid="1946" heatid="2852" lane="3" entrytime="00:00:50.00" />
                <RESULT eventid="1220" points="114" reactiontime="+97" swimtime="00:04:45.90" resultid="1947" heatid="2874" lane="6" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.25" />
                    <SPLIT distance="100" swimtime="00:02:16.55" />
                    <SPLIT distance="150" swimtime="00:03:31.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="104" reactiontime="+98" swimtime="00:00:50.24" resultid="1948" heatid="2887" lane="2" entrytime="00:00:45.00" />
                <RESULT eventid="1398" points="116" reactiontime="+96" swimtime="00:02:11.13" resultid="1949" heatid="2911" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="9999" agetotalmin="280" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1284" reactiontime="+101" swimtime="00:03:24.23" resultid="1979" heatid="3969" lane="0" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                    <SPLIT distance="100" swimtime="00:01:56.90" />
                    <SPLIT distance="150" swimtime="00:02:47.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1950" number="1" reactiontime="+101" />
                    <RELAYPOSITION athleteid="1931" number="2" />
                    <RELAYPOSITION athleteid="1945" number="3" />
                    <RELAYPOSITION athleteid="1957" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1494" reactiontime="+102" swimtime="00:03:07.34" resultid="1980" heatid="3988" lane="6" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.50" />
                    <SPLIT distance="100" swimtime="00:02:04.10" />
                    <SPLIT distance="150" swimtime="00:02:37.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1940" number="1" reactiontime="+102" />
                    <RELAYPOSITION athleteid="1945" number="2" />
                    <RELAYPOSITION athleteid="1970" number="3" />
                    <RELAYPOSITION athleteid="1974" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="1735" name="MOSiR Ostrowiec Św.">
          <ATHLETES>
            <ATHLETE firstname="Józef" lastname="Różalski" birthdate="1945-03-28" gender="M" nation="POL" license="501012700001" swrid="4216999" athleteid="1736">
              <RESULTS>
                <RESULT eventid="1108" points="78" reactiontime="+100" swimtime="00:02:01.01" resultid="1737" heatid="2848" lane="6" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="104" swimtime="00:00:55.05" resultid="1738" heatid="2856" lane="5" entrytime="00:00:50.00" />
                <RESULT eventid="1414" points="70" reactiontime="+102" swimtime="00:02:17.37" resultid="1739" heatid="2914" lane="2" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1382" points="99" reactiontime="+80" swimtime="00:00:51.33" resultid="1740" heatid="2908" lane="4" entrytime="00:00:52.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="1802" name="MKS Astoria Masters">
          <ATHLETES>
            <ATHLETE firstname="Wiktor" lastname="Michalski" birthdate="1982-02-13" gender="M" nation="POL" athleteid="1759">
              <RESULTS>
                <RESULT eventid="1172" points="290" reactiontime="+101" swimtime="00:01:10.87" resultid="1760" heatid="2868" lane="7" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="277" reactiontime="+88" swimtime="00:01:19.50" resultid="1761" heatid="2849" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1382" points="287" reactiontime="+72" swimtime="00:00:36.04" resultid="1762" heatid="2910" lane="0" entrytime="00:00:36.00" />
                <RESULT eventid="1478" points="211" reactiontime="+115" swimtime="00:03:07.79" resultid="1763" heatid="2930" lane="0" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.74" />
                    <SPLIT distance="100" swimtime="00:01:29.85" />
                    <SPLIT distance="150" swimtime="00:02:18.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="05" clubid="1809" name="MASTERS Łódź">
          <ATHLETES>
            <ATHLETE firstname="Michał" lastname="Woźniak" birthdate="1981-08-25" gender="M" nation="POL" license="503605700034" swrid="5484423" athleteid="1810">
              <RESULTS>
                <RESULT eventid="1108" points="443" reactiontime="+61" swimtime="00:01:07.99" resultid="1811" heatid="2850" lane="5" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1382" points="453" reactiontime="+53" swimtime="00:00:30.98" resultid="1812" heatid="2910" lane="4" entrytime="00:00:29.50" />
                <RESULT eventid="1478" points="355" reactiontime="+70" swimtime="00:02:38.02" resultid="1813" heatid="2930" lane="4" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                    <SPLIT distance="100" swimtime="00:01:18.51" />
                    <SPLIT distance="150" swimtime="00:01:58.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Lipka" birthdate="1980-12-18" gender="M" nation="POL" license="503605700025" athleteid="2073">
              <RESULTS>
                <RESULT eventid="1076" points="186" reactiontime="+90" swimtime="00:00:38.96" resultid="2074" heatid="2841" lane="1" />
                <RESULT eventid="1268" points="164" reactiontime="+97" swimtime="00:03:28.13" resultid="2075" heatid="2881" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.84" />
                    <SPLIT distance="100" swimtime="00:01:41.00" />
                    <SPLIT distance="150" swimtime="00:02:39.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="231" reactiontime="+91" swimtime="00:00:34.07" resultid="2076" heatid="2892" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewa" lastname="Adamska" birthdate="1984-09-25" gender="F" nation="POL" license="503605600036" swrid="5464086" athleteid="1829">
              <RESULTS>
                <RESULT eventid="1059" points="225" reactiontime="+88" swimtime="00:00:40.15" resultid="1830" heatid="2837" lane="6" entrytime="00:00:39.00" />
                <RESULT eventid="1156" points="304" reactiontime="+80" swimtime="00:01:16.83" resultid="1831" heatid="2861" lane="9" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="193" reactiontime="+83" swimtime="00:01:35.91" resultid="1832" heatid="2900" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1430" points="243" reactiontime="+85" swimtime="00:03:00.88" resultid="1833" heatid="2918" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.38" />
                    <SPLIT distance="150" swimtime="00:02:15.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Kruszyna-Kotulski" birthdate="1979-05-25" gender="M" nation="POL" license="503605700044" athleteid="1850">
              <RESULTS>
                <RESULT eventid="1076" points="371" reactiontime="+80" swimtime="00:00:30.98" resultid="1851" heatid="2843" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1140" points="248" reactiontime="+71" swimtime="00:00:41.25" resultid="1852" heatid="2857" lane="3" entrytime="00:00:41.00" />
                <RESULT eventid="1318" points="359" reactiontime="+72" swimtime="00:00:29.40" resultid="1853" heatid="2897" lane="1" entrytime="00:00:28.00" />
                <RESULT eventid="1382" points="226" reactiontime="+85" swimtime="00:00:39.04" resultid="1854" heatid="2909" lane="5" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Michniewski" birthdate="1983-04-11" gender="M" nation="POL" license="503605700012" athleteid="1845">
              <RESULTS>
                <RESULT eventid="1140" points="403" reactiontime="+80" swimtime="00:00:35.13" resultid="1846" heatid="2858" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1236" points="366" reactiontime="+87" swimtime="00:02:56.30" resultid="1847" heatid="2877" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                    <SPLIT distance="100" swimtime="00:01:21.29" />
                    <SPLIT distance="150" swimtime="00:02:09.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="418" reactiontime="+79" swimtime="00:00:27.96" resultid="1848" heatid="2898" lane="9" entrytime="00:00:27.00" />
                <RESULT eventid="1414" points="394" reactiontime="+79" swimtime="00:01:17.55" resultid="1849" heatid="2916" lane="0" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Olejarczyk" birthdate="1979-06-12" gender="M" nation="POL" license="503605700007" swrid="4992959" athleteid="1819">
              <RESULTS>
                <RESULT eventid="1076" points="418" reactiontime="+81" swimtime="00:00:29.78" resultid="1820" heatid="2843" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1172" points="450" reactiontime="+88" swimtime="00:01:01.18" resultid="1821" heatid="2868" lane="4" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="437" reactiontime="+81" swimtime="00:00:27.55" resultid="1822" heatid="2897" lane="4" entrytime="00:00:27.00" />
                <RESULT eventid="1350" points="338" reactiontime="+83" swimtime="00:01:10.93" resultid="1823" heatid="2903" lane="7" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Magdalena" lastname="Maciąg" birthdate="1987-03-12" gender="F" nation="POL" license="503605600031" swrid="5484414" athleteid="1824">
              <RESULTS>
                <RESULT eventid="1059" points="308" reactiontime="+81" swimtime="00:00:36.14" resultid="1825" heatid="2837" lane="3" entrytime="00:00:38.00" />
                <RESULT eventid="1156" points="328" reactiontime="+84" swimtime="00:01:14.94" resultid="1826" heatid="2861" lane="4" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="346" reactiontime="+89" swimtime="00:00:33.70" resultid="1827" heatid="2888" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1430" points="290" reactiontime="+91" swimtime="00:02:50.66" resultid="1828" heatid="2919" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.59" />
                    <SPLIT distance="100" swimtime="00:01:22.67" />
                    <SPLIT distance="150" swimtime="00:02:06.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Klarecka" birthdate="1977-06-06" gender="F" nation="POL" license="503605600029" swrid="5464091" athleteid="1814">
              <RESULTS>
                <RESULT eventid="1188" points="141" reactiontime="+110" swimtime="00:03:53.62" resultid="1815" heatid="2870" lane="3" entrytime="00:03:46.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.85" />
                    <SPLIT distance="100" swimtime="00:01:52.86" />
                    <SPLIT distance="150" swimtime="00:02:54.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1220" points="200" reactiontime="+114" swimtime="00:03:57.31" resultid="1816" heatid="2874" lane="3" entrytime="00:03:47.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.39" />
                    <SPLIT distance="100" swimtime="00:01:57.05" />
                    <SPLIT distance="150" swimtime="00:02:57.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1430" points="180" reactiontime="+117" swimtime="00:03:20.07" resultid="1817" heatid="2918" lane="5" entrytime="00:03:13.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.00" />
                    <SPLIT distance="100" swimtime="00:01:36.60" />
                    <SPLIT distance="150" swimtime="00:02:29.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="104" swimtime="00:04:21.53" resultid="1818" heatid="2927" lane="8" entrytime="00:04:08.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.36" />
                    <SPLIT distance="100" swimtime="00:02:11.15" />
                    <SPLIT distance="150" swimtime="00:03:18.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Kurstak-Jagiełło" birthdate="1981-06-30" gender="F" nation="POL" license="503605600022" athleteid="1834">
              <RESULTS>
                <RESULT eventid="1156" points="441" reactiontime="+90" swimtime="00:01:07.91" resultid="1835" heatid="2860" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="459" reactiontime="+80" swimtime="00:00:30.68" resultid="1836" heatid="2886" lane="2" />
                <RESULT eventid="1430" points="381" reactiontime="+83" swimtime="00:02:35.75" resultid="1837" heatid="2917" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.46" />
                    <SPLIT distance="100" swimtime="00:01:14.07" />
                    <SPLIT distance="150" swimtime="00:01:55.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artur" lastname="Frąckowiak" birthdate="1978-06-28" gender="M" nation="POL" license="503605700020" swrid="5279744" athleteid="1841">
              <RESULTS>
                <RESULT eventid="1076" points="372" reactiontime="+88" swimtime="00:00:30.96" resultid="1842" heatid="2841" lane="0" />
                <RESULT eventid="1172" points="355" reactiontime="+88" swimtime="00:01:06.25" resultid="1843" heatid="2865" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="389" reactiontime="+81" swimtime="00:00:28.63" resultid="1844" heatid="2891" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Babuchowski" birthdate="1984-06-08" gender="M" nation="POL" license="503605700040" swrid="4037687" athleteid="2077">
              <RESULTS>
                <RESULT eventid="1076" points="603" reactiontime="+75" swimtime="00:00:26.36" resultid="2078" heatid="2841" lane="4" />
                <RESULT eventid="1172" points="551" reactiontime="+72" swimtime="00:00:57.19" resultid="2079" heatid="2865" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="478" reactiontime="+74" swimtime="00:01:03.21" resultid="2080" heatid="2902" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Gurbski" birthdate="1976-06-09" gender="M" nation="POL" license="503605700026" athleteid="1838">
              <RESULTS>
                <RESULT eventid="1318" points="272" reactiontime="+90" swimtime="00:00:32.25" resultid="1839" heatid="2891" lane="3" />
                <RESULT eventid="1382" points="252" reactiontime="+87" swimtime="00:00:37.67" resultid="1840" heatid="2908" lane="9" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1494" reactiontime="+65" swimtime="00:02:20.37" resultid="1857" heatid="3989" lane="5" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                    <SPLIT distance="100" swimtime="00:01:21.38" />
                    <SPLIT distance="150" swimtime="00:01:50.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1810" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="1814" number="2" />
                    <RELAYPOSITION athleteid="1819" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="1834" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1284" reactiontime="+91" swimtime="00:01:59.42" resultid="2081" heatid="3970" lane="9" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                    <SPLIT distance="100" swimtime="00:00:58.17" />
                    <SPLIT distance="150" swimtime="00:01:32.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1834" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="1810" number="2" />
                    <RELAYPOSITION athleteid="1824" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="1819" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1284" reactiontime="+75" swimtime="00:02:10.44" resultid="1856" heatid="3970" lane="2" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.54" />
                    <SPLIT distance="100" swimtime="00:01:02.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1841" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="1829" number="2" />
                    <RELAYPOSITION athleteid="1814" number="3" reactiontime="+70" />
                    <RELAYPOSITION athleteid="1845" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1494" reactiontime="+90" swimtime="00:02:20.34" resultid="1858" heatid="3989" lane="9" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.29" />
                    <SPLIT distance="100" swimtime="00:01:15.94" />
                    <SPLIT distance="150" swimtime="00:01:46.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1829" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="1845" number="2" />
                    <RELAYPOSITION athleteid="1841" number="3" reactiontime="+67" />
                    <RELAYPOSITION athleteid="1824" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="TMT" nation="POL" clubid="1866" name="Toruń Multisport Team">
          <ATHLETES>
            <ATHLETE firstname="Lucyna" lastname="Serożyńska" birthdate="1955-06-29" gender="F" nation="POL" swrid="5469132" athleteid="1872">
              <RESULTS>
                <RESULT eventid="1092" points="82" reactiontime="+94" swimtime="00:02:11.83" resultid="1873" heatid="2845" lane="6" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="85" reactiontime="+127" swimtime="00:01:57.47" resultid="1874" heatid="2860" lane="2" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="82" reactiontime="+118" swimtime="00:00:54.27" resultid="1875" heatid="2886" lane="4" entrytime="00:00:55.70" />
                <RESULT eventid="1462" points="75" reactiontime="+111" swimtime="00:04:51.76" resultid="1876" heatid="2926" lane="4" entrytime="00:04:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.00" />
                    <SPLIT distance="150" swimtime="00:03:41.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kamil" lastname="Kordowski" birthdate="1997-10-11" gender="M" nation="POL" swrid="5506630" athleteid="1867">
              <RESULTS>
                <RESULT eventid="1076" points="444" reactiontime="+73" swimtime="00:00:29.19" resultid="1868" heatid="2843" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1172" points="439" reactiontime="+75" swimtime="00:01:01.71" resultid="1869" heatid="2869" lane="0" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="432" reactiontime="+84" swimtime="00:00:27.64" resultid="1870" heatid="2892" lane="6" />
                <RESULT eventid="1350" points="351" reactiontime="+77" swimtime="00:01:10.06" resultid="1871" heatid="2903" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Marchewka" birthdate="1981-02-04" gender="M" nation="POL" swrid="5506633" athleteid="1887">
              <RESULTS>
                <RESULT eventid="1108" points="393" reactiontime="+77" swimtime="00:01:10.75" resultid="1888" heatid="2850" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="1889" heatid="2883" lane="3" entrytime="00:02:40.00" />
                <RESULT eventid="1382" points="428" reactiontime="+68" swimtime="00:00:31.56" resultid="1890" heatid="2908" lane="1" />
                <RESULT eventid="1414" status="DNS" swimtime="00:00:00.00" resultid="1891" heatid="2916" lane="9" entrytime="00:01:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artur" lastname="Rybicki" birthdate="1984-01-15" gender="M" nation="POL" swrid="5506640" athleteid="1892">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="1893" heatid="2843" lane="8" entrytime="00:00:32.00" />
                <RESULT eventid="1172" status="DNS" swimtime="00:00:00.00" resultid="1894" heatid="2868" lane="3" entrytime="00:01:03.00" />
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="1895" heatid="2897" lane="2" entrytime="00:00:28.00" />
                <RESULT eventid="1446" status="DNS" swimtime="00:00:00.00" resultid="1896" heatid="2925" lane="9" entrytime="00:02:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Arentewicz" birthdate="1981-03-07" gender="M" nation="POL" swrid="4754686" athleteid="1882">
              <RESULTS>
                <RESULT eventid="1076" points="302" reactiontime="+79" swimtime="00:00:33.17" resultid="1883" heatid="2843" lane="9" entrytime="00:00:34.00" />
                <RESULT eventid="1172" points="272" reactiontime="+78" swimtime="00:01:12.36" resultid="1884" heatid="2867" lane="3" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="281" reactiontime="+85" swimtime="00:00:31.91" resultid="1885" heatid="2896" lane="9" entrytime="00:00:32.00" />
                <RESULT eventid="1446" status="DNS" swimtime="00:00:00.00" resultid="1886" heatid="2924" lane="7" entrytime="00:02:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anita" lastname="Śliwa" birthdate="1972-09-24" gender="F" nation="POL" athleteid="1877">
              <RESULTS>
                <RESULT eventid="1092" points="166" reactiontime="+93" swimtime="00:01:44.37" resultid="1878" heatid="2846" lane="0" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="146" reactiontime="+118" swimtime="00:03:59.25" resultid="1879" heatid="2879" lane="2" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.69" />
                    <SPLIT distance="100" swimtime="00:01:54.25" />
                    <SPLIT distance="150" swimtime="00:03:06.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="171" reactiontime="+96" swimtime="00:00:48.60" resultid="1880" heatid="2906" lane="0" entrytime="00:00:45.00" />
                <RESULT eventid="1462" points="152" reactiontime="+97" swimtime="00:03:50.66" resultid="1881" heatid="2927" lane="7" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.02" />
                    <SPLIT distance="100" swimtime="00:01:51.24" />
                    <SPLIT distance="150" swimtime="00:02:52.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="TMT - 1" number="1">
              <RESULTS>
                <RESULT eventid="1284" reactiontime="+78" swimtime="00:02:30.98" resultid="1897" heatid="3970" lane="7" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.18" />
                    <SPLIT distance="100" swimtime="00:01:19.73" />
                    <SPLIT distance="150" swimtime="00:01:59.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1867" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="1872" number="2" />
                    <RELAYPOSITION athleteid="1877" number="3" reactiontime="+103" />
                    <RELAYPOSITION athleteid="1882" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="TMT - 2" number="2">
              <RESULTS>
                <RESULT eventid="1494" status="DNS" swimtime="00:00:00.00" resultid="1898" heatid="3989" lane="0" entrytime="00:02:45.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1877" number="1" />
                    <RELAYPOSITION athleteid="1887" number="2" />
                    <RELAYPOSITION athleteid="1892" number="3" />
                    <RELAYPOSITION athleteid="1872" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="LTU" clubid="1585" name="Vandenis">
          <ATHLETES>
            <ATHLETE firstname="Sigitas" lastname="Katkevicius" birthdate="1957-08-05" gender="M" nation="LTU" swrid="4418116" athleteid="1586">
              <RESULTS>
                <RESULT eventid="1140" points="372" reactiontime="+83" swimtime="00:00:36.06" resultid="1587" heatid="2858" lane="9" entrytime="00:00:36.78" entrycourse="SCM" />
                <RESULT eventid="1172" points="372" reactiontime="+82" swimtime="00:01:05.20" resultid="1588" heatid="2868" lane="9" entrytime="00:01:05.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="358" reactiontime="+87" swimtime="00:00:29.44" resultid="1589" heatid="2896" lane="5" entrytime="00:00:29.95" entrycourse="SCM" />
                <RESULT eventid="1414" points="353" reactiontime="+90" swimtime="00:01:20.42" resultid="1590" heatid="2916" lane="8" entrytime="00:01:17.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2002" name="5 Styl Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Jakub" lastname="Niedźwiadek" birthdate="1993-10-18" gender="M" nation="POL" athleteid="2012">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="2013" heatid="2843" lane="2" entrytime="00:00:30.50" />
                <RESULT eventid="1172" points="338" reactiontime="+78" swimtime="00:01:07.30" resultid="2014" heatid="2867" lane="4" entrytime="00:01:07.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="338" reactiontime="+80" swimtime="00:00:30.01" resultid="2015" heatid="2897" lane="0" entrytime="00:00:28.00" />
                <RESULT eventid="1414" status="DNS" swimtime="00:00:00.00" resultid="2016" heatid="2916" lane="2" entrytime="00:01:16.00" />
                <RESULT eventid="1446" points="327" reactiontime="+93" swimtime="00:02:27.97" resultid="2826" heatid="2922" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                    <SPLIT distance="100" swimtime="00:01:12.68" />
                    <SPLIT distance="150" swimtime="00:01:50.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Dzikiewicz" birthdate="1990-10-27" gender="M" nation="POL" athleteid="2010">
              <RESULTS>
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="2011" heatid="2895" lane="8" entrytime="00:00:34.00" />
                <RESULT eventid="1140" status="DNS" swimtime="00:00:00.00" resultid="2022" heatid="2856" lane="8" />
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="2023" heatid="2881" lane="6" />
                <RESULT eventid="1446" status="DNS" swimtime="00:00:00.00" resultid="2024" heatid="2921" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Barnasiuk" birthdate="1992-02-04" gender="M" nation="POL" swrid="4273597" athleteid="2017">
              <RESULTS>
                <RESULT eventid="1076" points="431" reactiontime="+71" swimtime="00:00:29.48" resultid="2018" heatid="2843" lane="7" entrytime="00:00:30.50" />
                <RESULT eventid="1140" points="469" reactiontime="+69" swimtime="00:00:33.39" resultid="2019" heatid="2858" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="1318" points="434" reactiontime="+69" swimtime="00:00:27.60" resultid="2020" heatid="2897" lane="8" entrytime="00:00:28.00" />
                <RESULT eventid="1414" points="451" reactiontime="+71" swimtime="00:01:14.14" resultid="2021" heatid="2916" lane="6" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewa" lastname="Łatkowska" birthdate="1965-06-10" gender="F" nation="POL" athleteid="2005">
              <RESULTS>
                <RESULT eventid="1059" points="100" reactiontime="+97" swimtime="00:00:52.55" resultid="2006" heatid="2837" lane="0" entrytime="00:00:52.00" />
                <RESULT eventid="1252" points="135" reactiontime="+85" swimtime="00:04:05.38" resultid="2007" heatid="2879" lane="1" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.48" />
                    <SPLIT distance="100" swimtime="00:02:01.98" />
                    <SPLIT distance="150" swimtime="00:03:08.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="155" reactiontime="+76" swimtime="00:00:44.03" resultid="2008" heatid="2887" lane="7" entrytime="00:00:48.00" />
                <RESULT eventid="1366" points="139" reactiontime="+82" swimtime="00:00:52.06" resultid="2009" heatid="2905" lane="1" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ola" lastname="Dziewa" birthdate="1996-03-26" gender="F" nation="POL" athleteid="2003">
              <RESULTS>
                <RESULT eventid="1301" points="507" reactiontime="+71" swimtime="00:00:29.68" resultid="2004" heatid="2889" lane="3" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1494" reactiontime="+76" swimtime="00:02:28.77" resultid="3318" heatid="3989" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.13" />
                    <SPLIT distance="100" swimtime="00:01:25.48" />
                    <SPLIT distance="150" swimtime="00:01:02.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2005" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="2017" number="2" />
                    <RELAYPOSITION athleteid="2003" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="2012" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="O1" eventid="1284" reactiontime="+68" status="DSQ" swimtime="00:02:07.25" resultid="3319" heatid="3970" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.59" />
                    <SPLIT distance="100" swimtime="00:00:57.12" />
                    <SPLIT distance="150" swimtime="00:01:25.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2017" number="1" reactiontime="+68" status="DSQ" />
                    <RELAYPOSITION athleteid="2012" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="2003" number="3" reactiontime="-5" status="DSQ" />
                    <RELAYPOSITION athleteid="2005" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="01713" nation="POL" region="13" clubid="2130" name="Stow. Pływackie Masters Olsztyn">
          <ATHLETES>
            <ATHLETE firstname="Piotr" lastname="Konopacki" birthdate="1978-04-01" gender="M" nation="POL" license="501713700019" athleteid="2792">
              <RESULTS>
                <RESULT eventid="1108" points="324" reactiontime="+79" swimtime="00:01:15.44" resultid="2793" heatid="2848" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="435" reactiontime="+72" swimtime="00:01:01.87" resultid="2794" heatid="2864" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="416" reactiontime="+74" swimtime="00:02:16.63" resultid="2795" heatid="2921" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                    <SPLIT distance="100" swimtime="00:01:05.85" />
                    <SPLIT distance="150" swimtime="00:01:41.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1478" points="308" reactiontime="+72" swimtime="00:02:45.63" resultid="2796" heatid="2929" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.96" />
                    <SPLIT distance="100" swimtime="00:01:21.73" />
                    <SPLIT distance="150" swimtime="00:02:04.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Lemańczyk" birthdate="1977-10-01" gender="M" nation="POL" license="501713700050" athleteid="2802">
              <RESULTS>
                <RESULT eventid="1172" points="181" reactiontime="+83" swimtime="00:01:22.92" resultid="2803" heatid="2865" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="231" reactiontime="+97" swimtime="00:03:25.42" resultid="2804" heatid="2876" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.76" />
                    <SPLIT distance="100" swimtime="00:01:39.02" />
                    <SPLIT distance="150" swimtime="00:02:33.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1414" points="206" reactiontime="+89" swimtime="00:01:36.28" resultid="2805" heatid="2913" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="177" reactiontime="+91" swimtime="00:03:01.43" resultid="2806" heatid="2921" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.41" />
                    <SPLIT distance="100" swimtime="00:01:25.98" />
                    <SPLIT distance="150" swimtime="00:02:14.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mieszko" lastname="Palmi-Kukiełko" birthdate="1993-09-15" gender="M" nation="POL" license="101713700006" athleteid="2807">
              <RESULTS>
                <RESULT eventid="1204" points="431" reactiontime="+78" swimtime="00:02:26.53" resultid="2808" heatid="2872" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.58" />
                    <SPLIT distance="100" swimtime="00:01:07.41" />
                    <SPLIT distance="150" swimtime="00:01:46.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="513" reactiontime="+78" swimtime="00:02:22.33" resultid="2809" heatid="2881" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.78" />
                    <SPLIT distance="100" swimtime="00:01:06.32" />
                    <SPLIT distance="150" swimtime="00:01:48.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="525" reactiontime="+74" swimtime="00:01:01.26" resultid="2810" heatid="2902" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="470" reactiontime="+79" swimtime="00:02:11.19" resultid="2811" heatid="2922" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.83" />
                    <SPLIT distance="100" swimtime="00:01:03.77" />
                    <SPLIT distance="150" swimtime="00:01:38.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Gregorowicz" birthdate="1974-10-30" gender="M" nation="POL" license="101713700002" athleteid="2812">
              <RESULTS>
                <RESULT eventid="1204" points="434" reactiontime="+81" swimtime="00:02:26.18" resultid="2813" heatid="2872" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                    <SPLIT distance="100" swimtime="00:01:10.39" />
                    <SPLIT distance="150" swimtime="00:01:48.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="436" reactiontime="+75" swimtime="00:02:30.25" resultid="2814" heatid="2881" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.37" />
                    <SPLIT distance="100" swimtime="00:01:12.39" />
                    <SPLIT distance="150" swimtime="00:01:55.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="502" reactiontime="+75" swimtime="00:01:02.20" resultid="2815" heatid="2902" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="477" reactiontime="+74" swimtime="00:02:10.48" resultid="2816" heatid="2921" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.82" />
                    <SPLIT distance="100" swimtime="00:01:03.20" />
                    <SPLIT distance="150" swimtime="00:01:37.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Justyna" lastname="Łagowska" birthdate="1982-06-07" gender="F" nation="POL" license="501713600008" athleteid="2787">
              <RESULTS>
                <RESULT eventid="1092" points="132" swimtime="00:01:52.68" resultid="2788" heatid="2845" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="191" reactiontime="+114" swimtime="00:01:29.72" resultid="2789" heatid="2859" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="205" reactiontime="+134" swimtime="00:00:40.11" resultid="2790" heatid="2886" lane="9" />
                <RESULT eventid="1430" points="174" reactiontime="+118" swimtime="00:03:22.36" resultid="2791" heatid="2917" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.67" />
                    <SPLIT distance="100" swimtime="00:01:33.76" />
                    <SPLIT distance="150" swimtime="00:02:28.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Zaleska" birthdate="1988-01-17" gender="F" nation="POL" license="501713600012" athleteid="2782">
              <RESULTS>
                <RESULT eventid="1059" points="342" reactiontime="+82" swimtime="00:00:34.91" resultid="2783" heatid="2836" lane="4" />
                <RESULT eventid="1188" points="307" reactiontime="+83" swimtime="00:03:00.43" resultid="2784" heatid="2870" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.72" />
                    <SPLIT distance="100" swimtime="00:01:25.42" />
                    <SPLIT distance="150" swimtime="00:02:13.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="345" reactiontime="+87" swimtime="00:01:19.09" resultid="2785" heatid="2899" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1430" points="319" reactiontime="+81" swimtime="00:02:45.26" resultid="2786" heatid="2917" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                    <SPLIT distance="100" swimtime="00:01:18.64" />
                    <SPLIT distance="150" swimtime="00:02:01.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Mówiński" birthdate="1969-09-01" gender="M" nation="POL" license="501713700007" athleteid="2797">
              <RESULTS>
                <RESULT eventid="1140" points="197" reactiontime="+88" swimtime="00:00:44.59" resultid="2798" heatid="2856" lane="0" />
                <RESULT eventid="1268" points="188" reactiontime="+96" swimtime="00:03:18.90" resultid="2799" heatid="2882" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.21" />
                    <SPLIT distance="100" swimtime="00:01:39.38" />
                    <SPLIT distance="150" swimtime="00:02:37.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="174" reactiontime="+88" swimtime="00:01:28.53" resultid="2800" heatid="2902" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1382" points="147" reactiontime="+92" swimtime="00:00:45.04" resultid="2801" heatid="2907" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1284" reactiontime="+74" swimtime="00:02:05.56" resultid="2166" heatid="3970" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.09" />
                    <SPLIT distance="100" swimtime="00:00:52.69" />
                    <SPLIT distance="150" swimtime="00:01:25.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2807" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="2812" number="2" />
                    <RELAYPOSITION athleteid="2782" number="3" reactiontime="+16" />
                    <RELAYPOSITION athleteid="2787" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1494" reactiontime="+86" swimtime="00:02:18.04" resultid="2167" heatid="3989" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.79" />
                    <SPLIT distance="100" swimtime="00:01:03.83" />
                    <SPLIT distance="150" swimtime="00:01:38.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2807" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="2812" number="2" />
                    <RELAYPOSITION athleteid="2782" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="2787" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="EXOBO" nation="POL" clubid="1579" name="KS Extreme Team Oborniki">
          <ATHLETES>
            <ATHLETE firstname="Janusz" lastname="Wolniewicz" birthdate="1948-12-22" gender="M" nation="POL" swrid="4754624" athleteid="1580">
              <RESULTS>
                <RESULT eventid="1318" points="150" reactiontime="+101" swimtime="00:00:39.34" resultid="1581" heatid="2894" lane="7" entrytime="00:00:37.00" />
                <RESULT eventid="1446" points="87" reactiontime="+101" swimtime="00:03:49.35" resultid="1582" heatid="2923" lane="1" entrytime="00:03:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.25" />
                    <SPLIT distance="100" swimtime="00:01:48.87" />
                    <SPLIT distance="150" swimtime="00:02:51.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01709" nation="POL" region="09" clubid="2174" name="iSwim Białystok">
          <ATHLETES>
            <ATHLETE firstname="Dawid" lastname="Świderski" birthdate="1979-02-13" gender="M" nation="POL" license="517/09700108" swrid="5422007" athleteid="2175">
              <RESULTS>
                <RESULT eventid="1076" points="496" reactiontime="+79" swimtime="00:00:28.12" resultid="2176" heatid="2844" lane="1" entrytime="00:00:28.16" entrycourse="LCM" />
                <RESULT eventid="1318" points="475" reactiontime="+76" swimtime="00:00:26.79" resultid="2177" heatid="2898" lane="0" entrytime="00:00:26.54" entrycourse="LCM" />
                <RESULT eventid="1350" points="392" reactiontime="+85" swimtime="00:01:07.52" resultid="2178" heatid="2903" lane="6" entrytime="00:01:04.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Daszuta" birthdate="1973-03-12" gender="M" nation="POL" license="117/09700012" swrid="5421995" athleteid="2179">
              <RESULTS>
                <RESULT eventid="1076" points="432" reactiontime="+79" swimtime="00:00:29.44" resultid="2180" heatid="2841" lane="9" />
                <RESULT eventid="1140" points="419" reactiontime="+82" swimtime="00:00:34.66" resultid="2181" heatid="2855" lane="7" />
                <RESULT eventid="1382" points="288" reactiontime="+88" swimtime="00:00:36.03" resultid="2182" heatid="2907" lane="7" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00115" nation="POL" region="15" clubid="2359" name="KS Warta Poznań">
          <ATHLETES>
            <ATHLETE firstname="Małgorzata" lastname="Putowska" birthdate="1962-01-22" gender="F" nation="POL" license="500115600462" swrid="5416834" athleteid="2408">
              <RESULTS>
                <RESULT eventid="1220" points="171" reactiontime="+96" swimtime="00:04:10.09" resultid="2409" heatid="2874" lane="2" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.97" />
                    <SPLIT distance="100" swimtime="00:01:59.67" />
                    <SPLIT distance="150" swimtime="00:03:04.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="141" swimtime="00:04:02.08" resultid="2410" heatid="2879" lane="7" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.96" />
                    <SPLIT distance="100" swimtime="00:02:00.74" />
                    <SPLIT distance="150" swimtime="00:03:05.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="76" reactiontime="+92" swimtime="00:02:10.84" resultid="2411" heatid="2900" lane="8" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="121" reactiontime="+98" swimtime="00:04:08.82" resultid="2412" heatid="2927" lane="1" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.02" />
                    <SPLIT distance="100" swimtime="00:02:02.30" />
                    <SPLIT distance="150" swimtime="00:03:06.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewa" lastname="Szała" birthdate="1959-03-19" gender="F" nation="POL" license="500115600674" swrid="4302573" athleteid="2365">
              <RESULTS>
                <RESULT eventid="1092" points="227" reactiontime="+89" swimtime="00:01:34.16" resultid="2366" heatid="2845" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="237" reactiontime="+102" swimtime="00:03:23.52" resultid="2367" heatid="2878" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.87" />
                    <SPLIT distance="100" swimtime="00:01:37.95" />
                    <SPLIT distance="150" swimtime="00:02:35.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="239" reactiontime="+87" swimtime="00:00:43.44" resultid="2368" heatid="2904" lane="5" />
                <RESULT eventid="1462" points="225" reactiontime="+100" swimtime="00:03:22.61" resultid="2369" heatid="2926" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.54" />
                    <SPLIT distance="100" swimtime="00:01:39.91" />
                    <SPLIT distance="150" swimtime="00:02:32.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Janyga" birthdate="1966-03-27" gender="M" nation="POL" license="100115700346" swrid="4992782" athleteid="2375">
              <RESULTS>
                <RESULT eventid="1108" points="334" reactiontime="+71" swimtime="00:01:14.67" resultid="2376" heatid="2850" lane="1" entrytime="00:01:12.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1382" points="343" reactiontime="+76" swimtime="00:00:33.98" resultid="2377" heatid="2910" lane="2" entrytime="00:00:33.16" entrycourse="LCM" />
                <RESULT eventid="1446" points="321" reactiontime="+89" swimtime="00:02:28.93" resultid="2378" heatid="2924" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                    <SPLIT distance="100" swimtime="00:01:13.79" />
                    <SPLIT distance="150" swimtime="00:01:51.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Krupińska" birthdate="1953-05-24" gender="F" nation="POL" license="500115600520" swrid="4992790" athleteid="2384">
              <RESULTS>
                <RESULT eventid="1124" points="182" reactiontime="+99" swimtime="00:00:51.64" resultid="2385" heatid="2852" lane="2" entrytime="00:00:53.12" entrycourse="LCM" />
                <RESULT eventid="1220" points="160" reactiontime="+102" swimtime="00:04:15.57" resultid="2386" heatid="2874" lane="1" entrytime="00:04:18.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.31" />
                    <SPLIT distance="100" swimtime="00:02:06.07" />
                    <SPLIT distance="150" swimtime="00:03:12.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="110" reactiontime="+99" swimtime="00:00:49.36" resultid="2387" heatid="2887" lane="8" entrytime="00:00:49.85" entrycourse="LCM" />
                <RESULT eventid="1398" points="156" reactiontime="+109" swimtime="00:01:59.07" resultid="2388" heatid="2911" lane="6" entrytime="00:02:00.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Wieja" birthdate="1978-09-08" gender="M" nation="POL" license="500115700467" swrid="5331775" athleteid="2379">
              <RESULTS>
                <RESULT eventid="1108" points="338" reactiontime="+64" swimtime="00:01:14.42" resultid="2380" heatid="2850" lane="3" entrytime="00:01:09.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="2381" heatid="2883" lane="5" entrytime="00:02:30.00" />
                <RESULT eventid="1318" points="410" reactiontime="+64" swimtime="00:00:28.14" resultid="2382" heatid="2897" lane="5" entrytime="00:00:27.00" />
                <RESULT eventid="1382" points="385" reactiontime="+71" swimtime="00:00:32.69" resultid="2383" heatid="2910" lane="3" entrytime="00:00:32.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Waraczewski" birthdate="1962-04-19" gender="M" nation="POL" license="100115700344" swrid="4992781" athleteid="2399">
              <RESULTS>
                <RESULT eventid="1140" points="265" reactiontime="+96" swimtime="00:00:40.39" resultid="2400" heatid="2857" lane="6" entrytime="00:00:42.00" />
                <RESULT eventid="1236" points="257" reactiontime="+93" swimtime="00:03:18.34" resultid="2401" heatid="2877" lane="1" entrytime="00:03:21.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.08" />
                    <SPLIT distance="100" swimtime="00:01:34.56" />
                    <SPLIT distance="150" swimtime="00:02:26.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1414" points="248" reactiontime="+91" swimtime="00:01:30.49" resultid="2402" heatid="2915" lane="1" entrytime="00:01:31.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sylwia" lastname="Gorockiewicz" birthdate="1975-03-29" gender="F" nation="POL" license="500115600525" swrid="4837788" athleteid="2389">
              <RESULTS>
                <RESULT eventid="1124" points="91" reactiontime="+107" swimtime="00:01:05.08" resultid="2390" heatid="2852" lane="7" entrytime="00:00:59.00" />
                <RESULT eventid="1220" points="100" reactiontime="+93" swimtime="00:04:58.62" resultid="2391" heatid="2874" lane="8" entrytime="00:04:49.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.04" />
                    <SPLIT distance="100" swimtime="00:02:24.01" />
                    <SPLIT distance="150" swimtime="00:03:42.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="58" reactiontime="+139" swimtime="00:01:00.90" resultid="2392" heatid="2886" lane="5" entrytime="00:00:57.98" entrycourse="LCM" />
                <RESULT eventid="1398" points="92" reactiontime="+129" swimtime="00:02:21.57" resultid="2393" heatid="2911" lane="7" entrytime="00:02:18.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Kotecka" birthdate="1965-05-08" gender="F" nation="POL" license="100115600357" swrid="4754727" athleteid="2360">
              <RESULTS>
                <RESULT eventid="1092" points="172" reactiontime="+124" swimtime="00:01:43.29" resultid="2361" heatid="2846" lane="9" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="220" reactiontime="+105" swimtime="00:01:25.53" resultid="2362" heatid="2861" lane="1" entrytime="00:01:28.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1430" points="224" reactiontime="+106" swimtime="00:03:06.01" resultid="2363" heatid="2918" lane="4" entrytime="00:03:10.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.61" />
                    <SPLIT distance="100" swimtime="00:01:30.74" />
                    <SPLIT distance="150" swimtime="00:02:19.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="185" reactiontime="+103" swimtime="00:03:36.41" resultid="2364" heatid="2927" lane="2" entrytime="00:03:38.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.79" />
                    <SPLIT distance="100" swimtime="00:01:47.56" />
                    <SPLIT distance="150" swimtime="00:02:43.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Lesiński" birthdate="1944-04-13" gender="M" nation="POL" license="500115700616" swrid="4188190" athleteid="2370">
              <RESULTS>
                <RESULT eventid="1108" points="102" reactiontime="+85" swimtime="00:01:50.66" resultid="2371" heatid="2848" lane="4" entrytime="00:01:57.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="101" reactiontime="+108" swimtime="00:01:40.55" resultid="2372" heatid="2866" lane="9" entrytime="00:01:42.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1382" points="114" reactiontime="+83" swimtime="00:00:48.98" resultid="2373" heatid="2909" lane="0" entrytime="00:00:50.51" entrycourse="LCM" />
                <RESULT eventid="1478" points="96" reactiontime="+82" swimtime="00:04:03.61" resultid="2374" heatid="2929" lane="3" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.23" />
                    <SPLIT distance="100" swimtime="00:01:58.74" />
                    <SPLIT distance="150" swimtime="00:03:03.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Szymkowiak" birthdate="1980-04-12" gender="M" nation="POL" license="500115700523" swrid="5312534" athleteid="2403">
              <RESULTS>
                <RESULT eventid="1140" points="541" reactiontime="+78" swimtime="00:00:31.84" resultid="2404" heatid="2858" lane="5" entrytime="00:00:30.42" entrycourse="LCM" />
                <RESULT eventid="1172" points="454" reactiontime="+82" swimtime="00:01:01.03" resultid="2405" heatid="2869" lane="1" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="432" reactiontime="+76" swimtime="00:00:27.65" resultid="2406" heatid="2898" lane="8" entrytime="00:00:26.32" entrycourse="LCM" />
                <RESULT eventid="1414" points="497" reactiontime="+75" swimtime="00:01:11.80" resultid="2407" heatid="2916" lane="5" entrytime="00:01:07.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grażyna" lastname="Drela" birthdate="1957-10-01" gender="F" nation="POL" license="500115700493" swrid="4269916" athleteid="2394">
              <RESULTS>
                <RESULT eventid="1124" points="239" reactiontime="+106" swimtime="00:00:47.19" resultid="2395" heatid="2853" lane="0" entrytime="00:00:45.00" />
                <RESULT eventid="1156" points="215" reactiontime="+86" swimtime="00:01:26.24" resultid="2396" heatid="2861" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="240" reactiontime="+90" swimtime="00:00:38.05" resultid="2397" heatid="2887" lane="5" entrytime="00:00:41.00" />
                <RESULT eventid="1366" points="224" reactiontime="+85" swimtime="00:00:44.39" resultid="2398" heatid="2906" lane="8" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1284" reactiontime="+69" swimtime="00:02:15.07" resultid="2413" heatid="3969" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.85" />
                    <SPLIT distance="100" swimtime="00:01:06.98" />
                    <SPLIT distance="150" swimtime="00:01:36.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2379" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="2365" number="2" />
                    <RELAYPOSITION athleteid="2375" number="3" reactiontime="+18" />
                    <RELAYPOSITION athleteid="2360" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1494" reactiontime="+72" swimtime="00:02:31.53" resultid="2415" heatid="3988" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.85" />
                    <SPLIT distance="100" swimtime="00:01:05.22" />
                    <SPLIT distance="150" swimtime="00:01:52.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2379" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="2403" number="2" />
                    <RELAYPOSITION athleteid="2365" number="3" reactiontime="+67" />
                    <RELAYPOSITION athleteid="2360" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1284" reactiontime="+90" swimtime="00:03:12.60" resultid="2414" heatid="3969" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.06" />
                    <SPLIT distance="100" swimtime="00:01:27.81" />
                    <SPLIT distance="150" swimtime="00:02:27.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2399" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="2384" number="2" />
                    <RELAYPOSITION athleteid="2389" number="3" reactiontime="+100" />
                    <RELAYPOSITION athleteid="2370" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1494" reactiontime="+88" swimtime="00:03:05.32" resultid="2416" heatid="3987" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.05" />
                    <SPLIT distance="100" swimtime="00:01:31.40" />
                    <SPLIT distance="150" swimtime="00:02:26.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2370" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="2399" number="2" />
                    <RELAYPOSITION athleteid="2408" number="3" />
                    <RELAYPOSITION athleteid="2394" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="03503" nation="POL" region="03" clubid="2447" name="MASTERS Lublin">
          <ATHLETES>
            <ATHLETE firstname="Anna" lastname="Wójcicka" birthdate="1975-05-28" gender="F" nation="POL" license="103503600002" athleteid="2458">
              <RESULTS>
                <RESULT eventid="1092" points="276" reactiontime="+102" swimtime="00:01:28.14" resultid="2459" heatid="2845" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="308" reactiontime="+99" swimtime="00:00:39.94" resultid="2460" heatid="2904" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mirosław" lastname="Molenda" birthdate="1971-12-11" gender="M" nation="POL" license="103503700012" athleteid="2448">
              <RESULTS>
                <RESULT eventid="1076" points="178" reactiontime="+102" swimtime="00:00:39.56" resultid="2449" heatid="2840" lane="5" />
                <RESULT eventid="1172" points="197" reactiontime="+97" swimtime="00:01:20.54" resultid="2450" heatid="2864" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="207" reactiontime="+93" swimtime="00:00:35.33" resultid="2451" heatid="2891" lane="4" />
                <RESULT eventid="1446" points="178" reactiontime="+101" swimtime="00:03:01.30" resultid="2452" heatid="2921" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                    <SPLIT distance="100" swimtime="00:01:27.54" />
                    <SPLIT distance="150" swimtime="00:02:15.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Konrad" lastname="Ćwikła" birthdate="1975-11-07" gender="M" nation="POL" license="103503700005" swrid="5241236" athleteid="2461">
              <RESULTS>
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="2462" heatid="2848" lane="9" />
                <RESULT eventid="1318" points="334" reactiontime="+85" swimtime="00:00:30.13" resultid="2463" heatid="2892" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Wójcicki" birthdate="1975-04-28" gender="M" nation="POL" license="103503700001" swrid="5455050" athleteid="2469">
              <RESULTS>
                <RESULT eventid="1140" points="235" reactiontime="+84" swimtime="00:00:42.02" resultid="2470" heatid="2855" lane="5" />
                <RESULT eventid="1414" points="211" reactiontime="+94" swimtime="00:01:35.53" resultid="2471" heatid="2913" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Staszek" birthdate="1976-02-23" gender="M" nation="POL" license="103503700013" athleteid="2453">
              <RESULTS>
                <RESULT eventid="1076" points="155" reactiontime="+124" swimtime="00:00:41.44" resultid="2454" heatid="2840" lane="6" />
                <RESULT eventid="1172" points="224" reactiontime="+92" swimtime="00:01:17.19" resultid="2455" heatid="2864" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1382" points="180" reactiontime="+93" swimtime="00:00:42.12" resultid="2456" heatid="2908" lane="0" />
                <RESULT eventid="1414" points="215" reactiontime="+95" swimtime="00:01:34.89" resultid="2457" heatid="2913" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Pietrzak" birthdate="1988-10-21" gender="M" nation="POL" license="103503700011" athleteid="2464">
              <RESULTS>
                <RESULT eventid="1108" points="289" reactiontime="+91" swimtime="00:01:18.37" resultid="2465" heatid="2848" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="296" reactiontime="+74" swimtime="00:03:09.18" resultid="2466" heatid="2876" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.44" />
                    <SPLIT distance="100" swimtime="00:01:28.27" />
                    <SPLIT distance="150" swimtime="00:02:18.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1382" points="327" reactiontime="+86" swimtime="00:00:34.54" resultid="2467" heatid="2908" lane="7" />
                <RESULT eventid="1446" points="239" reactiontime="+79" swimtime="00:02:44.16" resultid="2468" heatid="2921" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                    <SPLIT distance="100" swimtime="00:01:18.06" />
                    <SPLIT distance="150" swimtime="00:02:02.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02202" nation="POL" region="02" clubid="2472" name="MKS Astoria Bydgoszcz">
          <ATHLETES>
            <ATHLETE firstname="Dariusz" lastname="Kostkowski" birthdate="1970-01-13" gender="M" nation="POL" license="102202700126" swrid="5471726" athleteid="2488">
              <RESULTS>
                <RESULT eventid="1140" points="173" reactiontime="+84" swimtime="00:00:46.52" resultid="2489" heatid="2856" lane="6" entrytime="00:00:52.86" entrycourse="LCM" />
                <RESULT eventid="1236" points="120" reactiontime="+76" swimtime="00:04:15.23" resultid="2490" heatid="2875" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.60" />
                    <SPLIT distance="100" swimtime="00:02:01.77" />
                    <SPLIT distance="150" swimtime="00:03:09.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1414" points="134" reactiontime="+74" swimtime="00:01:51.03" resultid="2491" heatid="2913" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1478" points="80" reactiontime="+104" swimtime="00:04:19.49" resultid="2492" heatid="2928" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.07" />
                    <SPLIT distance="100" swimtime="00:02:07.84" />
                    <SPLIT distance="150" swimtime="00:03:15.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Ciężki" birthdate="1994-09-30" gender="M" nation="POL" license="102202700137" swrid="4289450" athleteid="2483">
              <RESULTS>
                <RESULT eventid="1108" points="400" reactiontime="+75" swimtime="00:01:10.33" resultid="2484" heatid="2850" lane="4" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="499" reactiontime="+84" swimtime="00:00:59.14" resultid="2485" heatid="2865" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="487" reactiontime="+81" swimtime="00:00:26.57" resultid="2486" heatid="2892" lane="4" />
                <RESULT eventid="1478" points="370" reactiontime="+79" swimtime="00:02:35.85" resultid="2487" heatid="2930" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                    <SPLIT distance="100" swimtime="00:01:13.44" />
                    <SPLIT distance="150" swimtime="00:01:54.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Dudek" birthdate="2001-06-20" gender="F" nation="POL" license="102202600128" swrid="4001627" athleteid="2473">
              <RESULTS>
                <RESULT eventid="1059" points="475" reactiontime="+81" swimtime="00:00:31.31" resultid="2474" heatid="2838" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1156" points="537" reactiontime="+79" swimtime="00:01:03.61" resultid="2475" heatid="2862" lane="3" entrytime="00:01:03.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="540" reactiontime="+80" swimtime="00:00:29.06" resultid="2476" heatid="2889" lane="6" entrytime="00:00:28.50" />
                <RESULT eventid="1430" points="520" reactiontime="+78" swimtime="00:02:20.45" resultid="2477" heatid="2919" lane="5" entrytime="00:02:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                    <SPLIT distance="100" swimtime="00:01:08.06" />
                    <SPLIT distance="150" swimtime="00:01:44.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hanna" lastname="Bakuniak" birthdate="1996-03-25" gender="F" nation="POL" license="102202600136" swrid="4169734" athleteid="2478">
              <RESULTS>
                <RESULT eventid="1092" points="445" reactiontime="+82" swimtime="00:01:15.22" resultid="2479" heatid="2846" lane="6" entrytime="00:01:13.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="465" reactiontime="+70" swimtime="00:01:06.71" resultid="2480" heatid="2862" lane="6" entrytime="00:01:04.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1430" points="532" reactiontime="+71" swimtime="00:02:19.37" resultid="2481" heatid="2919" lane="3" entrytime="00:02:16.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                    <SPLIT distance="100" swimtime="00:01:07.26" />
                    <SPLIT distance="150" swimtime="00:01:44.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="425" reactiontime="+78" swimtime="00:02:44.06" resultid="2482" heatid="2927" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.91" />
                    <SPLIT distance="100" swimtime="00:01:17.40" />
                    <SPLIT distance="150" swimtime="00:01:59.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04303" nation="POL" region="03" clubid="2423" name="Masters Avia Świdnik">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Sitkowski" birthdate="1974-10-05" gender="M" nation="POL" license="504303700001" swrid="5439542" athleteid="2439">
              <RESULTS>
                <RESULT eventid="1108" points="304" reactiontime="+72" swimtime="00:01:17.09" resultid="2440" heatid="2850" lane="8" entrytime="00:01:14.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="271" reactiontime="+82" swimtime="00:02:56.14" resultid="2441" heatid="2883" lane="7" entrytime="00:02:56.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                    <SPLIT distance="100" swimtime="00:01:23.40" />
                    <SPLIT distance="150" swimtime="00:02:15.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1382" points="330" reactiontime="+70" swimtime="00:00:34.43" resultid="2442" heatid="2910" lane="1" entrytime="00:00:33.99" entrycourse="LCM" />
                <RESULT eventid="1478" points="268" reactiontime="+73" swimtime="00:02:53.57" resultid="2443" heatid="2930" lane="2" entrytime="00:02:48.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                    <SPLIT distance="100" swimtime="00:01:23.97" />
                    <SPLIT distance="150" swimtime="00:02:09.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Zielonka" birthdate="1986-05-26" gender="M" nation="POL" license="104303700006" swrid="4061691" athleteid="2424">
              <RESULTS>
                <RESULT eventid="1076" points="488" reactiontime="+82" swimtime="00:00:28.28" resultid="2425" heatid="2844" lane="8" entrytime="00:00:28.77" entrycourse="LCM" />
                <RESULT eventid="1172" points="523" reactiontime="+77" swimtime="00:00:58.20" resultid="2426" heatid="2869" lane="7" entrytime="00:00:58.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="479" reactiontime="+75" swimtime="00:00:26.71" resultid="2427" heatid="2898" lane="1" entrytime="00:00:26.31" entrycourse="LCM" />
                <RESULT eventid="1446" points="489" reactiontime="+77" swimtime="00:02:09.41" resultid="2428" heatid="2925" lane="3" entrytime="00:02:07.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.15" />
                    <SPLIT distance="100" swimtime="00:01:03.10" />
                    <SPLIT distance="150" swimtime="00:01:36.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cezary" lastname="Lipiński" birthdate="1972-04-11" gender="M" nation="POL" license="104303700002" swrid="5449345" athleteid="2429">
              <RESULTS>
                <RESULT eventid="1076" points="265" reactiontime="+72" swimtime="00:00:34.63" resultid="2430" heatid="2843" lane="0" entrytime="00:00:33.96" entrycourse="LCM" />
                <RESULT eventid="1204" reactiontime="+86" status="DNF" swimtime="00:00:00.00" resultid="2431" heatid="2872" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.20" />
                    <SPLIT distance="100" swimtime="00:01:41.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="340" reactiontime="+82" swimtime="00:00:29.94" resultid="2432" heatid="2896" lane="2" entrytime="00:00:30.43" entrycourse="LCM" />
                <RESULT eventid="1446" points="309" reactiontime="+84" swimtime="00:02:30.81" resultid="2433" heatid="2924" lane="5" entrytime="00:02:32.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.83" />
                    <SPLIT distance="100" swimtime="00:01:13.80" />
                    <SPLIT distance="150" swimtime="00:01:52.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Mazur" birthdate="1995-03-13" gender="M" nation="POL" license="104303700009" swrid="4195380" athleteid="2434">
              <RESULTS>
                <RESULT eventid="1076" points="523" reactiontime="+67" swimtime="00:00:27.64" resultid="2435" heatid="2844" lane="2" entrytime="00:00:27.50" />
                <RESULT eventid="1172" points="603" reactiontime="+67" swimtime="00:00:55.52" resultid="2436" heatid="2869" lane="6" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="568" reactiontime="+63" swimtime="00:00:25.24" resultid="2437" heatid="2898" lane="3" entrytime="00:00:26.00" />
                <RESULT eventid="1350" points="422" reactiontime="+66" swimtime="00:01:05.88" resultid="2438" heatid="2903" lane="2" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edyta" lastname="Lipiec" birthdate="1973-03-19" gender="F" nation="POL" license="504303600010" athleteid="2444">
              <RESULTS>
                <RESULT eventid="1156" points="248" swimtime="00:01:22.22" resultid="2445" heatid="2860" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="281" swimtime="00:00:36.12" resultid="2446" heatid="2886" lane="0" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="LTU" clubid="1764" name="Marijampoles TORPEDOS">
          <ATHLETES>
            <ATHLETE firstname="Jurate" lastname="Pranckeviciene" birthdate="1975-05-04" gender="F" nation="LTU" swrid="4754695" athleteid="1765">
              <RESULTS>
                <RESULT eventid="1156" status="DNS" swimtime="00:00:00.00" resultid="1766" heatid="2861" lane="6" entrytime="00:01:20.16" entrycourse="LCM" />
                <RESULT eventid="1301" status="DNS" swimtime="00:00:00.00" resultid="1767" heatid="2888" lane="8" entrytime="00:00:35.08" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Margarita" lastname="Cineliene" birthdate="1956-02-07" gender="F" nation="LTU" swrid="4301763" athleteid="1768">
              <RESULTS>
                <RESULT eventid="1124" points="186" reactiontime="+100" swimtime="00:00:51.31" resultid="1769" heatid="2852" lane="6" entrytime="00:00:50.35" entrycourse="LCM" />
                <RESULT eventid="1220" points="162" swimtime="00:04:14.63" resultid="1770" heatid="2874" lane="7" entrytime="00:04:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.10" />
                    <SPLIT distance="100" swimtime="00:02:00.46" />
                    <SPLIT distance="150" swimtime="00:03:07.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="137" reactiontime="+66" swimtime="00:00:45.88" resultid="1771" heatid="2887" lane="1" entrytime="00:00:48.00" entrycourse="LCM" />
                <RESULT eventid="1398" points="178" reactiontime="+73" swimtime="00:01:53.93" resultid="1772" heatid="2911" lane="3" entrytime="00:01:55.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vilmantas" lastname="Krasauskas" birthdate="1964-07-31" gender="M" nation="LTU" swrid="4199476" athleteid="1778">
              <RESULTS>
                <RESULT eventid="1172" points="351" reactiontime="+83" swimtime="00:01:06.47" resultid="1779" heatid="2868" lane="0" entrytime="00:01:05.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="332" reactiontime="+86" swimtime="00:00:30.18" resultid="1780" heatid="2896" lane="6" entrytime="00:00:30.11" entrycourse="LCM" />
                <RESULT eventid="1446" points="311" reactiontime="+81" swimtime="00:02:30.47" resultid="1781" heatid="2925" lane="1" entrytime="00:02:27.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.36" />
                    <SPLIT distance="100" swimtime="00:01:12.19" />
                    <SPLIT distance="150" swimtime="00:01:51.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Saulius" lastname="Brazukas" birthdate="1964-05-06" gender="M" nation="LTU" swrid="5186202" athleteid="1782">
              <RESULTS>
                <RESULT eventid="1108" points="101" reactiontime="+80" swimtime="00:01:51.22" resultid="1783" heatid="2849" lane="9" entrytime="00:01:53.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="102" reactiontime="+111" swimtime="00:04:03.54" resultid="1784" heatid="2882" lane="2" entrytime="00:04:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.93" />
                    <SPLIT distance="100" swimtime="00:01:55.21" />
                    <SPLIT distance="150" swimtime="00:03:03.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1382" points="111" reactiontime="+82" swimtime="00:00:49.46" resultid="1785" heatid="2909" lane="9" entrytime="00:00:51.93" entrycourse="LCM" />
                <RESULT eventid="1478" points="90" reactiontime="+81" swimtime="00:04:09.54" resultid="1786" heatid="2929" lane="1" entrytime="00:04:33.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.10" />
                    <SPLIT distance="100" swimtime="00:01:59.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stasys" lastname="Grigas" birthdate="1941-03-14" gender="M" nation="LTU" swrid="4777051" athleteid="1773">
              <RESULTS>
                <RESULT eventid="1108" points="32" reactiontime="+130" swimtime="00:02:42.79" resultid="1774" heatid="2848" lane="2" entrytime="00:02:39.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="25" reactiontime="+150" swimtime="00:07:07.42" resultid="1775" heatid="2876" lane="2" entrytime="00:06:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:42.59" />
                    <SPLIT distance="100" swimtime="00:03:34.63" />
                    <SPLIT distance="150" swimtime="00:05:23.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="22" swimtime="00:06:02.74" resultid="1776" heatid="2922" lane="7" entrytime="00:05:51.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:22.87" />
                    <SPLIT distance="100" swimtime="00:03:03.20" />
                    <SPLIT distance="150" swimtime="00:04:38.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1478" points="34" reactiontime="+132" swimtime="00:05:44.98" resultid="1777" heatid="2929" lane="0" entrytime="00:06:20.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:25.71" />
                    <SPLIT distance="100" swimtime="00:02:54.75" />
                    <SPLIT distance="150" swimtime="00:04:23.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00607" nation="POL" region="07" clubid="2619" name="TP Masters Opole">
          <ATHLETES>
            <ATHLETE firstname="Zbigniew" lastname="Januszkiewicz" birthdate="1962-08-18" gender="M" nation="POL" license="100607700003" swrid="4843497" athleteid="2627">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1108" points="410" reactiontime="+66" swimtime="00:01:09.77" resultid="2628" heatid="2850" lane="2" entrytime="00:01:10.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1382" points="404" reactiontime="+68" swimtime="00:00:32.17" resultid="2629" heatid="2910" lane="6" entrytime="00:00:32.47" entrycourse="LCM" />
                <RESULT comment="Rekord Polski Masters" eventid="1478" points="396" reactiontime="+68" swimtime="00:02:32.34" resultid="2630" heatid="2930" lane="3" entrytime="00:02:34.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                    <SPLIT distance="100" swimtime="00:01:15.17" />
                    <SPLIT distance="150" swimtime="00:01:54.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Bartnikowska" birthdate="1990-08-21" gender="F" nation="POL" license="100607600002" swrid="5295108" athleteid="2624">
              <RESULTS>
                <RESULT eventid="1092" points="435" reactiontime="+73" swimtime="00:01:15.79" resultid="2625" heatid="2846" lane="3" entrytime="00:01:12.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="512" reactiontime="+78" swimtime="00:00:33.72" resultid="2626" heatid="2906" lane="3" entrytime="00:00:33.01" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Vogel" birthdate="1981-09-20" gender="M" nation="POL" license="100607700016" swrid="5506641" athleteid="2620">
              <RESULTS>
                <RESULT eventid="1076" points="450" reactiontime="+76" swimtime="00:00:29.06" resultid="2621" heatid="2841" lane="2" />
                <RESULT eventid="1268" points="346" reactiontime="+83" swimtime="00:02:42.34" resultid="2622" heatid="2881" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.16" />
                    <SPLIT distance="100" swimtime="00:01:13.72" />
                    <SPLIT distance="150" swimtime="00:02:03.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="310" reactiontime="+77" swimtime="00:01:13.04" resultid="2623" heatid="2901" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06306" nation="POL" region="06" clubid="2271" name="KS Korona 1919">
          <ATHLETES>
            <ATHLETE firstname="Mariola" lastname="Kuliś" birthdate="1966-07-27" gender="F" nation="POL" license="506306600043" swrid="4992797" athleteid="2272">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1059" points="363" reactiontime="+80" swimtime="00:00:34.22" resultid="2273" heatid="2838" lane="8" entrytime="00:00:34.84" entrycourse="LCM" />
                <RESULT comment="Rekord Polski Masters" eventid="1124" points="415" reactiontime="+84" swimtime="00:00:39.27" resultid="2274" heatid="2853" lane="7" entrytime="00:00:40.53" entrycourse="LCM" />
                <RESULT comment="Rekord Polski Masters" eventid="1301" points="424" reactiontime="+72" swimtime="00:00:31.49" resultid="2275" heatid="2889" lane="1" entrytime="00:00:31.92" entrycourse="LCM" />
                <RESULT eventid="1398" points="343" reactiontime="+75" swimtime="00:01:31.57" resultid="2276" heatid="2912" lane="0" entrytime="00:01:41.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Pycia" birthdate="1966-02-21" gender="M" nation="POL" license="506306700057" swrid="4992712" athleteid="2336">
              <RESULTS>
                <RESULT eventid="1140" points="276" reactiontime="+89" swimtime="00:00:39.82" resultid="2337" heatid="2855" lane="4" />
                <RESULT eventid="1268" points="225" reactiontime="+105" swimtime="00:03:07.43" resultid="2338" heatid="2881" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.40" />
                    <SPLIT distance="150" swimtime="00:02:24.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="288" reactiontime="+95" swimtime="00:00:31.63" resultid="2339" heatid="2891" lane="5" />
                <RESULT eventid="1414" points="243" reactiontime="+98" swimtime="00:01:31.12" resultid="2340" heatid="2913" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Damian" lastname="Jośko" birthdate="1994-07-25" gender="M" nation="POL" license="506306700035" swrid="5484409" athleteid="2346">
              <RESULTS>
                <RESULT eventid="1172" points="336" reactiontime="+71" swimtime="00:01:07.42" resultid="2347" heatid="2864" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="373" reactiontime="+73" swimtime="00:00:29.04" resultid="2348" heatid="2892" lane="5" />
                <RESULT eventid="1382" points="299" reactiontime="+77" swimtime="00:00:35.57" resultid="2349" heatid="2908" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Łysiak" birthdate="1973-03-30" gender="M" nation="POL" license="506306700047" swrid="5468085" athleteid="2326">
              <RESULTS>
                <RESULT eventid="1140" points="274" reactiontime="+82" swimtime="00:00:39.93" resultid="2327" heatid="2855" lane="8" />
                <RESULT eventid="1236" points="311" reactiontime="+78" swimtime="00:03:05.96" resultid="2328" heatid="2877" lane="2" entrytime="00:03:10.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.82" />
                    <SPLIT distance="100" swimtime="00:01:31.03" />
                    <SPLIT distance="150" swimtime="00:02:17.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="260" reactiontime="+101" swimtime="00:00:32.76" resultid="2329" heatid="2893" lane="9" />
                <RESULT eventid="1414" points="263" reactiontime="+95" swimtime="00:01:28.69" resultid="2330" heatid="2915" lane="6" entrytime="00:01:25.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Leńczowska-Tomaszewska" birthdate="1982-01-15" gender="F" nation="POL" license="506306600071" swrid="4992907" athleteid="2302">
              <RESULTS>
                <RESULT eventid="1092" points="327" reactiontime="+79" swimtime="00:01:23.34" resultid="2303" heatid="2846" lane="7" entrytime="00:01:23.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="342" reactiontime="+85" swimtime="00:01:13.89" resultid="2304" heatid="2859" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="424" reactiontime="+84" swimtime="00:00:31.49" resultid="2305" heatid="2888" lane="3" entrytime="00:00:33.99" entrycourse="LCM" />
                <RESULT eventid="1366" points="352" reactiontime="+77" swimtime="00:00:38.19" resultid="2306" heatid="2906" lane="7" entrytime="00:00:38.42" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Borek" birthdate="1991-01-01" gender="M" nation="POL" license="506306700069" swrid="5468079" athleteid="2307">
              <RESULTS>
                <RESULT eventid="1108" points="326" reactiontime="+65" swimtime="00:01:15.30" resultid="2308" heatid="2849" lane="4" entrytime="00:01:17.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="297" reactiontime="+68" swimtime="00:00:38.86" resultid="2309" heatid="2857" lane="5" entrytime="00:00:38.36" entrycourse="LCM" />
                <RESULT eventid="1382" points="337" reactiontime="+68" swimtime="00:00:34.19" resultid="2310" heatid="2908" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Mleczko" birthdate="1947-08-26" gender="M" nation="POL" license="506306700050" swrid="4992812" athleteid="2297">
              <RESULTS>
                <RESULT eventid="1076" points="95" reactiontime="+110" swimtime="00:00:48.79" resultid="2298" heatid="2842" lane="8" entrytime="00:00:49.46" entrycourse="LCM" />
                <RESULT eventid="1172" points="171" reactiontime="+121" swimtime="00:01:24.46" resultid="2299" heatid="2866" lane="6" entrytime="00:01:23.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="188" reactiontime="+105" swimtime="00:00:36.47" resultid="2300" heatid="2894" lane="6" entrytime="00:00:36.58" entrycourse="LCM" />
                <RESULT eventid="1446" points="107" reactiontime="+125" swimtime="00:03:34.66" resultid="2301" heatid="2923" lane="7" entrytime="00:03:25.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.31" />
                    <SPLIT distance="100" swimtime="00:01:42.88" />
                    <SPLIT distance="150" swimtime="00:02:42.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariusz" lastname="Baranik" birthdate="1969-06-29" gender="M" nation="POL" license="506306700027" swrid="4992740" athleteid="2282">
              <RESULTS>
                <RESULT eventid="1076" points="439" reactiontime="+76" swimtime="00:00:29.30" resultid="2283" heatid="2844" lane="9" entrytime="00:00:29.15" entrycourse="LCM" />
                <RESULT eventid="1172" points="450" reactiontime="+73" swimtime="00:01:01.20" resultid="2284" heatid="2869" lane="9" entrytime="00:01:01.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="456" reactiontime="+72" swimtime="00:00:27.16" resultid="2285" heatid="2897" lane="3" entrytime="00:00:27.02" entrycourse="LCM" />
                <RESULT eventid="1414" points="336" reactiontime="+77" swimtime="00:01:21.76" resultid="2286" heatid="2915" lane="4" entrytime="00:01:20.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Waldemar" lastname="Piszczek" birthdate="1962-11-10" gender="M" nation="POL" license="506306700055" swrid="4992814" athleteid="2287">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1076" points="350" reactiontime="+86" swimtime="00:00:31.59" resultid="2288" heatid="2839" lane="3" />
                <RESULT eventid="1140" points="332" reactiontime="+94" swimtime="00:00:37.47" resultid="2289" heatid="2854" lane="3" />
                <RESULT eventid="1350" points="258" reactiontime="+99" swimtime="00:01:17.64" resultid="2290" heatid="2901" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1478" status="DNS" swimtime="00:00:00.00" resultid="2291" heatid="2928" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Jawień" birthdate="1971-06-11" gender="M" nation="POL" license="506306700034" swrid="5468083" athleteid="2316">
              <RESULTS>
                <RESULT eventid="1108" points="263" reactiontime="+76" swimtime="00:01:20.86" resultid="2317" heatid="2847" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="298" reactiontime="+83" swimtime="00:03:08.67" resultid="2318" heatid="2877" lane="6" entrytime="00:03:05.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.51" />
                    <SPLIT distance="100" swimtime="00:01:29.02" />
                    <SPLIT distance="150" swimtime="00:02:18.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1414" points="293" reactiontime="+81" swimtime="00:01:25.58" resultid="2319" heatid="2915" lane="3" entrytime="00:01:23.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1478" points="235" reactiontime="+82" swimtime="00:03:01.12" resultid="2320" heatid="2930" lane="8" entrytime="00:02:56.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.34" />
                    <SPLIT distance="100" swimtime="00:01:27.29" />
                    <SPLIT distance="150" swimtime="00:02:15.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Waga" birthdate="1940-07-04" gender="M" nation="POL" license="506306700064" swrid="4992823" athleteid="2331">
              <RESULTS>
                <RESULT eventid="1140" points="43" reactiontime="+116" swimtime="00:01:13.93" resultid="2332" heatid="2856" lane="1" entrytime="00:01:20.27" entrycourse="LCM" />
                <RESULT eventid="1172" points="59" reactiontime="+117" swimtime="00:01:59.95" resultid="2333" heatid="2865" lane="5" entrytime="00:02:00.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="72" reactiontime="+109" swimtime="00:00:50.26" resultid="2334" heatid="2893" lane="7" entrytime="00:00:52.12" entrycourse="LCM" />
                <RESULT eventid="1446" points="55" reactiontime="+91" swimtime="00:04:27.68" resultid="2335" heatid="2922" lane="2" entrytime="00:04:42.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.56" />
                    <SPLIT distance="100" swimtime="00:02:08.10" />
                    <SPLIT distance="150" swimtime="00:03:19.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Wysocka" birthdate="1988-10-27" gender="F" nation="POL" license="506306600075" swrid="4060957" athleteid="2277">
              <RESULTS>
                <RESULT eventid="1059" points="342" reactiontime="+90" swimtime="00:00:34.93" resultid="2278" heatid="2836" lane="3" />
                <RESULT eventid="1188" status="DNS" swimtime="00:00:00.00" resultid="2279" heatid="2870" lane="6" />
                <RESULT eventid="1334" points="295" reactiontime="+51" swimtime="00:01:23.29" resultid="2280" heatid="2899" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1430" points="376" reactiontime="+96" swimtime="00:02:36.43" resultid="2281" heatid="2917" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                    <SPLIT distance="100" swimtime="00:01:16.89" />
                    <SPLIT distance="150" swimtime="00:01:57.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Orlewicz- Musiał" birthdate="1960-05-29" gender="F" nation="POL" license="506306600054" swrid="5352178" athleteid="2350">
              <RESULTS>
                <RESULT eventid="1188" points="50" reactiontime="+106" swimtime="00:05:30.06" resultid="2351" heatid="2870" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.69" />
                    <SPLIT distance="100" swimtime="00:02:26.83" />
                    <SPLIT distance="150" swimtime="00:03:57.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" status="DNS" swimtime="00:00:00.00" resultid="2352" heatid="2878" lane="3" />
                <RESULT eventid="1334" points="57" swimtime="00:02:23.98" resultid="2353" heatid="2900" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="82" reactiontime="+101" swimtime="00:01:02.03" resultid="2354" heatid="2905" lane="7" entrytime="00:01:03.81" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulina" lastname="Bielańska-Bugiel" birthdate="1984-04-20" gender="F" nation="POL" license="506306600072" swrid="5468078" athleteid="2321">
              <RESULTS>
                <RESULT eventid="1124" points="96" reactiontime="+126" swimtime="00:01:03.79" resultid="2322" heatid="2851" lane="4" />
                <RESULT eventid="1220" points="104" swimtime="00:04:54.59" resultid="2323" heatid="2873" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.20" />
                    <SPLIT distance="100" swimtime="00:02:26.89" />
                    <SPLIT distance="150" swimtime="00:03:41.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="97" swimtime="00:00:51.47" resultid="2324" heatid="2886" lane="8" />
                <RESULT eventid="1366" points="104" reactiontime="+127" swimtime="00:00:57.34" resultid="2325" heatid="2905" lane="5" entrytime="00:00:53.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Macierzewska" birthdate="1960-04-20" gender="F" nation="POL" license="506306600048" swrid="4992827" athleteid="2341">
              <RESULTS>
                <RESULT eventid="1156" points="264" reactiontime="+90" swimtime="00:01:20.51" resultid="2342" heatid="2861" lane="3" entrytime="00:01:20.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="235" reactiontime="+82" swimtime="00:03:24.34" resultid="2343" heatid="2879" lane="3" entrytime="00:03:18.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.41" />
                    <SPLIT distance="100" swimtime="00:01:36.70" />
                    <SPLIT distance="150" swimtime="00:02:38.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="196" swimtime="00:01:35.45" resultid="2344" heatid="2900" lane="2" entrytime="00:01:32.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1430" points="241" reactiontime="+98" swimtime="00:03:01.45" resultid="2345" heatid="2919" lane="0" entrytime="00:02:55.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.76" />
                    <SPLIT distance="100" swimtime="00:01:27.40" />
                    <SPLIT distance="150" swimtime="00:02:15.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bogusław" lastname="Kwiatkowski" birthdate="1956-07-24" gender="M" nation="POL" license="506306700044" swrid="5468084" athleteid="2311">
              <RESULTS>
                <RESULT eventid="1108" points="58" reactiontime="+97" swimtime="00:02:13.85" resultid="2312" heatid="2847" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="43" reactiontime="+111" swimtime="00:05:59.36" resultid="2313" heatid="2876" lane="6" entrytime="00:05:54.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.77" />
                    <SPLIT distance="100" swimtime="00:02:52.21" />
                    <SPLIT distance="150" swimtime="00:04:25.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="74" reactiontime="+108" swimtime="00:00:49.71" resultid="2314" heatid="2893" lane="1" entrytime="00:00:52.70" entrycourse="LCM" />
                <RESULT eventid="1478" points="53" reactiontime="+103" swimtime="00:04:57.70" resultid="2315" heatid="2929" lane="8" entrytime="00:05:05.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.71" />
                    <SPLIT distance="100" swimtime="00:02:23.81" />
                    <SPLIT distance="150" swimtime="00:03:41.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Janusz" lastname="Toporski" birthdate="1959-10-20" gender="M" nation="POL" license="506306700060" swrid="5484421" athleteid="2292">
              <RESULTS>
                <RESULT eventid="1076" points="131" reactiontime="+82" swimtime="00:00:43.77" resultid="2293" heatid="2840" lane="1" />
                <RESULT eventid="1204" points="96" reactiontime="+90" swimtime="00:04:01.55" resultid="2294" heatid="2871" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.80" />
                    <SPLIT distance="100" swimtime="00:01:54.71" />
                    <SPLIT distance="150" swimtime="00:02:57.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="92" reactiontime="+98" swimtime="00:01:49.17" resultid="2295" heatid="2901" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1414" points="157" reactiontime="+98" swimtime="00:01:45.32" resultid="2296" heatid="2913" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1284" reactiontime="+81" swimtime="00:02:08.70" resultid="2355" heatid="3969" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.26" />
                    <SPLIT distance="100" swimtime="00:01:06.67" />
                    <SPLIT distance="150" swimtime="00:01:33.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2272" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="2341" number="2" />
                    <RELAYPOSITION athleteid="2282" number="3" reactiontime="+23" />
                    <RELAYPOSITION athleteid="2297" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1494" reactiontime="+74" swimtime="00:02:16.88" resultid="2357" heatid="3988" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.52" />
                    <SPLIT distance="100" swimtime="00:01:14.53" />
                    <SPLIT distance="150" swimtime="00:01:48.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2302" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="2287" number="2" />
                    <RELAYPOSITION athleteid="2277" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="2346" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1284" reactiontime="+98" swimtime="00:02:03.55" resultid="2356" heatid="3970" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.65" />
                    <SPLIT distance="100" swimtime="00:01:02.35" />
                    <SPLIT distance="150" swimtime="00:01:35.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2287" number="1" reactiontime="+98" />
                    <RELAYPOSITION athleteid="2302" number="2" />
                    <RELAYPOSITION athleteid="2277" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="2346" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1494" reactiontime="+97" swimtime="00:02:27.60" resultid="2358" heatid="3987" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.73" />
                    <SPLIT distance="100" swimtime="00:01:22.05" />
                    <SPLIT distance="150" swimtime="00:01:50.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2341" number="1" reactiontime="+97" />
                    <RELAYPOSITION athleteid="2272" number="2" />
                    <RELAYPOSITION athleteid="2282" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="2297" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02016" nation="POL" region="16" clubid="2232" name="Koszalińskie TKKF">
          <ATHLETES>
            <ATHLETE firstname="Roman" lastname="Pieślak" birthdate="1979-02-28" gender="M" nation="POL" license="102016700010" swrid="5506636" athleteid="2238">
              <RESULTS>
                <RESULT eventid="1140" points="354" reactiontime="+74" swimtime="00:00:36.66" resultid="2239" heatid="2858" lane="0" entrytime="00:00:36.50" />
                <RESULT eventid="1236" points="325" reactiontime="+83" swimtime="00:03:03.38" resultid="2240" heatid="2877" lane="3" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.90" />
                    <SPLIT distance="100" swimtime="00:01:27.10" />
                    <SPLIT distance="150" swimtime="00:02:14.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1414" points="327" reactiontime="+75" swimtime="00:01:22.56" resultid="2241" heatid="2915" lane="5" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="330" reactiontime="+83" swimtime="00:02:27.60" resultid="2242" heatid="2925" lane="8" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.65" />
                    <SPLIT distance="150" swimtime="00:01:49.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artur" lastname="Mamrot" birthdate="1972-12-10" gender="M" nation="POL" license="102016700007" swrid="5471728" athleteid="2243">
              <RESULTS>
                <RESULT eventid="1140" points="250" reactiontime="+82" swimtime="00:00:41.15" resultid="2244" heatid="2857" lane="1" entrytime="00:00:44.48" entrycourse="LCM" />
                <RESULT eventid="1236" points="229" reactiontime="+95" swimtime="00:03:25.93" resultid="2245" heatid="2877" lane="8" entrytime="00:03:21.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.67" />
                    <SPLIT distance="100" swimtime="00:01:33.82" />
                    <SPLIT distance="150" swimtime="00:02:28.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="231" reactiontime="+91" swimtime="00:00:34.07" resultid="2246" heatid="2894" lane="4" entrytime="00:00:35.01" entrycourse="LCM" />
                <RESULT eventid="1414" points="228" reactiontime="+84" swimtime="00:01:33.10" resultid="2247" heatid="2914" lane="5" entrytime="00:01:41.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Paziewska" birthdate="1974-09-05" gender="F" nation="POL" license="102016600012" swrid="5471732" athleteid="2233">
              <RESULTS>
                <RESULT eventid="1124" points="195" reactiontime="+102" swimtime="00:00:50.46" resultid="2234" heatid="2853" lane="8" entrytime="00:00:45.00" />
                <RESULT eventid="1156" status="DNS" swimtime="00:00:00.00" resultid="2235" heatid="2862" lane="0" entrytime="00:01:16.53" entrycourse="LCM" />
                <RESULT eventid="1301" points="318" reactiontime="+94" swimtime="00:00:34.66" resultid="2236" heatid="2888" lane="2" entrytime="00:00:34.68" entrycourse="LCM" />
                <RESULT eventid="1430" points="257" reactiontime="+98" swimtime="00:02:57.49" resultid="2237" heatid="2919" lane="8" entrytime="00:02:54.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.43" />
                    <SPLIT distance="100" swimtime="00:01:23.14" />
                    <SPLIT distance="150" swimtime="00:02:10.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lidia" lastname="Mikołajczyk" birthdate="1987-04-29" gender="F" nation="POL" license="102016600013" swrid="5471730" athleteid="2253">
              <RESULTS>
                <RESULT eventid="1156" points="408" reactiontime="+95" swimtime="00:01:09.69" resultid="2254" heatid="2862" lane="8" entrytime="00:01:14.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="332" reactiontime="+99" swimtime="00:03:02.12" resultid="2255" heatid="2879" lane="5" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                    <SPLIT distance="100" swimtime="00:01:24.95" />
                    <SPLIT distance="150" swimtime="00:02:17.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="424" reactiontime="+94" swimtime="00:00:31.49" resultid="2256" heatid="2888" lane="5" entrytime="00:00:33.96" entrycourse="LCM" />
                <RESULT eventid="1398" points="341" reactiontime="+97" swimtime="00:01:31.77" resultid="2257" heatid="2912" lane="7" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marian" lastname="Lasowy" birthdate="1955-07-15" gender="M" nation="POL" license="502016700001" swrid="4967127" athleteid="2248">
              <RESULTS>
                <RESULT eventid="1140" status="DNS" swimtime="00:00:00.00" resultid="2249" heatid="2856" lane="3" entrytime="00:00:50.50" />
                <RESULT eventid="1172" status="DNS" swimtime="00:00:00.00" resultid="2250" heatid="2863" lane="3" />
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="2251" heatid="2894" lane="0" entrytime="00:00:41.00" />
                <RESULT eventid="1446" status="DNS" swimtime="00:00:00.00" resultid="2252" heatid="2923" lane="0" entrytime="00:03:29.71" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1284" reactiontime="+80" swimtime="00:02:08.43" resultid="2258" heatid="3970" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.18" />
                    <SPLIT distance="100" swimtime="00:01:01.89" />
                    <SPLIT distance="150" swimtime="00:01:34.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2238" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="2253" number="2" />
                    <RELAYPOSITION athleteid="2243" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="2233" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1494" reactiontime="+91" swimtime="00:02:29.95" resultid="2259" heatid="3988" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.25" />
                    <SPLIT distance="100" swimtime="00:01:19.74" />
                    <SPLIT distance="150" swimtime="00:01:56.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2243" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="2238" number="2" />
                    <RELAYPOSITION athleteid="2253" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="2233" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="1534" name="Niezrzeszeni">
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Fajdasz" birthdate="1973-01-14" gender="M" nation="POL" swrid="4992689" athleteid="2068">
              <RESULTS>
                <RESULT eventid="1108" points="223" reactiontime="+84" swimtime="00:01:25.43" resultid="2069" heatid="2849" lane="6" entrytime="00:01:23.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="281" reactiontime="+80" swimtime="00:01:11.56" resultid="2070" heatid="2868" lane="8" entrytime="00:01:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1382" points="216" reactiontime="+84" swimtime="00:00:39.62" resultid="2071" heatid="2909" lane="3" entrytime="00:00:41.05" />
                <RESULT eventid="1478" points="207" reactiontime="+89" swimtime="00:03:08.98" resultid="2072" heatid="2930" lane="7" entrytime="00:02:50.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.18" />
                    <SPLIT distance="150" swimtime="00:02:20.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Kuśmider" birthdate="1989-01-01" gender="M" nation="POL" athleteid="2047">
              <RESULTS>
                <RESULT eventid="1172" points="383" reactiontime="+86" swimtime="00:01:04.55" resultid="2048" heatid="2867" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="361" reactiontime="+81" swimtime="00:00:29.34" resultid="2049" heatid="2896" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1446" points="339" reactiontime="+89" swimtime="00:02:26.24" resultid="2050" heatid="2924" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                    <SPLIT distance="100" swimtime="00:01:11.35" />
                    <SPLIT distance="150" swimtime="00:01:49.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabela" lastname="Pietrusińska" birthdate="1970-01-01" gender="F" nation="POL" athleteid="1545">
              <RESULTS>
                <RESULT eventid="1059" points="88" swimtime="00:00:54.86" resultid="1546" heatid="2837" lane="1" entrytime="00:00:47.00" />
                <RESULT eventid="1156" points="108" reactiontime="+120" swimtime="00:01:48.34" resultid="1547" heatid="2860" lane="6" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="138" reactiontime="+111" swimtime="00:00:45.75" resultid="1548" heatid="2887" lane="6" entrytime="00:00:45.00" />
                <RESULT eventid="1430" points="105" reactiontime="+104" swimtime="00:03:58.73" resultid="1549" heatid="2918" lane="2" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.26" />
                    <SPLIT distance="100" swimtime="00:01:54.40" />
                    <SPLIT distance="150" swimtime="00:02:59.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Boruch" birthdate="1978-08-25" gender="F" nation="POL" athleteid="1859">
              <RESULTS>
                <RESULT eventid="1059" points="190" reactiontime="+80" swimtime="00:00:42.43" resultid="1860" heatid="2837" lane="8" entrytime="00:00:50.00" />
                <RESULT eventid="1156" points="218" reactiontime="+89" swimtime="00:01:25.80" resultid="1861" heatid="2861" lane="8" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="104" swimtime="00:01:57.95" resultid="1862" heatid="2900" lane="7" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robert" lastname="Brus" birthdate="1967-04-30" gender="M" nation="POL" swrid="4218696" athleteid="1863">
              <RESULTS>
                <RESULT eventid="1140" points="183" swimtime="00:00:45.63" resultid="1864" heatid="2857" lane="9" entrytime="00:00:48.00" />
                <RESULT eventid="1382" points="212" reactiontime="+80" swimtime="00:00:39.91" resultid="1865" heatid="2909" lane="4" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Olborski" birthdate="1997-09-06" gender="M" nation="POL" swrid="4261737" athleteid="1572">
              <RESULTS>
                <RESULT eventid="1076" points="614" reactiontime="+73" swimtime="00:00:26.20" resultid="1573" heatid="2844" lane="6" entrytime="00:00:27.00" />
                <RESULT eventid="1172" points="571" reactiontime="+77" swimtime="00:00:56.52" resultid="1574" heatid="2869" lane="5" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Kopeć" birthdate="1978-01-01" gender="M" nation="POL" athleteid="2036">
              <RESULTS>
                <RESULT eventid="1076" points="103" reactiontime="+82" swimtime="00:00:47.37" resultid="2037" heatid="2842" lane="6" entrytime="00:00:40.00" />
                <RESULT eventid="1172" points="159" reactiontime="+73" swimtime="00:01:26.48" resultid="2038" heatid="2866" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="209" reactiontime="+78" swimtime="00:00:35.19" resultid="2039" heatid="2895" lane="5" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Demczuk" birthdate="1982-06-15" gender="M" nation="POL" athleteid="2025">
              <RESULTS>
                <RESULT eventid="1172" points="225" reactiontime="+85" swimtime="00:01:17.03" resultid="2026" heatid="2866" lane="3" entrytime="00:01:22.00" />
                <RESULT eventid="1318" points="272" reactiontime="+84" swimtime="00:00:32.25" resultid="2027" heatid="2895" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="1446" points="169" reactiontime="+89" swimtime="00:03:04.42" resultid="2028" heatid="2923" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.62" />
                    <SPLIT distance="100" swimtime="00:01:27.92" />
                    <SPLIT distance="150" swimtime="00:02:16.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartłomiej" lastname="Lassek" birthdate="1994-01-01" gender="M" nation="POL" swrid="4181299" athleteid="2051">
              <RESULTS>
                <RESULT eventid="1076" points="696" reactiontime="+74" swimtime="00:00:25.12" resultid="2052" heatid="2844" lane="4" entrytime="00:00:24.50" />
                <RESULT comment="Rekord Polski Masters" eventid="1446" points="660" reactiontime="+74" swimtime="00:01:57.15" resultid="2053" heatid="2925" lane="4" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.21" />
                    <SPLIT distance="100" swimtime="00:00:56.93" />
                    <SPLIT distance="150" swimtime="00:01:27.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Grzelczak" birthdate="1985-01-11" gender="M" nation="POL" athleteid="1535">
              <RESULTS>
                <RESULT eventid="1140" points="245" reactiontime="+98" swimtime="00:00:41.44" resultid="1536" heatid="2857" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="1236" points="201" reactiontime="+98" swimtime="00:03:34.96" resultid="1537" heatid="2877" lane="9" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.16" />
                    <SPLIT distance="100" swimtime="00:01:40.86" />
                    <SPLIT distance="150" swimtime="00:02:38.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1414" points="202" reactiontime="+106" swimtime="00:01:36.80" resultid="1538" heatid="2915" lane="8" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="117" reactiontime="+108" swimtime="00:03:27.98" resultid="1539" heatid="2923" lane="2" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.03" />
                    <SPLIT distance="100" swimtime="00:01:36.48" />
                    <SPLIT distance="150" swimtime="00:02:33.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Gołębiowski" birthdate="1996-05-20" gender="M" nation="POL" swrid="4115580" athleteid="1698">
              <RESULTS>
                <RESULT eventid="1140" points="411" reactiontime="+67" swimtime="00:00:34.88" resultid="1699" heatid="2858" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="1318" points="452" reactiontime="+67" swimtime="00:00:27.23" resultid="1700" heatid="2896" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="1414" points="370" reactiontime="+71" swimtime="00:01:19.19" resultid="1701" heatid="2916" lane="3" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="455" reactiontime="+71" swimtime="00:01:00.96" resultid="1702" heatid="2867" lane="5" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sławomir" lastname="Formas" birthdate="1969-11-05" gender="M" nation="POL" swrid="4292540" athleteid="1603">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1140" points="512" reactiontime="+77" swimtime="00:00:32.43" resultid="1604" heatid="2858" lane="7" entrytime="00:00:33.00" />
                <RESULT comment="Rekord Polski Masters" eventid="1236" points="479" reactiontime="+86" swimtime="00:02:41.10" resultid="1605" heatid="2877" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.90" />
                    <SPLIT distance="100" swimtime="00:01:17.06" />
                    <SPLIT distance="150" swimtime="00:01:59.18" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1414" points="494" reactiontime="+79" swimtime="00:01:11.93" resultid="1606" heatid="2916" lane="7" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robert" lastname="Pietrusiński" birthdate="1962-01-01" gender="M" nation="POL" athleteid="1550">
              <RESULTS>
                <RESULT eventid="1076" points="176" reactiontime="+94" swimtime="00:00:39.67" resultid="1551" heatid="2842" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1268" points="129" reactiontime="+102" swimtime="00:03:45.40" resultid="1552" heatid="2883" lane="9" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.66" />
                    <SPLIT distance="100" swimtime="00:01:43.25" />
                    <SPLIT distance="150" swimtime="00:02:54.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="187" reactiontime="+111" swimtime="00:00:36.52" resultid="1553" heatid="2895" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="1382" points="182" reactiontime="+83" swimtime="00:00:41.97" resultid="1554" heatid="2910" lane="9" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Roksela" birthdate="1981-01-01" gender="M" nation="POL" athleteid="2044">
              <RESULTS>
                <RESULT eventid="1076" points="123" reactiontime="+81" swimtime="00:00:44.73" resultid="2045" heatid="2842" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1172" points="176" reactiontime="+100" swimtime="00:01:23.59" resultid="2046" heatid="2866" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krystian" lastname="Bator" birthdate="1981-03-09" gender="M" nation="POL" swrid="5394192" athleteid="1591">
              <RESULTS>
                <RESULT eventid="1076" points="425" reactiontime="+70" swimtime="00:00:29.62" resultid="1592" heatid="2844" lane="0" entrytime="00:00:29.00" />
                <RESULT eventid="1172" points="415" reactiontime="+71" swimtime="00:01:02.88" resultid="1593" heatid="2869" lane="8" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="399" reactiontime="+68" swimtime="00:00:28.39" resultid="1594" heatid="2897" lane="6" entrytime="00:00:27.49" />
                <RESULT eventid="1350" points="279" reactiontime="+77" swimtime="00:01:15.62" resultid="1595" heatid="2903" lane="8" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Woźniak" birthdate="1986-08-22" gender="M" nation="POL" athleteid="1583">
              <RESULTS>
                <RESULT eventid="1140" points="95" reactiontime="+112" swimtime="00:00:56.82" resultid="1584" heatid="2856" lane="7" entrytime="00:00:57.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dorota" lastname="Bartniak" birthdate="1997-01-01" gender="F" nation="POL" swrid="4287745" athleteid="2054">
              <RESULTS>
                <RESULT eventid="1156" points="445" reactiontime="+78" swimtime="00:01:07.71" resultid="2055" heatid="2862" lane="9" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="426" reactiontime="+77" swimtime="00:02:47.55" resultid="2056" heatid="2879" lane="4" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                    <SPLIT distance="100" swimtime="00:01:18.60" />
                    <SPLIT distance="150" swimtime="00:02:05.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1430" points="358" reactiontime="+85" swimtime="00:02:39.00" resultid="2057" heatid="2919" lane="9" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.78" />
                    <SPLIT distance="100" swimtime="00:01:18.83" />
                    <SPLIT distance="150" swimtime="00:02:00.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1398" points="450" reactiontime="+82" swimtime="00:01:23.68" resultid="2058" heatid="2912" lane="5" entrytime="00:01:21.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jarosław" lastname="Guziński" birthdate="1966-01-01" gender="M" nation="POL" swrid="5484405" athleteid="1611">
              <RESULTS>
                <RESULT eventid="1076" points="146" reactiontime="+98" swimtime="00:00:42.20" resultid="1612" heatid="2840" lane="2" />
                <RESULT eventid="1172" points="171" reactiontime="+91" swimtime="00:01:24.49" resultid="1613" heatid="2864" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="1614" heatid="2892" lane="0" />
                <RESULT eventid="1350" status="DNS" swimtime="00:00:00.00" resultid="1615" heatid="2902" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jarek" lastname="Kopeć" birthdate="1969-01-01" gender="M" nation="POL" athleteid="2032">
              <RESULTS>
                <RESULT eventid="1172" points="209" reactiontime="+89" swimtime="00:01:18.97" resultid="2033" heatid="2866" lane="5" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="245" reactiontime="+97" swimtime="00:00:33.39" resultid="2034" heatid="2895" lane="7" entrytime="00:00:34.00" />
                <RESULT eventid="1446" points="177" reactiontime="+89" swimtime="00:03:01.53" resultid="2035" heatid="2924" lane="9" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.67" />
                    <SPLIT distance="100" swimtime="00:01:23.01" />
                    <SPLIT distance="150" swimtime="00:02:11.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Kędzior" birthdate="1973-12-08" gender="M" nation="POL" athleteid="1797">
              <RESULTS>
                <RESULT eventid="1108" points="177" reactiontime="+79" swimtime="00:01:32.27" resultid="1798" heatid="2849" lane="7" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="252" reactiontime="+95" swimtime="00:01:14.19" resultid="1799" heatid="2867" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="250" reactiontime="+89" swimtime="00:00:33.18" resultid="1800" heatid="2895" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="1478" points="145" reactiontime="+91" swimtime="00:03:32.90" resultid="1801" heatid="2929" lane="5" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.77" />
                    <SPLIT distance="100" swimtime="00:01:43.20" />
                    <SPLIT distance="150" swimtime="00:02:40.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Janczewski" birthdate="1990-12-06" gender="M" nation="POL" athleteid="1994">
              <RESULTS>
                <RESULT eventid="1318" points="582" reactiontime="+82" swimtime="00:00:25.04" resultid="1995" heatid="2898" lane="6" entrytime="00:00:26.00" />
                <RESULT eventid="1446" points="519" reactiontime="+89" swimtime="00:02:06.90" resultid="1996" heatid="2925" lane="2" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.94" />
                    <SPLIT distance="100" swimtime="00:01:02.33" />
                    <SPLIT distance="150" swimtime="00:01:34.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Syska" birthdate="2002-03-05" gender="M" nation="POL" swrid="4852151" athleteid="1787">
              <RESULTS>
                <RESULT eventid="1076" points="512" reactiontime="+63" swimtime="00:00:27.83" resultid="1788" heatid="2844" lane="3" entrytime="00:00:27.00" />
                <RESULT eventid="1318" points="473" reactiontime="+65" swimtime="00:00:26.82" resultid="1789" heatid="2898" lane="7" entrytime="00:00:26.00" />
                <RESULT eventid="1172" points="496" reactiontime="+63" swimtime="00:00:59.25" resultid="1790" heatid="2869" lane="2" entrytime="00:00:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="492" reactiontime="+66" swimtime="00:01:02.63" resultid="1791" heatid="2903" lane="4" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabela" lastname="Wypych-Staszewska" birthdate="1970-01-01" gender="F" nation="POL" athleteid="1575">
              <RESULTS>
                <RESULT eventid="1059" points="211" reactiontime="+67" swimtime="00:00:41.01" resultid="1576" heatid="2837" lane="7" entrytime="00:00:42.00" />
                <RESULT eventid="1156" points="246" reactiontime="+66" swimtime="00:01:22.51" resultid="1577" heatid="2860" lane="5" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="227" reactiontime="+75" swimtime="00:00:38.76" resultid="1578" heatid="2888" lane="9" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Kubiak" birthdate="1989-07-05" gender="M" nation="POL" athleteid="1792">
              <RESULTS>
                <RESULT eventid="1204" points="139" swimtime="00:03:33.70" resultid="1793" heatid="2872" lane="6" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.59" />
                    <SPLIT distance="100" swimtime="00:01:41.43" />
                    <SPLIT distance="150" swimtime="00:02:38.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="133" swimtime="00:04:06.54" resultid="1794" heatid="2876" lane="5" entrytime="00:04:00.00" />
                <RESULT eventid="1350" points="121" swimtime="00:01:39.77" resultid="1795" heatid="2902" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1478" points="116" reactiontime="+96" swimtime="00:03:49.28" resultid="1796" heatid="2929" lane="7" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.30" />
                    <SPLIT distance="100" swimtime="00:01:54.34" />
                    <SPLIT distance="150" swimtime="00:02:53.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artur" lastname="Malina" birthdate="1970-02-10" gender="M" nation="POL" athleteid="2100">
              <RESULTS>
                <RESULT eventid="1140" status="DNS" swimtime="00:00:00.00" resultid="2101" heatid="2856" lane="4" entrytime="00:00:49.00" />
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="2102" heatid="2893" lane="4" entrytime="00:00:42.00" />
                <RESULT eventid="1236" status="DNS" swimtime="00:00:00.00" resultid="2103" heatid="2876" lane="3" entrytime="00:05:00.00" />
                <RESULT eventid="1414" status="DNS" swimtime="00:00:00.00" resultid="2104" heatid="2916" lane="4" entrytime="00:00:54.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Bartoszewski" birthdate="1994-03-09" gender="M" nation="POL" swrid="4181340" athleteid="2126">
              <RESULTS>
                <RESULT eventid="1140" points="525" reactiontime="+78" swimtime="00:00:32.15" resultid="2127" heatid="2858" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="1318" points="531" reactiontime="+69" swimtime="00:00:25.81" resultid="2128" heatid="2898" lane="2" entrytime="00:00:26.00" />
                <RESULT eventid="1382" points="508" reactiontime="+64" swimtime="00:00:29.82" resultid="2129" heatid="2910" lane="5" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Wypych" birthdate="1991-01-01" gender="M" nation="POL" swrid="4072458" athleteid="2029">
              <RESULTS>
                <RESULT eventid="1140" points="657" reactiontime="+71" swimtime="00:00:29.85" resultid="2030" heatid="2858" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1318" points="699" reactiontime="+67" swimtime="00:00:23.55" resultid="2031" heatid="2898" lane="4" entrytime="00:00:24.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Kotulski" birthdate="1981-01-01" gender="M" nation="POL" athleteid="2040">
              <RESULTS>
                <RESULT eventid="1076" points="262" reactiontime="+87" swimtime="00:00:34.76" resultid="2041" heatid="2842" lane="5" entrytime="00:00:37.00" />
                <RESULT eventid="1172" points="213" reactiontime="+87" swimtime="00:01:18.48" resultid="2042" heatid="2867" lane="9" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="232" reactiontime="+81" swimtime="00:00:33.99" resultid="2043" heatid="2895" lane="4" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Zieliński" birthdate="2000-06-03" gender="M" nation="POL" swrid="4639122" athleteid="1607">
              <RESULTS>
                <RESULT eventid="1140" points="340" reactiontime="+78" swimtime="00:00:37.17" resultid="1608" heatid="2856" lane="9" />
                <RESULT eventid="1414" points="287" reactiontime="+86" swimtime="00:01:26.17" resultid="1609" heatid="2914" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="412" reactiontime="+81" swimtime="00:00:28.08" resultid="1610" heatid="2893" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Łopuszyński" birthdate="1969-11-10" gender="M" nation="POL" athleteid="1540">
              <RESULTS>
                <RESULT eventid="1204" points="96" reactiontime="+113" swimtime="00:04:01.65" resultid="1541" heatid="2872" lane="7" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.34" />
                    <SPLIT distance="100" swimtime="00:01:51.66" />
                    <SPLIT distance="150" swimtime="00:02:56.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="99" reactiontime="+110" swimtime="00:04:05.88" resultid="1542" heatid="2882" lane="3" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.55" />
                    <SPLIT distance="100" swimtime="00:02:00.90" />
                    <SPLIT distance="150" swimtime="00:03:08.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="110" reactiontime="+112" swimtime="00:00:43.59" resultid="1543" heatid="2893" lane="6" entrytime="00:00:45.00" />
                <RESULT eventid="1350" points="90" reactiontime="+106" swimtime="00:01:50.12" resultid="1544" heatid="2902" lane="6" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Zrobek" birthdate="1999-11-10" gender="F" nation="POL" swrid="4493371" athleteid="2109">
              <RESULTS>
                <RESULT eventid="1059" points="513" reactiontime="+77" swimtime="00:00:30.50" resultid="2110" heatid="2838" lane="4" entrytime="00:00:30.80" />
                <RESULT eventid="1156" points="609" reactiontime="+76" swimtime="00:01:00.99" resultid="2111" heatid="2862" lane="5" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="604" reactiontime="+74" swimtime="00:00:27.99" resultid="2112" heatid="2889" lane="5" entrytime="00:00:27.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Bogusiak" birthdate="1982-05-30" gender="M" nation="POL" athleteid="2832">
              <RESULTS>
                <RESULT eventid="1318" points="215" reactiontime="+95" swimtime="00:00:34.90" resultid="2833" heatid="2895" lane="0" entrytime="00:00:34.50" />
                <RESULT eventid="1172" points="212" reactiontime="+78" swimtime="00:01:18.60" resultid="2834" heatid="2866" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="180" reactiontime="+97" swimtime="00:03:00.60" resultid="2835" heatid="2923" lane="3" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.98" />
                    <SPLIT distance="150" swimtime="00:02:14.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Malicki" birthdate="1984-02-12" gender="M" nation="POL" athleteid="1730">
              <RESULTS>
                <RESULT eventid="1172" points="381" reactiontime="+97" swimtime="00:01:04.69" resultid="1731" heatid="2868" lane="1" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="379" reactiontime="+95" swimtime="00:00:28.88" resultid="1732" heatid="2897" lane="7" entrytime="00:00:28.00" />
                <RESULT eventid="1268" points="268" reactiontime="+94" swimtime="00:02:56.78" resultid="1733" heatid="2883" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.04" />
                    <SPLIT distance="100" swimtime="00:01:21.03" />
                    <SPLIT distance="150" swimtime="00:02:15.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="311" reactiontime="+95" swimtime="00:02:30.54" resultid="1734" heatid="2925" lane="7" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                    <SPLIT distance="100" swimtime="00:01:09.98" />
                    <SPLIT distance="150" swimtime="00:01:50.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Pawiński" birthdate="1984-01-01" gender="M" nation="POL" athleteid="2059">
              <RESULTS>
                <RESULT eventid="1318" points="276" reactiontime="+79" swimtime="00:00:32.11" resultid="2060" heatid="2896" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="1446" status="DNS" swimtime="00:00:00.00" resultid="2061" heatid="2924" lane="8" entrytime="00:02:50.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="1928" name="MUKS Zgierz">
          <ATHLETES>
            <ATHLETE firstname="Robert" lastname="Szalbierz" birthdate="1968-08-06" gender="M" nation="POL" license="502805700034" swrid="5373990" athleteid="2524">
              <RESULTS>
                <RESULT eventid="1076" points="288" reactiontime="+92" swimtime="00:00:33.69" resultid="2525" heatid="2840" lane="7" />
                <RESULT eventid="1172" points="284" reactiontime="+89" swimtime="00:01:11.34" resultid="2526" heatid="2865" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="305" reactiontime="+91" swimtime="00:00:31.05" resultid="2527" heatid="2891" lane="6" />
                <RESULT eventid="1446" points="247" reactiontime="+97" swimtime="00:02:42.37" resultid="2528" heatid="2921" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                    <SPLIT distance="100" swimtime="00:01:18.24" />
                    <SPLIT distance="150" swimtime="00:02:00.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Jasiński" birthdate="1969-01-02" gender="M" nation="POL" athleteid="2086">
              <RESULTS>
                <RESULT eventid="1172" points="134" reactiontime="+111" swimtime="00:01:31.57" resultid="2087" heatid="2866" lane="0" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="2088" heatid="2894" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1446" status="DNS" swimtime="00:00:00.00" resultid="2089" heatid="2923" lane="9" entrytime="00:03:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zdzisław" lastname="Jasiński" birthdate="1960-07-23" gender="M" nation="POL" license="502805700027" swrid="5374015" athleteid="2579">
              <RESULTS>
                <RESULT eventid="1172" points="212" reactiontime="+84" swimtime="00:01:18.55" resultid="2580" heatid="2863" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="177" reactiontime="+122" swimtime="00:03:44.58" resultid="2581" heatid="2875" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.49" />
                    <SPLIT distance="100" swimtime="00:01:47.59" />
                    <SPLIT distance="150" swimtime="00:02:46.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="199" reactiontime="+89" swimtime="00:00:35.80" resultid="2582" heatid="2890" lane="3" />
                <RESULT eventid="1446" points="126" reactiontime="+116" swimtime="00:03:23.20" resultid="2583" heatid="2920" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                    <SPLIT distance="100" swimtime="00:01:30.87" />
                    <SPLIT distance="150" swimtime="00:02:26.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Rembowska-Świeboda" birthdate="1968-06-27" gender="F" nation="POL" athleteid="2827">
              <RESULTS>
                <RESULT eventid="1301" points="345" reactiontime="+76" swimtime="00:00:33.74" resultid="2828" heatid="2888" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1366" points="308" reactiontime="+77" swimtime="00:00:39.92" resultid="2829" heatid="2906" lane="1" entrytime="00:00:39.00" />
                <RESULT eventid="1156" points="287" reactiontime="+81" swimtime="00:01:18.36" resultid="2830" heatid="2861" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="289" reactiontime="+70" swimtime="00:01:26.88" resultid="2831" heatid="2846" lane="8" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Węgrzycka" birthdate="1977-01-26" gender="F" nation="POL" license="502805600056" swrid="5464095" athleteid="2570">
              <RESULTS>
                <RESULT eventid="1156" points="138" reactiontime="+101" swimtime="00:01:40.06" resultid="2571" heatid="2860" lane="3" entrytime="00:01:39.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="156" reactiontime="+94" swimtime="00:00:43.97" resultid="2572" heatid="2887" lane="3" entrytime="00:00:43.22" entrycourse="LCM" />
                <RESULT eventid="1430" points="121" reactiontime="+117" swimtime="00:03:47.91" resultid="2573" heatid="2917" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.79" />
                    <SPLIT distance="100" swimtime="00:01:44.83" />
                    <SPLIT distance="150" swimtime="00:02:46.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Justyna" lastname="Barańska" birthdate="1984-02-23" gender="F" nation="POL" license="102805600050" athleteid="2565">
              <RESULTS>
                <RESULT eventid="1156" points="265" reactiontime="+87" swimtime="00:01:20.46" resultid="2566" heatid="2859" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1220" points="271" reactiontime="+86" swimtime="00:03:34.50" resultid="2567" heatid="2873" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.01" />
                    <SPLIT distance="100" swimtime="00:01:42.60" />
                    <SPLIT distance="150" swimtime="00:02:38.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1398" points="262" reactiontime="+104" swimtime="00:01:40.11" resultid="2568" heatid="2911" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1430" points="235" reactiontime="+89" swimtime="00:03:02.99" resultid="2569" heatid="2917" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.19" />
                    <SPLIT distance="100" swimtime="00:01:26.45" />
                    <SPLIT distance="150" swimtime="00:02:15.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Włodzimierz" lastname="Przytulski" birthdate="1957-01-09" gender="M" nation="POL" license="502805700049" swrid="4754657" athleteid="2516">
              <RESULTS>
                <RESULT eventid="1076" points="290" reactiontime="+93" swimtime="00:00:33.61" resultid="2517" heatid="2839" lane="4" />
                <RESULT eventid="1204" points="167" reactiontime="+104" swimtime="00:03:21.05" resultid="2518" heatid="2871" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.52" />
                    <SPLIT distance="100" swimtime="00:01:37.00" />
                    <SPLIT distance="150" swimtime="00:02:29.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="192" reactiontime="+100" swimtime="00:01:25.64" resultid="2519" heatid="2901" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jarosław" lastname="Woźniak" birthdate="1980-09-30" gender="M" nation="POL" swrid="5506643" athleteid="2082">
              <RESULTS>
                <RESULT eventid="1172" points="150" reactiontime="+100" swimtime="00:01:28.17" resultid="2083" heatid="2866" lane="2" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="215" reactiontime="+110" swimtime="00:00:34.86" resultid="2084" heatid="2894" lane="1" entrytime="00:00:39.00" />
                <RESULT eventid="1414" points="160" reactiontime="+117" swimtime="00:01:44.56" resultid="2085" heatid="2915" lane="9" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roman" lastname="Wiczel" birthdate="1948-01-22" gender="M" nation="POL" license="502805700021" swrid="4876444" athleteid="2597">
              <RESULTS>
                <RESULT eventid="1236" points="190" reactiontime="+98" swimtime="00:03:39.35" resultid="2598" heatid="2875" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.79" />
                    <SPLIT distance="100" swimtime="00:01:48.36" />
                    <SPLIT distance="150" swimtime="00:02:46.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1414" points="184" reactiontime="+101" swimtime="00:01:39.86" resultid="2599" heatid="2914" lane="4" entrytime="00:01:40.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="203" reactiontime="+96" swimtime="00:00:44.11" resultid="2758" heatid="2857" lane="7" entrytime="00:00:42.05" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Justyna" lastname="Barańska" birthdate="1977-01-05" gender="F" nation="POL" license="502805600055" swrid="4655158" athleteid="2532">
              <RESULTS>
                <RESULT eventid="1124" points="252" reactiontime="+97" swimtime="00:00:46.38" resultid="2533" heatid="2852" lane="4" entrytime="00:00:47.83" entrycourse="LCM" />
                <RESULT eventid="1220" points="250" reactiontime="+80" swimtime="00:03:40.28" resultid="2534" heatid="2874" lane="5" entrytime="00:03:47.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.67" />
                    <SPLIT distance="100" swimtime="00:01:49.42" />
                    <SPLIT distance="150" swimtime="00:02:46.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1398" points="236" swimtime="00:01:43.72" resultid="2535" heatid="2912" lane="9" entrytime="00:01:46.17" entrycourse="LCM" />
                <RESULT eventid="1462" points="154" swimtime="00:03:50.11" resultid="2536" heatid="2926" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.96" />
                    <SPLIT distance="100" swimtime="00:01:55.81" />
                    <SPLIT distance="150" swimtime="00:02:56.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Morozowski" birthdate="1973-05-09" gender="M" nation="POL" license="102805700051" swrid="5416829" athleteid="2550">
              <RESULTS>
                <RESULT eventid="1140" points="269" reactiontime="+96" swimtime="00:00:40.17" resultid="2551" heatid="2855" lane="1" />
                <RESULT eventid="1236" points="209" swimtime="00:03:32.38" resultid="2552" heatid="2876" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.14" />
                    <SPLIT distance="100" swimtime="00:01:41.24" />
                    <SPLIT distance="150" swimtime="00:02:36.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1414" points="214" reactiontime="+109" swimtime="00:01:35.06" resultid="2553" heatid="2914" lane="9" />
                <RESULT eventid="1446" points="187" reactiontime="+105" swimtime="00:02:58.30" resultid="2554" heatid="2921" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.53" />
                    <SPLIT distance="100" swimtime="00:01:22.41" />
                    <SPLIT distance="150" swimtime="00:02:10.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Piekarski" birthdate="1986-04-22" gender="M" nation="POL" license="502805700144" athleteid="2589">
              <RESULTS>
                <RESULT eventid="1172" points="120" reactiontime="+143" swimtime="00:01:34.91" resultid="2590" heatid="2865" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="160" reactiontime="+100" swimtime="00:00:38.49" resultid="2591" heatid="2891" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Kaczmarek" birthdate="1976-11-27" gender="F" nation="POL" athleteid="2759">
              <RESULTS>
                <RESULT eventid="1124" points="109" swimtime="00:01:01.25" resultid="2760" heatid="2852" lane="5" entrytime="00:00:50.00" />
                <RESULT eventid="1301" status="DNS" swimtime="00:00:00.00" resultid="2761" heatid="2887" lane="4" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Gajda" birthdate="1978-02-23" gender="M" nation="POL" athleteid="2817">
              <RESULTS>
                <RESULT eventid="1318" points="276" reactiontime="+84" swimtime="00:00:32.10" resultid="2818" heatid="2895" lane="1" entrytime="00:00:34.00" />
                <RESULT eventid="1414" points="218" reactiontime="+94" swimtime="00:01:34.41" resultid="2819" heatid="2915" lane="2" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Janusz" lastname="Błasiak" birthdate="1955-03-16" gender="M" nation="POL" license="502805700037" swrid="5464088" athleteid="2584">
              <RESULTS>
                <RESULT eventid="1172" points="106" reactiontime="+89" swimtime="00:01:38.89" resultid="2585" heatid="2863" lane="8" />
                <RESULT eventid="1268" points="59" reactiontime="+97" swimtime="00:04:52.15" resultid="2586" heatid="2882" lane="7" entrytime="00:04:48.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.98" />
                    <SPLIT distance="100" swimtime="00:02:29.87" />
                    <SPLIT distance="150" swimtime="00:03:55.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="107" reactiontime="+93" swimtime="00:00:43.94" resultid="2587" heatid="2890" lane="7" />
                <RESULT eventid="1446" points="87" reactiontime="+98" swimtime="00:03:49.82" resultid="2588" heatid="2922" lane="5" entrytime="00:03:47.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:51.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Włodzimierz" lastname="Łatecki" birthdate="1957-05-25" gender="M" nation="POL" license="502805700022" swrid="5464093" athleteid="2592">
              <RESULTS>
                <RESULT eventid="1204" points="31" swimtime="00:05:49.54" resultid="2593" heatid="2871" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.17" />
                    <SPLIT distance="100" swimtime="00:02:44.84" />
                    <SPLIT distance="150" swimtime="00:04:18.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="40" reactiontime="+119" swimtime="00:05:33.14" resultid="2594" heatid="2880" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.69" />
                    <SPLIT distance="150" swimtime="00:04:28.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="55" reactiontime="+129" swimtime="00:04:27.97" resultid="2595" heatid="2922" lane="6" entrytime="00:04:22.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.66" />
                    <SPLIT distance="150" swimtime="00:03:17.69" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G4" eventid="1478" status="DSQ" swimtime="00:00:00.00" resultid="2596" heatid="2928" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Lis - Piwowarski" birthdate="1984-05-29" gender="M" nation="POL" license="502805700146" swrid="5506632" athleteid="2520">
              <RESULTS>
                <RESULT eventid="1076" points="58" reactiontime="+91" swimtime="00:00:57.48" resultid="2521" heatid="2841" lane="6" />
                <RESULT eventid="1172" points="126" reactiontime="+97" swimtime="00:01:33.41" resultid="2522" heatid="2864" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="175" reactiontime="+85" swimtime="00:00:37.34" resultid="2523" heatid="2892" lane="7" />
                <RESULT eventid="1446" points="79" reactiontime="+104" swimtime="00:03:57.63" resultid="2934" heatid="2920" lane="0" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.24" />
                    <SPLIT distance="100" swimtime="00:01:40.35" />
                    <SPLIT distance="150" swimtime="00:02:46.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Sypniewski" birthdate="1957-02-01" gender="M" nation="POL" license="102805700035" swrid="5373999" athleteid="2555">
              <RESULTS>
                <RESULT eventid="1140" points="236" reactiontime="+74" swimtime="00:00:41.99" resultid="2556" heatid="2854" lane="5" />
                <RESULT eventid="1268" points="158" reactiontime="+82" swimtime="00:03:30.58" resultid="2557" heatid="2880" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.31" />
                    <SPLIT distance="100" swimtime="00:01:44.10" />
                    <SPLIT distance="150" swimtime="00:02:41.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1382" points="210" reactiontime="+77" swimtime="00:00:40.04" resultid="2558" heatid="2907" lane="5" />
                <RESULT eventid="1414" points="188" reactiontime="+78" swimtime="00:01:39.23" resultid="2559" heatid="2913" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Wiśniewska" birthdate="1981-02-26" gender="F" nation="POL" license="502805600123" swrid="5464096" athleteid="2537">
              <RESULTS>
                <RESULT eventid="1124" points="94" reactiontime="+125" swimtime="00:01:04.36" resultid="2538" heatid="2851" lane="2" />
                <RESULT eventid="1220" points="96" reactiontime="+134" swimtime="00:05:02.47" resultid="2539" heatid="2873" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.78" />
                    <SPLIT distance="100" swimtime="00:02:27.01" />
                    <SPLIT distance="150" swimtime="00:03:45.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="82" reactiontime="+136" swimtime="00:00:54.35" resultid="2540" heatid="2886" lane="6" entrytime="00:01:02.85" entrycourse="LCM" />
                <RESULT eventid="1398" points="82" reactiontime="+131" swimtime="00:02:27.45" resultid="2541" heatid="2911" lane="1" entrytime="00:02:19.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daria" lastname="Fajkowska" birthdate="1973-03-18" gender="F" nation="POL" license="502805600044" swrid="4992744" athleteid="2506">
              <RESULTS>
                <RESULT eventid="1059" points="402" reactiontime="+81" swimtime="00:00:33.09" resultid="2507" heatid="2836" lane="2" />
                <RESULT eventid="1124" points="349" reactiontime="+85" swimtime="00:00:41.58" resultid="2508" heatid="2852" lane="9" />
                <RESULT eventid="1301" points="472" reactiontime="+94" swimtime="00:00:30.38" resultid="2509" heatid="2886" lane="7" />
                <RESULT eventid="1366" points="478" reactiontime="+81" swimtime="00:00:34.49" resultid="2510" heatid="2905" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Szczęsnowicz" birthdate="1986-07-27" gender="F" nation="POL" athleteid="2093">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="2094" heatid="2838" lane="9" entrytime="00:00:37.00" />
                <RESULT eventid="1301" status="DNS" swimtime="00:00:00.00" resultid="2095" heatid="2889" lane="0" entrytime="00:00:32.00" />
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="2096" heatid="2853" lane="3" entrytime="00:00:38.00" />
                <RESULT eventid="1398" status="DNS" swimtime="00:00:00.00" resultid="2097" heatid="2912" lane="6" entrytime="00:01:27.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tadeusz" lastname="Obiedziński" birthdate="1959-05-12" gender="M" nation="POL" license="502805700040" swrid="4992722" athleteid="2542">
              <RESULTS>
                <RESULT eventid="1140" points="213" reactiontime="+90" swimtime="00:00:43.40" resultid="2543" heatid="2854" lane="4" />
                <RESULT eventid="1236" points="142" reactiontime="+108" swimtime="00:04:01.23" resultid="2544" heatid="2875" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.22" />
                    <SPLIT distance="100" swimtime="00:01:57.54" />
                    <SPLIT distance="150" swimtime="00:03:02.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1414" points="145" reactiontime="+92" swimtime="00:01:48.08" resultid="2545" heatid="2914" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Bednarek" birthdate="1951-03-24" gender="M" nation="POL" license="502805700052" swrid="5464087" athleteid="2574">
              <RESULTS>
                <RESULT eventid="1172" points="180" reactiontime="+84" swimtime="00:01:23.06" resultid="2575" heatid="2863" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="118" swimtime="00:03:52.33" resultid="2576" heatid="2880" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.89" />
                    <SPLIT distance="100" swimtime="00:01:53.85" />
                    <SPLIT distance="150" swimtime="00:03:02.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="187" swimtime="00:00:36.54" resultid="2577" heatid="2894" lane="2" entrytime="00:00:36.84" entrycourse="LCM" />
                <RESULT eventid="1446" points="147" reactiontime="+120" swimtime="00:03:13.17" resultid="2578" heatid="2920" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.68" />
                    <SPLIT distance="100" swimtime="00:01:31.30" />
                    <SPLIT distance="150" swimtime="00:02:22.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Klusek" birthdate="1975-01-12" gender="F" nation="POL" license="502805600030" swrid="5464092" athleteid="2511">
              <RESULTS>
                <RESULT eventid="1059" points="266" reactiontime="+101" swimtime="00:00:37.96" resultid="2512" heatid="2837" lane="5" entrytime="00:00:37.66" entrycourse="LCM" />
                <RESULT eventid="1188" points="229" reactiontime="+109" swimtime="00:03:19.06" resultid="2513" heatid="2870" lane="5" entrytime="00:03:16.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.29" />
                    <SPLIT distance="100" swimtime="00:01:31.87" />
                    <SPLIT distance="150" swimtime="00:02:24.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="251" reactiontime="+107" swimtime="00:01:27.92" resultid="2514" heatid="2900" lane="3" entrytime="00:01:28.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1430" points="293" reactiontime="+104" swimtime="00:02:50.07" resultid="2515" heatid="2917" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                    <SPLIT distance="100" swimtime="00:01:20.71" />
                    <SPLIT distance="150" swimtime="00:02:05.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Waldemar" lastname="Jagiełło" birthdate="1979-03-01" gender="M" nation="POL" license="502805700042" swrid="4541616" athleteid="2560">
              <RESULTS>
                <RESULT eventid="1140" points="464" reactiontime="+89" swimtime="00:00:33.51" resultid="2561" heatid="2855" lane="6" />
                <RESULT eventid="1172" points="454" reactiontime="+84" swimtime="00:01:01.02" resultid="2562" heatid="2864" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="448" reactiontime="+79" swimtime="00:00:27.32" resultid="2563" heatid="2891" lane="1" />
                <RESULT eventid="1414" points="411" reactiontime="+86" swimtime="00:01:16.50" resultid="2564" heatid="2914" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dagmara" lastname="Luzniakowska" birthdate="1980-04-29" gender="F" nation="POL" athleteid="2090">
              <RESULTS>
                <RESULT eventid="1059" points="110" reactiontime="+101" swimtime="00:00:50.89" resultid="2091" heatid="2837" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1156" points="190" reactiontime="+98" swimtime="00:01:29.81" resultid="2092" heatid="2861" lane="7" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Urszula" lastname="Mróz" birthdate="1962-03-03" gender="F" nation="POL" license="502805600024" swrid="4754660" athleteid="2497">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1059" points="294" reactiontime="+85" swimtime="00:00:36.70" resultid="2498" heatid="2838" lane="0" entrytime="00:00:36.30" entrycourse="LCM" />
                <RESULT eventid="1124" points="249" reactiontime="+104" swimtime="00:00:46.57" resultid="2499" heatid="2851" lane="5" />
                <RESULT eventid="1301" points="315" reactiontime="+93" swimtime="00:00:34.76" resultid="2500" heatid="2888" lane="6" entrytime="00:00:34.31" entrycourse="LCM" />
                <RESULT eventid="1366" points="254" reactiontime="+78" swimtime="00:00:42.55" resultid="2501" heatid="2904" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Chwiałkowski" birthdate="1985-11-09" gender="M" nation="POL" license="502805700033" swrid="5464089" athleteid="2600">
              <RESULTS>
                <RESULT eventid="1382" points="206" reactiontime="+99" swimtime="00:00:40.27" resultid="2601" heatid="2908" lane="2" />
                <RESULT eventid="1446" points="249" reactiontime="+109" swimtime="00:02:42.00" resultid="2602" heatid="2924" lane="3" entrytime="00:02:44.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.52" />
                    <SPLIT distance="100" swimtime="00:01:17.52" />
                    <SPLIT distance="150" swimtime="00:02:00.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrian" lastname="Styrzyński" birthdate="1987-02-16" gender="M" nation="POL" license="502805700147" swrid="4041266" athleteid="2529">
              <RESULTS>
                <RESULT eventid="1076" points="550" reactiontime="+75" swimtime="00:00:27.17" resultid="2530" heatid="2841" lane="5" />
                <RESULT eventid="1140" points="550" reactiontime="+77" swimtime="00:00:31.66" resultid="2531" heatid="2855" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Ścibiorek" birthdate="1971-09-12" gender="F" nation="POL" license="502805600026" swrid="4992745" athleteid="2502">
              <RESULTS>
                <RESULT eventid="1059" points="413" reactiontime="+75" swimtime="00:00:32.78" resultid="2503" heatid="2838" lane="2" entrytime="00:00:32.06" entrycourse="LCM" />
                <RESULT comment="Rekord Polski Masters" eventid="1252" points="398" reactiontime="+85" swimtime="00:02:51.36" resultid="2504" heatid="2878" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                    <SPLIT distance="100" swimtime="00:01:19.83" />
                    <SPLIT distance="150" swimtime="00:02:10.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="421" reactiontime="+83" swimtime="00:01:13.98" resultid="2505" heatid="2900" lane="4" entrytime="00:01:12.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1284" reactiontime="+99" swimtime="00:02:09.37" resultid="2603" heatid="3969" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                    <SPLIT distance="100" swimtime="00:01:09.40" />
                    <SPLIT distance="150" swimtime="00:01:42.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2550" number="1" reactiontime="+99" />
                    <RELAYPOSITION athleteid="2565" number="2" />
                    <RELAYPOSITION athleteid="2827" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="2560" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1494" swimtime="00:02:25.36" resultid="2607" heatid="3989" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.98" />
                    <SPLIT distance="100" swimtime="00:01:19.63" />
                    <SPLIT distance="150" swimtime="00:01:49.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2827" number="1" />
                    <RELAYPOSITION athleteid="2550" number="2" />
                    <RELAYPOSITION athleteid="2560" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="2565" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1284" reactiontime="+94" swimtime="00:02:36.24" resultid="2604" heatid="3970" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.71" />
                    <SPLIT distance="100" swimtime="00:01:19.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2520" number="1" reactiontime="+94" />
                    <RELAYPOSITION athleteid="2532" number="2" />
                    <RELAYPOSITION athleteid="2570" number="3" reactiontime="+90" />
                    <RELAYPOSITION athleteid="2579" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1494" reactiontime="+83" swimtime="00:03:08.19" resultid="2608" heatid="3988" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.98" />
                    <SPLIT distance="100" swimtime="00:01:35.27" />
                    <SPLIT distance="150" swimtime="00:02:23.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2579" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="2532" number="2" />
                    <RELAYPOSITION athleteid="2520" number="3" reactiontime="+2" />
                    <RELAYPOSITION athleteid="2570" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="3">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1284" reactiontime="+85" swimtime="00:01:59.46" resultid="2605" heatid="3969" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                    <SPLIT distance="100" swimtime="00:01:04.24" />
                    <SPLIT distance="150" swimtime="00:01:34.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2502" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="2516" number="2" />
                    <RELAYPOSITION athleteid="2506" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="2529" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1494" reactiontime="+95" swimtime="00:02:13.02" resultid="2609" heatid="3988" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.68" />
                    <SPLIT distance="100" swimtime="00:01:09.40" />
                    <SPLIT distance="150" swimtime="00:01:42.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2516" number="1" reactiontime="+95" />
                    <RELAYPOSITION athleteid="2529" number="2" />
                    <RELAYPOSITION athleteid="2502" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="2506" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="1284" reactiontime="+103" swimtime="00:02:20.16" resultid="2606" heatid="3969" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                    <SPLIT distance="100" swimtime="00:01:10.72" />
                    <SPLIT distance="150" swimtime="00:01:45.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2511" number="1" reactiontime="+103" />
                    <RELAYPOSITION athleteid="2574" number="2" />
                    <RELAYPOSITION athleteid="2555" number="3" reactiontime="+22" />
                    <RELAYPOSITION athleteid="2497" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1494" swimtime="00:02:40.38" resultid="2610" heatid="3987" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.63" />
                    <SPLIT distance="100" swimtime="00:01:25.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2497" number="1" />
                    <RELAYPOSITION athleteid="2555" number="2" />
                    <RELAYPOSITION athleteid="2511" number="3" reactiontime="+69" />
                    <RELAYPOSITION athleteid="2574" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="1747" name="UKS Dwójeczka Częstochowa">
          <ATHLETES>
            <ATHLETE firstname="Ireneusz" lastname="Stachurski" birthdate="1969-07-22" gender="M" nation="POL" license="107311700001" swrid="5464094" athleteid="1748">
              <RESULTS>
                <RESULT eventid="1076" points="118" reactiontime="+101" swimtime="00:00:45.32" resultid="1749" heatid="2842" lane="1" entrytime="00:00:46.00" entrycourse="LCM" />
                <RESULT eventid="1172" points="221" reactiontime="+105" swimtime="00:01:17.53" resultid="1750" heatid="2868" lane="5" entrytime="00:01:02.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="204" reactiontime="+102" swimtime="00:00:35.52" resultid="1751" heatid="2895" lane="9" entrytime="00:00:35.00" entrycourse="LCM" />
                <RESULT eventid="1446" points="197" reactiontime="+101" swimtime="00:02:55.05" resultid="1752" heatid="2921" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                    <SPLIT distance="100" swimtime="00:01:21.07" />
                    <SPLIT distance="150" swimtime="00:02:08.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2062" name="Swim Club Masters Ślęza">
          <ATHLETES>
            <ATHLETE firstname="Joanna" lastname="Chojcan" birthdate="1986-08-04" gender="F" nation="POL" athleteid="2063">
              <RESULTS>
                <RESULT eventid="1092" points="303" reactiontime="+70" swimtime="00:01:25.51" resultid="2064" heatid="2846" lane="1" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="257" reactiontime="+48" swimtime="00:01:27.23" resultid="2065" heatid="2900" lane="5" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="197" reactiontime="+85" swimtime="00:03:29.11" resultid="2066" heatid="2870" lane="4" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                    <SPLIT distance="100" swimtime="00:01:30.63" />
                    <SPLIT distance="150" swimtime="00:02:28.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="289" reactiontime="+77" swimtime="00:03:06.49" resultid="2067" heatid="2927" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.64" />
                    <SPLIT distance="100" swimtime="00:01:30.54" />
                    <SPLIT distance="150" swimtime="00:02:19.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="11514" nation="POL" region="14" clubid="2615" name="Stow. Pływackie Sebastiana Karasia">
          <ATHLETES>
            <ATHLETE firstname="Piotr" lastname="Fuliński" birthdate="1982-06-03" gender="M" nation="POL" license="111514700186" swrid="4992686" athleteid="2616">
              <RESULTS>
                <RESULT eventid="1172" points="502" reactiontime="+80" swimtime="00:00:59.01" resultid="2617" heatid="2864" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="478" reactiontime="+80" swimtime="00:00:26.73" resultid="2618" heatid="2892" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="1899" name="Gdynia Masters">
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Skwarło" birthdate="1939-01-01" gender="M" nation="POL" swrid="4302086" athleteid="1900">
              <RESULTS>
                <RESULT eventid="1140" points="93" reactiontime="+112" swimtime="00:00:57.19" resultid="1901" heatid="2856" lane="2" entrytime="00:00:56.50" />
                <RESULT eventid="1268" points="40" reactiontime="+106" swimtime="00:05:31.45" resultid="1902" heatid="2882" lane="1" entrytime="00:04:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:27.44" />
                    <SPLIT distance="100" swimtime="00:02:57.67" />
                    <SPLIT distance="150" swimtime="00:04:20.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="55" reactiontime="+133" swimtime="00:00:54.73" resultid="1903" heatid="2893" lane="8" entrytime="00:00:53.50" />
                <RESULT eventid="1414" points="66" reactiontime="+155" swimtime="00:02:20.45" resultid="1904" heatid="2914" lane="7" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="12914" nation="POL" region="14" clubid="2708" name="Water Squad">
          <ATHLETES>
            <ATHLETE firstname="Agnieszka" lastname="Kaczmarek" birthdate="1985-05-07" gender="F" nation="POL" license="512914600004" swrid="5240932" athleteid="2709">
              <RESULTS>
                <RESULT eventid="1059" points="415" reactiontime="+85" swimtime="00:00:32.73" resultid="2710" heatid="2836" lane="7" />
                <RESULT eventid="1156" points="418" reactiontime="+82" swimtime="00:01:09.15" resultid="2711" heatid="2859" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="465" reactiontime="+86" swimtime="00:00:30.55" resultid="2712" heatid="2886" lane="1" />
                <RESULT eventid="1366" points="496" reactiontime="+78" swimtime="00:00:34.08" resultid="2713" heatid="2906" lane="2" entrytime="00:00:36.22" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrian" lastname="Kulisz" birthdate="1977-06-16" gender="M" nation="POL" license="512914700002" swrid="5416809" athleteid="2719">
              <RESULTS>
                <RESULT eventid="1076" points="291" reactiontime="+80" swimtime="00:00:33.58" resultid="2720" heatid="2840" lane="8" />
                <RESULT eventid="1172" points="302" reactiontime="+80" swimtime="00:01:09.89" resultid="2721" heatid="2867" lane="6" entrytime="00:01:12.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="263" reactiontime="+108" swimtime="00:00:32.60" resultid="2722" heatid="2896" lane="8" entrytime="00:00:31.48" entrycourse="LCM" />
                <RESULT eventid="1414" points="209" reactiontime="+88" swimtime="00:01:35.72" resultid="2723" heatid="2915" lane="0" entrytime="00:01:35.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Kotlarski" birthdate="1989-05-02" gender="M" nation="POL" license="512914700025" swrid="4071566" athleteid="2750">
              <RESULTS>
                <RESULT eventid="1172" points="451" reactiontime="+75" swimtime="00:01:01.16" resultid="2751" heatid="2865" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="398" reactiontime="+76" swimtime="00:02:34.92" resultid="2752" heatid="2881" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                    <SPLIT distance="100" swimtime="00:01:12.25" />
                    <SPLIT distance="150" swimtime="00:01:57.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Korpetta" birthdate="1959-12-27" gender="M" nation="POL" license="112914700013" swrid="4754654" athleteid="2745">
              <RESULTS>
                <RESULT eventid="1172" points="203" reactiontime="+102" swimtime="00:01:19.74" resultid="2746" heatid="2863" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="133" reactiontime="+112" swimtime="00:03:43.17" resultid="2747" heatid="2882" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.50" />
                    <SPLIT distance="100" swimtime="00:01:51.93" />
                    <SPLIT distance="150" swimtime="00:02:59.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="196" reactiontime="+96" swimtime="00:00:35.96" resultid="2748" heatid="2890" lane="5" />
                <RESULT eventid="1446" points="196" reactiontime="+101" swimtime="00:02:55.53" resultid="2749" heatid="2920" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.71" />
                    <SPLIT distance="100" swimtime="00:01:23.88" />
                    <SPLIT distance="150" swimtime="00:02:10.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Brożyna" birthdate="1980-04-28" gender="M" nation="POL" license="512914700006" swrid="5312396" athleteid="2732">
              <RESULTS>
                <RESULT eventid="1108" points="330" reactiontime="+71" swimtime="00:01:15.03" resultid="2733" heatid="2850" lane="9" entrytime="00:01:16.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="283" reactiontime="+85" swimtime="00:02:53.52" resultid="2734" heatid="2882" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.81" />
                    <SPLIT distance="100" swimtime="00:01:22.76" />
                    <SPLIT distance="150" swimtime="00:02:14.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1382" points="308" reactiontime="+71" swimtime="00:00:35.21" resultid="2735" heatid="2910" lane="8" entrytime="00:00:35.40" entrycourse="LCM" />
                <RESULT eventid="1478" points="307" reactiontime="+73" swimtime="00:02:45.87" resultid="2736" heatid="2930" lane="6" entrytime="00:02:41.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.94" />
                    <SPLIT distance="150" swimtime="00:02:04.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Kaczmarek" birthdate="1977-06-25" gender="M" nation="POL" license="512914700003" swrid="4043251" athleteid="2724">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1076" points="612" reactiontime="+80" swimtime="00:00:26.22" resultid="2725" heatid="2841" lane="3" />
                <RESULT eventid="1172" points="569" reactiontime="+83" swimtime="00:00:56.59" resultid="2726" heatid="2869" lane="4" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.28" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1382" points="611" reactiontime="+70" swimtime="00:00:28.04" resultid="2727" heatid="2907" lane="4" />
                <RESULT eventid="1446" status="DNS" swimtime="00:00:00.00" resultid="2728" heatid="2925" lane="5" entrytime="00:02:02.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Szyszkowska" birthdate="1996-11-05" gender="F" nation="POL" license="512914600054" swrid="4282341" athleteid="2714">
              <RESULTS>
                <RESULT eventid="1059" points="449" reactiontime="+88" swimtime="00:00:31.90" resultid="2715" heatid="2838" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="1124" points="539" reactiontime="+93" swimtime="00:00:36.00" resultid="2716" heatid="2853" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="1301" points="528" reactiontime="+83" swimtime="00:00:29.28" resultid="2717" heatid="2889" lane="2" entrytime="00:00:28.50" />
                <RESULT eventid="1398" points="485" reactiontime="+88" swimtime="00:01:21.58" resultid="2718" heatid="2912" lane="4" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hubert" lastname="Markowski" birthdate="1976-01-04" gender="M" nation="POL" license="512914700011" swrid="5471789" athleteid="2729">
              <RESULTS>
                <RESULT eventid="1076" points="386" reactiontime="+80" swimtime="00:00:30.56" resultid="2730" heatid="2843" lane="1" entrytime="00:00:31.47" entrycourse="LCM" />
                <RESULT eventid="1204" points="282" reactiontime="+92" swimtime="00:02:48.82" resultid="2731" heatid="2872" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                    <SPLIT distance="100" swimtime="00:01:18.36" />
                    <SPLIT distance="150" swimtime="00:02:02.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Romuald" lastname="Kozłowski" birthdate="1966-08-13" gender="M" nation="POL" license="512914700012" swrid="5425564" athleteid="2741">
              <RESULTS>
                <RESULT eventid="1140" points="396" reactiontime="+78" swimtime="00:00:35.33" resultid="2742" heatid="2858" lane="1" entrytime="00:00:34.92" entrycourse="LCM" />
                <RESULT eventid="1318" points="384" reactiontime="+73" swimtime="00:00:28.75" resultid="2743" heatid="2892" lane="1" />
                <RESULT eventid="1414" points="333" reactiontime="+82" swimtime="00:01:22.05" resultid="2744" heatid="2916" lane="1" entrytime="00:01:17.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Kośmider" birthdate="1966-03-01" gender="M" nation="POL" license="512914700009" swrid="4992964" athleteid="2753">
              <RESULTS>
                <RESULT eventid="1236" points="292" reactiontime="+85" swimtime="00:03:10.00" resultid="2754" heatid="2877" lane="7" entrytime="00:03:17.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.18" />
                    <SPLIT distance="100" swimtime="00:01:29.33" />
                    <SPLIT distance="150" swimtime="00:02:18.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="315" reactiontime="+79" swimtime="00:02:29.78" resultid="2755" heatid="2924" lane="4" entrytime="00:02:31.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                    <SPLIT distance="100" swimtime="00:01:13.57" />
                    <SPLIT distance="150" swimtime="00:01:51.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1284" reactiontime="+84" swimtime="00:01:52.52" resultid="2756" heatid="3969" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.82" />
                    <SPLIT distance="100" swimtime="00:00:55.37" />
                    <SPLIT distance="150" swimtime="00:01:23.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2724" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="2709" number="2" />
                    <RELAYPOSITION athleteid="2714" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="2741" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1494" reactiontime="+74" swimtime="00:02:04.98" resultid="2757" heatid="3989" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.13" />
                    <SPLIT distance="100" swimtime="00:01:03.93" />
                    <SPLIT distance="150" swimtime="00:01:36.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2724" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="2741" number="2" />
                    <RELAYPOSITION athleteid="2709" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="2714" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="UKR" clubid="2762" name="Ukraine Swim Team">
          <ATHLETES>
            <ATHLETE firstname="Valeriia" lastname="Khokhol" birthdate="1996-08-21" gender="F" nation="UKR" athleteid="2778">
              <RESULTS>
                <RESULT eventid="1301" points="368" reactiontime="+97" swimtime="00:00:33.03" resultid="2779" heatid="2889" lane="9" entrytime="00:00:32.01" />
                <RESULT eventid="1124" points="309" reactiontime="+106" swimtime="00:00:43.33" resultid="2780" heatid="2853" lane="6" entrytime="00:00:39.02" />
                <RESULT eventid="1398" points="310" reactiontime="+96" swimtime="00:01:34.75" resultid="2781" heatid="2912" lane="2" entrytime="00:01:28.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yevgeniya" lastname="Motrych" birthdate="1983-11-07" gender="F" nation="UKR" athleteid="2773">
              <RESULTS>
                <RESULT eventid="1124" points="228" reactiontime="+115" swimtime="00:00:47.91" resultid="2774" heatid="2853" lane="9" entrytime="00:00:47.19" />
                <RESULT eventid="1156" points="156" reactiontime="+104" swimtime="00:01:35.89" resultid="2775" heatid="2861" lane="0" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1398" points="224" reactiontime="+99" swimtime="00:01:45.46" resultid="2776" heatid="2911" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1430" points="162" reactiontime="+101" swimtime="00:03:26.87" resultid="2777" heatid="2918" lane="6" entrytime="00:03:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.24" />
                    <SPLIT distance="100" swimtime="00:01:36.79" />
                    <SPLIT distance="150" swimtime="00:02:32.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nataliia" lastname="Boryshkevych" birthdate="1976-04-15" gender="F" nation="UKR" swrid="5241793" athleteid="2763">
              <RESULTS>
                <RESULT eventid="1059" points="212" reactiontime="+86" swimtime="00:00:40.96" resultid="2764" heatid="2837" lane="4" entrytime="00:00:37.00" />
                <RESULT eventid="1156" points="362" reactiontime="+88" swimtime="00:01:12.49" resultid="2765" heatid="2862" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="196" reactiontime="+90" swimtime="00:01:35.45" resultid="2766" heatid="2900" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1430" points="329" reactiontime="+89" swimtime="00:02:43.58" resultid="2767" heatid="2919" lane="7" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                    <SPLIT distance="100" swimtime="00:01:19.13" />
                    <SPLIT distance="150" swimtime="00:02:02.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Iryna" lastname="Oriekhova" birthdate="1988-05-19" gender="F" nation="UKR" athleteid="2768">
              <RESULTS>
                <RESULT eventid="1156" points="235" reactiontime="+104" swimtime="00:01:23.71" resultid="2769" heatid="2860" lane="4" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="238" reactiontime="+104" swimtime="00:03:23.34" resultid="2770" heatid="2879" lane="6" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.03" />
                    <SPLIT distance="100" swimtime="00:01:36.90" />
                    <SPLIT distance="150" swimtime="00:02:33.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="257" reactiontime="+107" swimtime="00:00:42.43" resultid="2771" heatid="2905" lane="4" entrytime="00:00:50.00" />
                <RESULT eventid="1430" points="223" reactiontime="+98" swimtime="00:03:06.28" resultid="2772" heatid="2918" lane="3" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.47" />
                    <SPLIT distance="100" swimtime="00:01:29.22" />
                    <SPLIT distance="150" swimtime="00:02:18.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="14" clubid="3975" name="LEGIA Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Bogdan" lastname="Dubiński" birthdate="1953-05-05" gender="M" nation="POL" swrid="4992696" athleteid="1923">
              <RESULTS>
                <RESULT eventid="1172" points="186" reactiontime="+96" swimtime="00:01:22.08" resultid="1924" heatid="2863" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="118" reactiontime="+102" swimtime="00:03:51.88" resultid="1925" heatid="2880" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.45" />
                    <SPLIT distance="100" swimtime="00:01:55.72" />
                    <SPLIT distance="150" swimtime="00:03:04.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="192" reactiontime="+90" swimtime="00:00:36.24" resultid="1926" heatid="2894" lane="3" entrytime="00:00:36.00" />
                <RESULT eventid="1382" points="159" reactiontime="+75" swimtime="00:00:43.91" resultid="1927" heatid="2909" lane="2" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="1916" name="UKS TRÓJKA Puławy">
          <ATHLETES>
            <ATHLETE firstname="Sebastian" lastname="Gogacz" birthdate="1976-10-28" gender="M" nation="POL" license="501203700057" swrid="4754646" athleteid="1917">
              <RESULTS>
                <RESULT eventid="1204" points="360" reactiontime="+83" swimtime="00:02:35.54" resultid="1918" heatid="2872" lane="4" entrytime="00:02:39.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                    <SPLIT distance="100" swimtime="00:01:15.32" />
                    <SPLIT distance="150" swimtime="00:01:55.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="324" reactiontime="+87" swimtime="00:02:45.82" resultid="1919" heatid="2883" lane="6" entrytime="00:02:44.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                    <SPLIT distance="100" swimtime="00:01:23.16" />
                    <SPLIT distance="150" swimtime="00:02:08.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="tomasz" lastname="bielawski" birthdate="1976-09-22" gender="M" nation="POL" license="501203700070" athleteid="1920">
              <RESULTS>
                <RESULT eventid="1108" points="255" reactiontime="+102" swimtime="00:01:21.74" resultid="1921" heatid="2850" lane="0" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="358" reactiontime="+102" swimtime="00:01:06.03" resultid="1922" heatid="2868" lane="2" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00309" nation="POL" region="09" clubid="2493" name="MKS Juvenia Białystok">
          <ATHLETES>
            <ATHLETE firstname="Dominika" lastname="Michalik" birthdate="1979-07-14" gender="F" nation="POL" license="500309600228" swrid="4595750" athleteid="2494">
              <RESULTS>
                <RESULT eventid="1156" points="462" reactiontime="+78" swimtime="00:01:06.88" resultid="2495" heatid="2862" lane="2" entrytime="00:01:07.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1430" points="442" reactiontime="+82" swimtime="00:02:28.27" resultid="2496" heatid="2919" lane="6" entrytime="00:02:26.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                    <SPLIT distance="100" swimtime="00:01:10.05" />
                    <SPLIT distance="150" swimtime="00:01:48.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02906" nation="POL" region="06" clubid="2611" name="SSKSiT GLOSATOR Kraków">
          <ATHLETES>
            <ATHLETE firstname="Elżbieta" lastname="Hamowska" birthdate="1960-03-20" gender="F" nation="POL" license="502906600058" swrid="5297381" athleteid="2612">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="2613" heatid="2845" lane="0" />
                <RESULT eventid="1156" status="DNS" swimtime="00:00:00.00" resultid="2614" heatid="2859" lane="7" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="01" clubid="1555" name="Masters Wrocław">
          <ATHLETES>
            <ATHLETE firstname="Piotr" lastname="Krzekotowski" birthdate="1966-01-01" gender="M" nation="POL" swrid="5416779" athleteid="1561">
              <RESULTS>
                <RESULT eventid="1108" points="88" reactiontime="+93" swimtime="00:01:56.49" resultid="1562" heatid="2848" lane="5" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="120" reactiontime="+95" swimtime="00:03:50.62" resultid="1563" heatid="2882" lane="4" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.63" />
                    <SPLIT distance="100" swimtime="00:01:57.78" />
                    <SPLIT distance="150" swimtime="00:03:01.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="69" reactiontime="+88" swimtime="00:02:00.54" resultid="1564" heatid="2902" lane="2" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="115" reactiontime="+97" swimtime="00:03:29.54" resultid="1565" heatid="2923" lane="8" entrytime="00:03:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.90" />
                    <SPLIT distance="150" swimtime="00:02:35.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Marszałek" birthdate="1954-01-01" gender="M" nation="POL" athleteid="1556">
              <RESULTS>
                <RESULT eventid="1076" points="73" swimtime="00:00:53.17" resultid="1557" heatid="2842" lane="0" entrytime="00:00:51.00" />
                <RESULT eventid="1268" points="90" reactiontime="+104" swimtime="00:04:14.13" resultid="1558" heatid="2882" lane="6" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.32" />
                    <SPLIT distance="100" swimtime="00:02:07.88" />
                    <SPLIT distance="150" swimtime="00:03:18.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="127" swimtime="00:00:41.55" resultid="1559" heatid="2893" lane="5" entrytime="00:00:43.00" />
                <RESULT eventid="1446" points="98" reactiontime="+96" swimtime="00:03:40.99" resultid="1560" heatid="2922" lane="4" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.50" />
                    <SPLIT distance="100" swimtime="00:01:49.34" />
                    <SPLIT distance="150" swimtime="00:02:46.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00211" nation="POL" clubid="1803" name="KS. Górnik Radlin">
          <ATHLETES>
            <ATHLETE firstname="Ryszard" lastname="Kubica" birthdate="1972-02-22" gender="M" nation="POL" license="100211700343" swrid="5398297" athleteid="1804">
              <RESULTS>
                <RESULT eventid="1108" points="251" reactiontime="+78" swimtime="00:01:22.10" resultid="1805" heatid="2849" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="212" reactiontime="+102" swimtime="00:03:05.70" resultid="1806" heatid="2872" lane="3" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.67" />
                    <SPLIT distance="100" swimtime="00:01:23.67" />
                    <SPLIT distance="150" swimtime="00:02:13.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="281" reactiontime="+98" swimtime="00:01:15.45" resultid="1807" heatid="2903" lane="0" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1478" points="235" reactiontime="+82" swimtime="00:03:01.27" resultid="1808" heatid="2930" lane="9" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.60" />
                    <SPLIT distance="100" swimtime="00:01:27.42" />
                    <SPLIT distance="150" swimtime="00:02:16.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="1753" name="IKS DSS Kraków">
          <ATHLETES>
            <ATHLETE firstname="Ewa" lastname="Rupp" birthdate="1956-03-06" gender="F" nation="POL" license="505806600021" swrid="5484417" athleteid="1754">
              <RESULTS>
                <RESULT eventid="1092" points="68" reactiontime="+81" swimtime="00:02:20.50" resultid="1755" heatid="2845" lane="4" entrytime="00:02:11.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="88" reactiontime="+121" swimtime="00:01:55.89" resultid="1756" heatid="2860" lane="1" entrytime="00:01:58.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="30" reactiontime="+122" swimtime="00:02:56.95" resultid="1757" heatid="2900" lane="1" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="85" reactiontime="+84" swimtime="00:04:40.46" resultid="1758" heatid="2927" lane="0" entrytime="00:04:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.39" />
                    <SPLIT distance="100" swimtime="00:02:19.04" />
                    <SPLIT distance="150" swimtime="00:03:32.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="1981" name="Klub Sportowy Mako">
          <ATHLETES>
            <ATHLETE firstname="Marek" lastname="Piórkowski" birthdate="1965-07-28" gender="M" nation="POL" license="510414700072" swrid="5506637" athleteid="2188">
              <RESULTS>
                <RESULT eventid="1108" points="109" reactiontime="+79" swimtime="00:01:48.51" resultid="2214" heatid="2847" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="132" reactiontime="+100" swimtime="00:01:31.90" resultid="2215" heatid="2864" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1382" points="116" reactiontime="+74" swimtime="00:00:48.76" resultid="2216" heatid="2907" lane="1" />
                <RESULT eventid="1478" points="93" reactiontime="+79" swimtime="00:04:06.87" resultid="2217" heatid="2928" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.19" />
                    <SPLIT distance="100" swimtime="00:02:00.37" />
                    <SPLIT distance="150" swimtime="00:03:06.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Matusiewicz" birthdate="1998-04-12" gender="M" nation="POL" swrid="5058424" athleteid="1982">
              <RESULTS>
                <RESULT eventid="1108" points="124" reactiontime="+116" swimtime="00:01:43.90" resultid="1983" heatid="2849" lane="0" entrytime="00:01:50.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="118" reactiontime="+114" swimtime="00:03:51.91" resultid="1984" heatid="2883" lane="0" entrytime="00:03:46.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.61" />
                    <SPLIT distance="100" swimtime="00:01:49.94" />
                    <SPLIT distance="150" swimtime="00:02:55.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="116" reactiontime="+86" swimtime="00:00:42.79" resultid="1985" heatid="2894" lane="9" entrytime="00:00:41.23" />
                <RESULT eventid="1414" points="103" reactiontime="+86" swimtime="00:02:01.00" resultid="1986" heatid="2914" lane="6" entrytime="00:01:55.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Adamowicz" birthdate="1967-07-11" gender="M" nation="POL" license="510414700009" swrid="4655152" athleteid="2198">
              <RESULTS>
                <RESULT eventid="1318" points="156" reactiontime="+71" swimtime="00:00:38.78" resultid="2201" heatid="2890" lane="4" />
                <RESULT eventid="1140" points="200" reactiontime="+77" swimtime="00:00:44.35" resultid="2222" heatid="2857" lane="8" entrytime="00:00:45.48" entrycourse="LCM" />
                <RESULT eventid="1236" points="145" reactiontime="+80" swimtime="00:03:59.84" resultid="2223" heatid="2875" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.62" />
                    <SPLIT distance="100" swimtime="00:01:55.73" />
                    <SPLIT distance="150" swimtime="00:03:01.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="89" reactiontime="+89" swimtime="00:03:47.79" resultid="2225" heatid="2920" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.39" />
                    <SPLIT distance="100" swimtime="00:01:45.97" />
                    <SPLIT distance="150" swimtime="00:02:47.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Timea" lastname="Balajcza" birthdate="1971-09-22" gender="F" nation="POL" license="510414600003" swrid="5240601" athleteid="2193">
              <RESULTS>
                <RESULT eventid="1124" points="435" reactiontime="+92" swimtime="00:00:38.66" resultid="2194" heatid="2853" lane="2" entrytime="00:00:39.14" entrycourse="LCM" />
                <RESULT comment="Rekord Polski Masters" eventid="1220" points="386" reactiontime="+84" swimtime="00:03:10.80" resultid="2219" heatid="2874" lane="4" entrytime="00:03:18.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.75" />
                    <SPLIT distance="100" swimtime="00:01:32.21" />
                    <SPLIT distance="150" swimtime="00:02:22.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1398" points="397" reactiontime="+78" swimtime="00:01:27.19" resultid="2220" heatid="2912" lane="1" entrytime="00:01:31.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1430" points="293" reactiontime="+87" swimtime="00:02:50.08" resultid="2221" heatid="2918" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.25" />
                    <SPLIT distance="100" swimtime="00:01:22.29" />
                    <SPLIT distance="150" swimtime="00:02:07.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Rudziński" birthdate="1966-05-10" gender="M" nation="POL" license="510414700010" swrid="4934041" athleteid="2203">
              <RESULTS>
                <RESULT eventid="1382" points="87" reactiontime="+108" swimtime="00:00:53.61" resultid="2207" heatid="2907" lane="3" />
                <RESULT eventid="1204" points="101" reactiontime="+104" swimtime="00:03:57.21" resultid="2226" heatid="2872" lane="1" entrytime="00:04:08.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.25" />
                    <SPLIT distance="100" swimtime="00:01:47.71" />
                    <SPLIT distance="150" swimtime="00:02:51.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="199" reactiontime="+111" swimtime="00:03:35.82" resultid="2227" heatid="2875" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.96" />
                    <SPLIT distance="100" swimtime="00:01:42.06" />
                    <SPLIT distance="150" swimtime="00:02:39.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1318" points="141" reactiontime="+112" swimtime="00:00:40.11" resultid="2228" heatid="2891" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Dąbrowska" birthdate="1987-05-20" gender="F" nation="POL" license="510414600006" swrid="4655165" athleteid="2183">
              <RESULTS>
                <RESULT eventid="1156" points="172" reactiontime="+104" swimtime="00:01:32.92" resultid="2185" heatid="2859" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1430" points="143" reactiontime="+116" swimtime="00:03:36.03" resultid="2187" heatid="2917" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.16" />
                    <SPLIT distance="100" swimtime="00:01:43.52" />
                    <SPLIT distance="150" swimtime="00:02:40.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="104" reactiontime="+101" swimtime="00:02:02.12" resultid="2210" heatid="2845" lane="2" />
                <RESULT eventid="1366" points="123" swimtime="00:00:54.15" resultid="2212" heatid="2904" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sebastian" lastname="Ostapczuk" birthdate="1970-07-13" gender="M" nation="POL" athleteid="1987">
              <RESULTS>
                <RESULT eventid="1172" status="DNS" swimtime="00:00:00.00" resultid="1988" heatid="2866" lane="7" entrytime="00:01:29.00" />
                <RESULT eventid="1236" status="DNS" swimtime="00:00:00.00" resultid="1989" heatid="2876" lane="4" entrytime="00:03:35.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1494" reactiontime="+88" swimtime="00:02:51.08" resultid="2209" heatid="3989" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.05" />
                    <SPLIT distance="100" swimtime="00:01:27.36" />
                    <SPLIT distance="150" swimtime="00:02:09.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2188" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="2193" number="2" />
                    <RELAYPOSITION athleteid="2203" number="3" reactiontime="+78" />
                    <RELAYPOSITION athleteid="2183" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1284" reactiontime="+108" swimtime="00:02:34.44" resultid="2230" heatid="3969" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.32" />
                    <SPLIT distance="100" swimtime="00:01:22.74" />
                    <SPLIT distance="150" swimtime="00:02:00.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2183" number="1" reactiontime="+108" />
                    <RELAYPOSITION athleteid="2188" number="2" />
                    <RELAYPOSITION athleteid="2198" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="2193" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="1741" name="Motyl MOSiR Stalowa Wola">
          <ATHLETES>
            <ATHLETE firstname="Arkadiusz" lastname="Berwecki" birthdate="1973-01-14" gender="M" nation="POL" swrid="4791744" athleteid="1742">
              <RESULTS>
                <RESULT eventid="1076" points="462" reactiontime="+82" swimtime="00:00:28.79" resultid="1743" heatid="2844" lane="7" entrytime="00:00:27.89" />
                <RESULT eventid="1268" points="423" reactiontime="+80" swimtime="00:02:31.85" resultid="1744" heatid="2883" lane="4" entrytime="00:02:24.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                    <SPLIT distance="100" swimtime="00:01:12.31" />
                    <SPLIT distance="150" swimtime="00:01:54.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="461" reactiontime="+78" swimtime="00:01:03.99" resultid="1745" heatid="2903" lane="3" entrytime="00:01:02.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="438" reactiontime="+82" swimtime="00:02:14.23" resultid="1746" heatid="2925" lane="6" entrytime="00:02:07.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                    <SPLIT distance="100" swimtime="00:01:04.39" />
                    <SPLIT distance="150" swimtime="00:01:39.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02706" nation="POL" region="06" clubid="2631" name="UKS Jasień Sucha Beskidzka">
          <ATHLETES>
            <ATHLETE firstname="Sabina" lastname="Sikora" birthdate="1984-10-03" gender="F" nation="POL" license="102706600159" swrid="5468086" athleteid="2632">
              <RESULTS>
                <RESULT eventid="1124" points="460" reactiontime="+89" swimtime="00:00:37.94" resultid="2633" heatid="2853" lane="1" entrytime="00:00:42.21" entrycourse="LCM" />
                <RESULT eventid="1220" points="334" reactiontime="+90" swimtime="00:03:20.19" resultid="2634" heatid="2874" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.16" />
                    <SPLIT distance="100" swimtime="00:01:38.07" />
                    <SPLIT distance="150" swimtime="00:02:29.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1301" points="469" reactiontime="+82" swimtime="00:00:30.46" resultid="2635" heatid="2888" lane="4" entrytime="00:00:32.31" entrycourse="LCM" />
                <RESULT eventid="1398" points="359" reactiontime="+84" swimtime="00:01:30.23" resultid="2636" heatid="2912" lane="8" entrytime="00:01:34.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03315" nation="POL" region="15" clubid="2417" name="KU AZS UAM Poznań">
          <ATHLETES>
            <ATHLETE firstname="Jacek" lastname="Thiem" birthdate="1963-02-17" gender="M" nation="POL" license="503315700211" swrid="4754725" athleteid="2418">
              <RESULTS>
                <RESULT eventid="1076" points="173" reactiontime="+98" swimtime="00:00:39.90" resultid="2419" heatid="2840" lane="4" />
                <RESULT eventid="1204" points="139" reactiontime="+113" swimtime="00:03:33.30" resultid="2420" heatid="2871" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.74" />
                    <SPLIT distance="100" swimtime="00:01:46.39" />
                    <SPLIT distance="150" swimtime="00:02:42.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="162" reactiontime="+107" swimtime="00:01:30.68" resultid="2421" heatid="2902" lane="5" entrytime="00:01:30.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="157" reactiontime="+113" swimtime="00:03:08.91" resultid="2422" heatid="2923" lane="4" entrytime="00:03:08.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.28" />
                    <SPLIT distance="100" swimtime="00:01:35.09" />
                    <SPLIT distance="150" swimtime="00:02:24.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>

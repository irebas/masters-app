<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="SiKReT Gliwice" version="11.51721">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" phone="+41 99 999 99 99" fax="+41 99 999 99 99" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Gliwice" name="Zimowe Mistrzostwa Polski w Pływaniu Masters" course="SCM" hostclub="SiKReT Gliwice" hostclub.url="http://www.sikret-plywanie.pl" organizer="Samorząd Miasta Gliwice, MZUK Gliwice, PZP,SLOZP,SiKReT Gliwice" reservecount="2" result.url="http://www.megatiming.pl" startmethod="1" timing="AUTOMATIC" nation="POL">
      <AGEDATE value="2017-11-17" type="YEAR" />
      <POOL name="Olimpijczyk Gliwice" lanemax="9" />
      <FACILITY city="Gliwice" name="Olimpijczyk Gliwice" nation="POL" />
      <POINTTABLE pointtableid="3010" name="FINA Point Scoring" version="2017" />
      <CONTACT email="wisniowicz@interia.pl" name="Wojciech Wiśniowicz" phone="500193225" />
      <FEES>
        <FEE currency="PLN" type="ATHLETE" value="11000" />
        <FEE currency="PLN" type="LATEENTRY.INDIVIDUAL" value="15000" />
      </FEES>
      <SESSIONS>
        <SESSION date="2017-11-17" daytime="14:45" endtime="21:41" name="BLOK I" number="1" warmupfrom="13:30">
          <EVENTS>
            <EVENT eventid="14189" daytime="18:05" gender="M" number="7" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="19641" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="16620" />
                    <RANKING order="2" place="-1" resultid="17989" />
                    <RANKING order="3" place="-1" resultid="18613" />
                    <RANKING order="4" place="-1" resultid="18337" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19642" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18499" />
                    <RANKING order="2" place="-1" resultid="15388" />
                    <RANKING order="3" place="-1" resultid="17975" />
                    <RANKING order="4" place="-1" resultid="16631" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19643" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14430" />
                    <RANKING order="2" place="2" resultid="16545" />
                    <RANKING order="3" place="3" resultid="15757" />
                    <RANKING order="4" place="4" resultid="14945" />
                    <RANKING order="5" place="5" resultid="14447" />
                    <RANKING order="6" place="-1" resultid="15897" />
                    <RANKING order="7" place="-1" resultid="18952" />
                    <RANKING order="8" place="-1" resultid="18153" />
                    <RANKING order="9" place="-1" resultid="17935" />
                    <RANKING order="10" place="-1" resultid="17984" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19644" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17170" />
                    <RANKING order="2" place="2" resultid="18205" />
                    <RANKING order="3" place="-1" resultid="18969" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19645" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18182" />
                    <RANKING order="2" place="2" resultid="16837" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19646" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14861" />
                    <RANKING order="2" place="2" resultid="18221" />
                    <RANKING order="3" place="3" resultid="14706" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19647" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17221" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19648" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18213" />
                    <RANKING order="2" place="2" resultid="17309" />
                    <RANKING order="3" place="3" resultid="16228" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19649" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17747" />
                    <RANKING order="2" place="2" resultid="14438" />
                    <RANKING order="3" place="-1" resultid="18437" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19650" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17108" />
                    <RANKING order="2" place="2" resultid="17733" />
                    <RANKING order="3" place="3" resultid="15215" />
                    <RANKING order="4" place="4" resultid="15825" />
                    <RANKING order="5" place="5" resultid="14656" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19651" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18330" />
                    <RANKING order="2" place="-1" resultid="17284" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19652" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="14927" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19653" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="19654" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="19655" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="19656" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19614" daytime="18:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19615" daytime="18:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19616" daytime="18:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19617" daytime="18:55" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1130" daytime="16:45" gender="X" number="5" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="12486" agemax="99" agemin="80" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16644" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1182" agemax="119" agemin="100" calculate="TOTAL" />
                <AGEGROUP agegroupid="1183" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17512" />
                    <RANKING order="2" place="2" resultid="16886" />
                    <RANKING order="3" place="3" resultid="18399" />
                    <RANKING order="4" place="4" resultid="18010" />
                    <RANKING order="5" place="5" resultid="18012" />
                    <RANKING order="6" place="6" resultid="17117" />
                    <RANKING order="7" place="7" resultid="18226" />
                    <RANKING order="8" place="8" resultid="17869" />
                    <RANKING order="9" place="9" resultid="15912" />
                    <RANKING order="10" place="10" resultid="16642" />
                    <RANKING order="11" place="11" resultid="16304" />
                    <RANKING order="12" place="-1" resultid="17717" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1184" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17653" />
                    <RANKING order="2" place="2" resultid="15302" />
                    <RANKING order="3" place="3" resultid="16087" />
                    <RANKING order="4" place="4" resultid="17866" />
                    <RANKING order="5" place="5" resultid="17513" />
                    <RANKING order="6" place="6" resultid="17240" />
                    <RANKING order="7" place="7" resultid="18225" />
                    <RANKING order="8" place="8" resultid="15965" />
                    <RANKING order="9" place="-1" resultid="15366" />
                    <RANKING order="10" place="-1" resultid="17867" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1185" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16479" />
                    <RANKING order="2" place="2" resultid="14718" />
                    <RANKING order="3" place="3" resultid="16206" />
                    <RANKING order="4" place="-1" resultid="17239" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1186" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15303" />
                    <RANKING order="2" place="2" resultid="14533" />
                    <RANKING order="3" place="3" resultid="16480" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1145" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14532" />
                    <RANKING order="2" place="2" resultid="16481" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19319" daytime="16:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19320" daytime="16:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19321" daytime="16:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19322" daytime="16:55" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1147" daytime="17:10" gender="F" number="6" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="19625" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14984" />
                    <RANKING order="2" place="-1" resultid="16964" />
                    <RANKING order="3" place="-1" resultid="18200" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19626" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="14646" />
                    <RANKING order="2" place="-1" resultid="18095" />
                    <RANKING order="3" place="-1" resultid="18411" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19627" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17709" />
                    <RANKING order="2" place="2" resultid="18361" />
                    <RANKING order="3" place="-1" resultid="18424" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19628" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15852" />
                    <RANKING order="2" place="2" resultid="17928" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19629" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16007" />
                    <RANKING order="2" place="-1" resultid="14890" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19630" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14526" />
                    <RANKING order="2" place="2" resultid="17329" />
                    <RANKING order="3" place="3" resultid="17099" />
                    <RANKING order="4" place="-1" resultid="15338" />
                    <RANKING order="5" place="-1" resultid="14808" />
                    <RANKING order="6" place="-1" resultid="14799" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19631" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15795" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19632" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16466" />
                    <RANKING order="2" place="-1" resultid="16349" />
                    <RANKING order="3" place="-1" resultid="14508" />
                    <RANKING order="4" place="-1" resultid="16157" />
                    <RANKING order="5" place="-1" resultid="14487" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19633" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16388" />
                    <RANKING order="2" place="-1" resultid="19742" />
                    <RANKING order="3" place="-1" resultid="17189" />
                    <RANKING order="4" place="-1" resultid="14844" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19634" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17435" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19635" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="14403" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19636" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="19637" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="19638" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18310" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19639" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="19640" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19594" daytime="17:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19595" daytime="17:35" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="19606" daytime="19:40" gender="M" number="9" order="12" round="FHT" preveventid="14207">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="19623" daytime="19:40" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1113" daytime="16:10" gender="M" number="4" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1114" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17323" />
                    <RANKING order="2" place="2" resultid="16213" />
                    <RANKING order="3" place="3" resultid="18052" />
                    <RANKING order="4" place="4" resultid="16266" />
                    <RANKING order="5" place="-1" resultid="15015" />
                    <RANKING order="6" place="-1" resultid="18567" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1115" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16741" />
                    <RANKING order="2" place="2" resultid="18165" />
                    <RANKING order="3" place="3" resultid="18498" />
                    <RANKING order="4" place="4" resultid="15749" />
                    <RANKING order="5" place="5" resultid="17293" />
                    <RANKING order="6" place="6" resultid="15889" />
                    <RANKING order="7" place="7" resultid="15387" />
                    <RANKING order="8" place="8" resultid="18347" />
                    <RANKING order="9" place="9" resultid="16276" />
                    <RANKING order="10" place="-1" resultid="15436" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1116" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15756" />
                    <RANKING order="2" place="2" resultid="15896" />
                    <RANKING order="3" place="3" resultid="16879" />
                    <RANKING order="4" place="4" resultid="17303" />
                    <RANKING order="5" place="5" resultid="15443" />
                    <RANKING order="6" place="6" resultid="18387" />
                    <RANKING order="7" place="7" resultid="18124" />
                    <RANKING order="8" place="-1" resultid="17353" />
                    <RANKING order="9" place="-1" resultid="16614" />
                    <RANKING order="10" place="-1" resultid="18585" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1117" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17169" />
                    <RANKING order="2" place="2" resultid="17019" />
                    <RANKING order="3" place="3" resultid="15293" />
                    <RANKING order="4" place="4" resultid="17370" />
                    <RANKING order="5" place="5" resultid="16824" />
                    <RANKING order="6" place="6" resultid="17272" />
                    <RANKING order="7" place="7" resultid="17577" />
                    <RANKING order="8" place="8" resultid="16857" />
                    <RANKING order="9" place="-1" resultid="15905" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1118" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16970" />
                    <RANKING order="2" place="2" resultid="15056" />
                    <RANKING order="3" place="3" resultid="18554" />
                    <RANKING order="4" place="4" resultid="16023" />
                    <RANKING order="5" place="5" resultid="18046" />
                    <RANKING order="6" place="6" resultid="18417" />
                    <RANKING order="7" place="7" resultid="18527" />
                    <RANKING order="8" place="8" resultid="16041" />
                    <RANKING order="9" place="9" resultid="17792" />
                    <RANKING order="10" place="10" resultid="17757" />
                    <RANKING order="11" place="11" resultid="14421" />
                    <RANKING order="12" place="12" resultid="16587" />
                    <RANKING order="13" place="-1" resultid="14635" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1119" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18561" />
                    <RANKING order="2" place="2" resultid="14965" />
                    <RANKING order="3" place="3" resultid="16067" />
                    <RANKING order="4" place="4" resultid="16032" />
                    <RANKING order="5" place="5" resultid="17670" />
                    <RANKING order="6" place="6" resultid="15988" />
                    <RANKING order="7" place="7" resultid="16074" />
                    <RANKING order="8" place="8" resultid="17649" />
                    <RANKING order="9" place="-1" resultid="18447" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1120" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17338" />
                    <RANKING order="2" place="2" resultid="18456" />
                    <RANKING order="3" place="3" resultid="14908" />
                    <RANKING order="4" place="4" resultid="18535" />
                    <RANKING order="5" place="5" resultid="15924" />
                    <RANKING order="6" place="6" resultid="17679" />
                    <RANKING order="7" place="7" resultid="16125" />
                    <RANKING order="8" place="8" resultid="15857" />
                    <RANKING order="9" place="9" resultid="16430" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1121" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15741" />
                    <RANKING order="2" place="2" resultid="17178" />
                    <RANKING order="3" place="3" resultid="14348" />
                    <RANKING order="4" place="4" resultid="16322" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1122" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17410" />
                    <RANKING order="2" place="2" resultid="15397" />
                    <RANKING order="3" place="3" resultid="17746" />
                    <RANKING order="4" place="4" resultid="15936" />
                    <RANKING order="5" place="5" resultid="16245" />
                    <RANKING order="6" place="6" resultid="15255" />
                    <RANKING order="7" place="-1" resultid="14394" />
                    <RANKING order="8" place="-1" resultid="14727" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1123" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17449" />
                    <RANKING order="2" place="2" resultid="18266" />
                    <RANKING order="3" place="3" resultid="14655" />
                    <RANKING order="4" place="4" resultid="17053" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1124" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14358" />
                    <RANKING order="2" place="2" resultid="17739" />
                    <RANKING order="3" place="3" resultid="16330" />
                    <RANKING order="4" place="4" resultid="14412" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1125" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14453" />
                    <RANKING order="2" place="2" resultid="15808" />
                    <RANKING order="3" place="3" resultid="14379" />
                    <RANKING order="4" place="-1" resultid="14926" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1126" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1127" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14824" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1128" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1129" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19310" daytime="16:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19311" daytime="16:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19312" daytime="16:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19313" daytime="16:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19314" daytime="16:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19315" daytime="16:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19316" daytime="16:35" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19317" daytime="16:35" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="19318" daytime="16:40" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1079" daytime="15:15" gender="M" number="2" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1080" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14763" />
                    <RANKING order="2" place="2" resultid="16619" />
                    <RANKING order="3" place="3" resultid="18336" />
                    <RANKING order="4" place="4" resultid="18051" />
                    <RANKING order="5" place="5" resultid="17838" />
                    <RANKING order="6" place="6" resultid="17829" />
                    <RANKING order="7" place="7" resultid="16705" />
                    <RANKING order="8" place="8" resultid="18612" />
                    <RANKING order="9" place="9" resultid="14771" />
                    <RANKING order="10" place="10" resultid="16717" />
                    <RANKING order="11" place="11" resultid="17027" />
                    <RANKING order="12" place="12" resultid="16628" />
                    <RANKING order="13" place="-1" resultid="15014" />
                    <RANKING order="14" place="-1" resultid="17279" />
                    <RANKING order="15" place="-1" resultid="18058" />
                    <RANKING order="16" place="-1" resultid="18566" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1081" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16929" />
                    <RANKING order="2" place="2" resultid="16923" />
                    <RANKING order="3" place="3" resultid="16725" />
                    <RANKING order="4" place="4" resultid="16711" />
                    <RANKING order="5" place="5" resultid="15973" />
                    <RANKING order="6" place="6" resultid="15748" />
                    <RANKING order="7" place="7" resultid="15724" />
                    <RANKING order="8" place="8" resultid="16740" />
                    <RANKING order="9" place="9" resultid="16630" />
                    <RANKING order="10" place="10" resultid="17485" />
                    <RANKING order="11" place="11" resultid="14607" />
                    <RANKING order="12" place="12" resultid="17292" />
                    <RANKING order="13" place="13" resultid="16222" />
                    <RANKING order="14" place="14" resultid="18491" />
                    <RANKING order="15" place="15" resultid="17974" />
                    <RANKING order="16" place="16" resultid="16833" />
                    <RANKING order="17" place="17" resultid="16755" />
                    <RANKING order="18" place="18" resultid="15456" />
                    <RANKING order="19" place="-1" resultid="15381" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1082" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16683" />
                    <RANKING order="2" place="2" resultid="14446" />
                    <RANKING order="3" place="3" resultid="18369" />
                    <RANKING order="4" place="4" resultid="17915" />
                    <RANKING order="5" place="5" resultid="15275" />
                    <RANKING order="6" place="6" resultid="18386" />
                    <RANKING order="7" place="7" resultid="18381" />
                    <RANKING order="8" place="8" resultid="14481" />
                    <RANKING order="9" place="9" resultid="16864" />
                    <RANKING order="10" place="10" resultid="17909" />
                    <RANKING order="11" place="11" resultid="17079" />
                    <RANKING order="12" place="12" resultid="17302" />
                    <RANKING order="13" place="13" resultid="17859" />
                    <RANKING order="14" place="14" resultid="15442" />
                    <RANKING order="15" place="15" resultid="15044" />
                    <RANKING order="16" place="16" resultid="17352" />
                    <RANKING order="17" place="17" resultid="18152" />
                    <RANKING order="18" place="18" resultid="15678" />
                    <RANKING order="19" place="19" resultid="18001" />
                    <RANKING order="20" place="20" resultid="14502" />
                    <RANKING order="21" place="21" resultid="14629" />
                    <RANKING order="22" place="22" resultid="17983" />
                    <RANKING order="23" place="-1" resultid="17696" />
                    <RANKING order="24" place="-1" resultid="18584" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1083" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15292" />
                    <RANKING order="2" place="2" resultid="17692" />
                    <RANKING order="3" place="3" resultid="17492" />
                    <RANKING order="4" place="4" resultid="17369" />
                    <RANKING order="5" place="5" resultid="16417" />
                    <RANKING order="6" place="5" resultid="17196" />
                    <RANKING order="7" place="7" resultid="16797" />
                    <RANKING order="8" place="8" resultid="16809" />
                    <RANKING order="9" place="9" resultid="16823" />
                    <RANKING order="10" place="10" resultid="17183" />
                    <RANKING order="11" place="11" resultid="14990" />
                    <RANKING order="12" place="12" resultid="16803" />
                    <RANKING order="13" place="13" resultid="17228" />
                    <RANKING order="14" place="14" resultid="16856" />
                    <RANKING order="15" place="15" resultid="16815" />
                    <RANKING order="16" place="16" resultid="17271" />
                    <RANKING order="17" place="17" resultid="17806" />
                    <RANKING order="18" place="18" resultid="16819" />
                    <RANKING order="19" place="19" resultid="16730" />
                    <RANKING order="20" place="20" resultid="17040" />
                    <RANKING order="21" place="21" resultid="16845" />
                    <RANKING order="22" place="22" resultid="17834" />
                    <RANKING order="23" place="23" resultid="16869" />
                    <RANKING order="24" place="24" resultid="16939" />
                    <RANKING order="25" place="25" resultid="16874" />
                    <RANKING order="26" place="26" resultid="16190" />
                    <RANKING order="27" place="27" resultid="16300" />
                    <RANKING order="28" place="28" resultid="16762" />
                    <RANKING order="29" place="29" resultid="16280" />
                    <RANKING order="30" place="-1" resultid="16851" />
                    <RANKING order="31" place="-1" resultid="17473" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1084" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17003" />
                    <RANKING order="2" place="2" resultid="17586" />
                    <RANKING order="3" place="3" resultid="16022" />
                    <RANKING order="4" place="4" resultid="18181" />
                    <RANKING order="5" place="5" resultid="15055" />
                    <RANKING order="6" place="6" resultid="17466" />
                    <RANKING order="7" place="7" resultid="17777" />
                    <RANKING order="8" place="8" resultid="16769" />
                    <RANKING order="9" place="9" resultid="16040" />
                    <RANKING order="10" place="10" resultid="14420" />
                    <RANKING order="11" place="11" resultid="17862" />
                    <RANKING order="12" place="12" resultid="14953" />
                    <RANKING order="13" place="13" resultid="17403" />
                    <RANKING order="14" place="14" resultid="18174" />
                    <RANKING order="15" place="15" resultid="17953" />
                    <RANKING order="16" place="16" resultid="16049" />
                    <RANKING order="17" place="17" resultid="16836" />
                    <RANKING order="18" place="18" resultid="16688" />
                    <RANKING order="19" place="19" resultid="14721" />
                    <RANKING order="20" place="20" resultid="17397" />
                    <RANKING order="21" place="21" resultid="16586" />
                    <RANKING order="22" place="22" resultid="18190" />
                    <RANKING order="23" place="23" resultid="16933" />
                    <RANKING order="24" place="24" resultid="15451" />
                    <RANKING order="25" place="-1" resultid="15343" />
                    <RANKING order="26" place="-1" resultid="15356" />
                    <RANKING order="27" place="-1" resultid="16316" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1085" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18414" />
                    <RANKING order="2" place="2" resultid="17614" />
                    <RANKING order="3" place="3" resultid="17608" />
                    <RANKING order="4" place="4" resultid="18446" />
                    <RANKING order="5" place="5" resultid="14860" />
                    <RANKING order="6" place="6" resultid="17669" />
                    <RANKING order="7" place="7" resultid="16031" />
                    <RANKING order="8" place="8" resultid="17563" />
                    <RANKING order="9" place="9" resultid="15987" />
                    <RANKING order="10" place="10" resultid="17623" />
                    <RANKING order="11" place="11" resultid="16083" />
                    <RANKING order="12" place="12" resultid="14705" />
                    <RANKING order="13" place="13" resultid="18138" />
                    <RANKING order="14" place="14" resultid="14284" />
                    <RANKING order="15" place="-1" resultid="14895" />
                    <RANKING order="16" place="-1" resultid="16079" />
                    <RANKING order="17" place="-1" resultid="16236" />
                    <RANKING order="18" place="-1" resultid="16983" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1086" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14297" />
                    <RANKING order="2" place="2" resultid="18455" />
                    <RANKING order="3" place="3" resultid="15923" />
                    <RANKING order="4" place="4" resultid="17337" />
                    <RANKING order="5" place="5" resultid="17678" />
                    <RANKING order="6" place="6" resultid="18507" />
                    <RANKING order="7" place="7" resultid="14907" />
                    <RANKING order="8" place="8" resultid="15210" />
                    <RANKING order="9" place="9" resultid="18534" />
                    <RANKING order="10" place="10" resultid="18293" />
                    <RANKING order="11" place="11" resultid="18274" />
                    <RANKING order="12" place="12" resultid="15008" />
                    <RANKING order="13" place="13" resultid="18547" />
                    <RANKING order="14" place="14" resultid="16124" />
                    <RANKING order="15" place="15" resultid="16411" />
                    <RANKING order="16" place="16" resultid="15942" />
                    <RANKING order="17" place="17" resultid="16429" />
                    <RANKING order="18" place="18" resultid="16944" />
                    <RANKING order="19" place="-1" resultid="17220" />
                    <RANKING order="20" place="-1" resultid="14618" />
                    <RANKING order="21" place="-1" resultid="15005" />
                    <RANKING order="22" place="-1" resultid="16989" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1087" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15740" />
                    <RANKING order="2" place="2" resultid="14922" />
                    <RANKING order="3" place="3" resultid="18212" />
                    <RANKING order="4" place="4" resultid="18318" />
                    <RANKING order="5" place="5" resultid="16362" />
                    <RANKING order="6" place="6" resultid="16227" />
                    <RANKING order="7" place="7" resultid="14512" />
                    <RANKING order="8" place="8" resultid="15270" />
                    <RANKING order="9" place="9" resultid="17308" />
                    <RANKING order="10" place="10" resultid="16321" />
                    <RANKING order="11" place="-1" resultid="15771" />
                    <RANKING order="12" place="-1" resultid="15361" />
                    <RANKING order="13" place="-1" resultid="17317" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1088" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17409" />
                    <RANKING order="2" place="2" resultid="17572" />
                    <RANKING order="3" place="3" resultid="14273" />
                    <RANKING order="4" place="4" resultid="14437" />
                    <RANKING order="5" place="5" resultid="15396" />
                    <RANKING order="6" place="6" resultid="18633" />
                    <RANKING order="7" place="7" resultid="18961" />
                    <RANKING order="8" place="8" resultid="16700" />
                    <RANKING order="9" place="9" resultid="15935" />
                    <RANKING order="10" place="10" resultid="16182" />
                    <RANKING order="11" place="11" resultid="15254" />
                    <RANKING order="12" place="12" resultid="16252" />
                    <RANKING order="13" place="13" resultid="16244" />
                    <RANKING order="14" place="14" resultid="16421" />
                    <RANKING order="15" place="-1" resultid="14666" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1089" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14700" />
                    <RANKING order="2" place="2" resultid="17107" />
                    <RANKING order="3" place="3" resultid="18265" />
                    <RANKING order="4" place="4" resultid="14521" />
                    <RANKING order="5" place="5" resultid="14742" />
                    <RANKING order="6" place="6" resultid="15801" />
                    <RANKING order="7" place="7" resultid="18520" />
                    <RANKING order="8" place="8" resultid="17732" />
                    <RANKING order="9" place="9" resultid="14463" />
                    <RANKING order="10" place="10" resultid="17602" />
                    <RANKING order="11" place="11" resultid="14851" />
                    <RANKING order="12" place="12" resultid="16384" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1090" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14357" />
                    <RANKING order="2" place="2" resultid="15263" />
                    <RANKING order="3" place="3" resultid="18329" />
                    <RANKING order="4" place="4" resultid="14411" />
                    <RANKING order="5" place="5" resultid="16453" />
                    <RANKING order="6" place="-1" resultid="17072" />
                    <RANKING order="7" place="-1" resultid="17283" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1091" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15807" />
                    <RANKING order="2" place="2" resultid="16177" />
                    <RANKING order="3" place="3" resultid="16442" />
                    <RANKING order="4" place="4" resultid="14378" />
                    <RANKING order="5" place="-1" resultid="17061" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1092" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15762" />
                    <RANKING order="2" place="2" resultid="18297" />
                    <RANKING order="3" place="-1" resultid="17068" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1093" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14823" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1095" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19284" daytime="15:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19285" daytime="15:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19286" daytime="15:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19287" daytime="15:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19288" daytime="15:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19289" daytime="15:25" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19290" daytime="15:25" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19291" daytime="15:25" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="19292" daytime="15:25" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="19293" daytime="15:30" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="19294" daytime="15:30" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="19295" daytime="15:30" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="19296" daytime="15:35" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="19297" daytime="15:35" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="19298" daytime="15:35" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="19299" daytime="15:35" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="19300" daytime="15:40" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="19301" daytime="15:40" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="19302" daytime="15:40" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="19303" daytime="15:40" number="20" order="20" status="OFFICIAL" />
                <HEAT heatid="19304" daytime="15:45" number="21" order="21" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1165" daytime="19:05" gender="F" number="8" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="19657" agemax="24" agemin="20" />
                <AGEGROUP agegroupid="19658" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="19659" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14869" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19660" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="19661" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17388" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19662" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="19663" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18104" />
                    <RANKING order="2" place="2" resultid="17203" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19664" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17813" />
                    <RANKING order="2" place="2" resultid="16148" />
                    <RANKING order="3" place="3" resultid="18430" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19665" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14370" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19666" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="19667" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14478" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19668" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="19669" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="19670" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="19671" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="19672" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19624" daytime="19:05" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="14207" daytime="20:05" gender="M" number="9" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="19673" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16267" />
                    <RANKING order="2" place="-1" resultid="16260" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19674" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16693" />
                    <RANKING order="2" place="2" resultid="14988" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19675" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17084" />
                    <RANKING order="2" place="2" resultid="15679" />
                    <RANKING order="3" place="-1" resultid="14630" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19676" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17578" />
                    <RANKING order="2" place="-1" resultid="15333" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19677" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16527" />
                    <RANKING order="2" place="2" resultid="14636" />
                    <RANKING order="3" place="3" resultid="14366" />
                    <RANKING order="4" place="4" resultid="17758" />
                    <RANKING order="5" place="5" resultid="16050" />
                    <RANKING order="6" place="-1" resultid="14783" />
                    <RANKING order="7" place="-1" resultid="18191" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19678" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16133" />
                    <RANKING order="2" place="2" resultid="14694" />
                    <RANKING order="3" place="-1" resultid="14896" />
                    <RANKING order="4" place="-1" resultid="16084" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19679" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16995" />
                    <RANKING order="2" place="2" resultid="18275" />
                    <RANKING order="3" place="3" resultid="18111" />
                    <RANKING order="4" place="4" resultid="16412" />
                    <RANKING order="5" place="5" resultid="17146" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19680" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15772" />
                    <RANKING order="2" place="2" resultid="14349" />
                    <RANKING order="3" place="3" resultid="18116" />
                    <RANKING order="4" place="4" resultid="14977" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19681" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14749" />
                    <RANKING order="2" place="2" resultid="14395" />
                    <RANKING order="3" place="3" resultid="18634" />
                    <RANKING order="4" place="4" resultid="18629" />
                    <RANKING order="5" place="5" resultid="18962" />
                    <RANKING order="6" place="6" resultid="14433" />
                    <RANKING order="7" place="-1" resultid="14667" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19682" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14743" />
                    <RANKING order="2" place="-1" resultid="14852" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19683" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16331" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19684" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19685" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="19686" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="19687" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="19688" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19620" daytime="20:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19621" daytime="20:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19622" daytime="21:10" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1062" daytime="15:00" gender="F" number="1" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1064" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16579" />
                    <RANKING order="2" place="2" resultid="17902" />
                    <RANKING order="3" place="3" resultid="14611" />
                    <RANKING order="4" place="4" resultid="14876" />
                    <RANKING order="5" place="5" resultid="16538" />
                    <RANKING order="6" place="6" resultid="18199" />
                    <RANKING order="7" place="7" resultid="16593" />
                    <RANKING order="8" place="8" resultid="14790" />
                    <RANKING order="9" place="-1" resultid="16636" />
                    <RANKING order="10" place="-1" resultid="18575" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16748" />
                    <RANKING order="2" place="2" resultid="14834" />
                    <RANKING order="3" place="3" resultid="15230" />
                    <RANKING order="4" place="4" resultid="17377" />
                    <RANKING order="5" place="5" resultid="17854" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14997" />
                    <RANKING order="2" place="2" resultid="17031" />
                    <RANKING order="3" place="3" resultid="17425" />
                    <RANKING order="4" place="4" resultid="14777" />
                    <RANKING order="5" place="5" resultid="16598" />
                    <RANKING order="6" place="6" resultid="17686" />
                    <RANKING order="7" place="7" resultid="15427" />
                    <RANKING order="8" place="8" resultid="18352" />
                    <RANKING order="9" place="9" resultid="16917" />
                    <RANKING order="10" place="10" resultid="18423" />
                    <RANKING order="11" place="11" resultid="14755" />
                    <RANKING order="12" place="-1" resultid="18953" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14588" />
                    <RANKING order="2" place="2" resultid="14713" />
                    <RANKING order="3" place="3" resultid="16830" />
                    <RANKING order="4" place="4" resultid="17644" />
                    <RANKING order="5" place="5" resultid="18132" />
                    <RANKING order="6" place="6" resultid="16058" />
                    <RANKING order="7" place="7" resultid="15873" />
                    <RANKING order="8" place="8" resultid="15412" />
                    <RANKING order="9" place="9" resultid="17851" />
                    <RANKING order="10" place="-1" resultid="15417" />
                    <RANKING order="11" place="-1" resultid="16165" />
                    <RANKING order="12" place="-1" resultid="16999" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1068" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16014" />
                    <RANKING order="2" place="2" resultid="15346" />
                    <RANKING order="3" place="3" resultid="14281" />
                    <RANKING order="4" place="4" resultid="17461" />
                    <RANKING order="5" place="5" resultid="14940" />
                    <RANKING order="6" place="6" resultid="17771" />
                    <RANKING order="7" place="7" resultid="17800" />
                    <RANKING order="8" place="8" resultid="18089" />
                    <RANKING order="9" place="9" resultid="14889" />
                    <RANKING order="10" place="10" resultid="18144" />
                    <RANKING order="11" place="11" resultid="16612" />
                    <RANKING order="12" place="12" resultid="16976" />
                    <RANKING order="13" place="13" resultid="16292" />
                    <RANKING order="14" place="-1" resultid="15422" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16460" />
                    <RANKING order="2" place="2" resultid="14678" />
                    <RANKING order="3" place="3" resultid="15199" />
                    <RANKING order="4" place="4" resultid="17556" />
                    <RANKING order="5" place="5" resultid="16370" />
                    <RANKING order="6" place="6" resultid="16378" />
                    <RANKING order="7" place="7" resultid="16288" />
                    <RANKING order="8" place="8" resultid="15930" />
                    <RANKING order="9" place="9" resultid="15945" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16309" />
                    <RANKING order="2" place="2" resultid="17596" />
                    <RANKING order="3" place="3" resultid="18103" />
                    <RANKING order="4" place="4" resultid="15064" />
                    <RANKING order="5" place="5" resultid="16531" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15223" />
                    <RANKING order="2" place="2" resultid="16465" />
                    <RANKING order="3" place="3" resultid="16147" />
                    <RANKING order="4" place="4" resultid="17548" />
                    <RANKING order="5" place="5" resultid="17619" />
                    <RANKING order="6" place="6" resultid="16156" />
                    <RANKING order="7" place="7" resultid="14486" />
                    <RANKING order="8" place="8" resultid="16348" />
                    <RANKING order="9" place="9" resultid="16296" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1072" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17153" />
                    <RANKING order="2" place="2" resultid="16387" />
                    <RANKING order="3" place="3" resultid="17628" />
                    <RANKING order="4" place="4" resultid="17091" />
                    <RANKING order="5" place="5" resultid="14843" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1073" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15204" />
                    <RANKING order="2" place="2" resultid="17723" />
                    <RANKING order="3" place="3" resultid="14492" />
                    <RANKING order="4" place="4" resultid="17639" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1074" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14457" />
                    <RANKING order="2" place="2" resultid="16339" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1075" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1076" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1077" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18309" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1078" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1063" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19275" daytime="15:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19276" daytime="15:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19277" daytime="15:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19278" daytime="15:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19279" daytime="15:05" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19280" daytime="15:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19281" daytime="15:10" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19282" daytime="15:10" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="19283" daytime="15:15" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="19612" daytime="17:00" gender="F" number="6" order="7" round="FHT" preveventid="1147">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="19596" daytime="17:00" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="19610" daytime="17:50" gender="M" number="7" order="9" round="FHT" preveventid="14189">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="19618" daytime="17:50" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1096" daytime="15:45" gender="F" number="3" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1097" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17233" />
                    <RANKING order="2" place="2" resultid="17941" />
                    <RANKING order="3" place="3" resultid="15729" />
                    <RANKING order="4" place="4" resultid="18159" />
                    <RANKING order="5" place="5" resultid="14791" />
                    <RANKING order="6" place="6" resultid="16539" />
                    <RANKING order="7" place="-1" resultid="15405" />
                    <RANKING order="8" place="-1" resultid="18576" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14835" />
                    <RANKING order="2" place="2" resultid="17591" />
                    <RANKING order="3" place="3" resultid="18410" />
                    <RANKING order="4" place="-1" resultid="17506" />
                    <RANKING order="5" place="-1" resultid="14645" />
                    <RANKING order="6" place="-1" resultid="18094" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1099" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14998" />
                    <RANKING order="2" place="2" resultid="17032" />
                    <RANKING order="3" place="3" resultid="17785" />
                    <RANKING order="4" place="4" resultid="17708" />
                    <RANKING order="5" place="5" resultid="18360" />
                    <RANKING order="6" place="6" resultid="17961" />
                    <RANKING order="7" place="7" resultid="17479" />
                    <RANKING order="8" place="-1" resultid="18481" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1100" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14589" />
                    <RANKING order="2" place="2" resultid="17927" />
                    <RANKING order="3" place="3" resultid="14714" />
                    <RANKING order="4" place="4" resultid="16059" />
                    <RANKING order="5" place="5" resultid="18133" />
                    <RANKING order="6" place="6" resultid="15949" />
                    <RANKING order="7" place="7" resultid="15874" />
                    <RANKING order="8" place="8" resultid="16284" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1101" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15282" />
                    <RANKING order="2" place="2" resultid="14282" />
                    <RANKING order="3" place="3" resultid="15882" />
                    <RANKING order="4" place="-1" resultid="17632" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15236" />
                    <RANKING order="2" place="2" resultid="18514" />
                    <RANKING order="3" place="3" resultid="17328" />
                    <RANKING order="4" place="4" resultid="17098" />
                    <RANKING order="5" place="5" resultid="16379" />
                    <RANKING order="6" place="-1" resultid="14807" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1103" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16399" />
                    <RANKING order="2" place="2" resultid="15065" />
                    <RANKING order="3" place="3" resultid="16532" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1104" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18621" />
                    <RANKING order="2" place="2" resultid="14686" />
                    <RANKING order="3" place="3" resultid="17549" />
                    <RANKING order="4" place="4" resultid="18429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1105" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14623" />
                    <RANKING order="2" place="2" resultid="14369" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1106" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17724" />
                    <RANKING order="2" place="2" resultid="16405" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1107" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16340" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1108" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1109" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1110" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1111" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1112" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19305" daytime="15:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19306" daytime="15:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19307" daytime="15:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19308" daytime="16:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19309" daytime="16:05" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2017-11-18" daytime="09:00" endtime="12:24" name="BLOK II" number="2" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="1341" daytime="12:35" gender="M" number="19" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1342" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17324" />
                    <RANKING order="2" place="2" resultid="18615" />
                    <RANKING order="3" place="-1" resultid="18060" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1343" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16694" />
                    <RANKING order="2" place="2" resultid="18501" />
                    <RANKING order="3" place="3" resultid="15891" />
                    <RANKING order="4" place="4" resultid="14672" />
                    <RANKING order="5" place="5" resultid="15390" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1344" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15899" />
                    <RANKING order="2" place="2" resultid="18587" />
                    <RANKING order="3" place="3" resultid="18126" />
                    <RANKING order="4" place="4" resultid="15045" />
                    <RANKING order="5" place="-1" resultid="16881" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1345" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17172" />
                    <RANKING order="2" place="2" resultid="15907" />
                    <RANKING order="3" place="3" resultid="17705" />
                    <RANKING order="4" place="4" resultid="17457" />
                    <RANKING order="5" place="-1" resultid="16799" />
                    <RANKING order="6" place="-1" resultid="17042" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1346" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15058" />
                    <RANKING order="2" place="2" resultid="16971" />
                    <RANKING order="3" place="3" resultid="16528" />
                    <RANKING order="4" place="4" resultid="17794" />
                    <RANKING order="5" place="5" resultid="16052" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1347" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17610" />
                    <RANKING order="2" place="2" resultid="14695" />
                    <RANKING order="3" place="3" resultid="16075" />
                    <RANKING order="4" place="4" resultid="15039" />
                    <RANKING order="5" place="5" resultid="18222" />
                    <RANKING order="6" place="6" resultid="16094" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1348" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17147" />
                    <RANKING order="2" place="2" resultid="17392" />
                    <RANKING order="3" place="3" resultid="15859" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1349" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15743" />
                    <RANKING order="2" place="2" resultid="18215" />
                    <RANKING order="3" place="3" resultid="14350" />
                    <RANKING order="4" place="4" resultid="16230" />
                    <RANKING order="5" place="-1" resultid="14978" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1350" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15248" />
                    <RANKING order="2" place="2" resultid="14729" />
                    <RANKING order="3" place="3" resultid="14397" />
                    <RANKING order="4" place="4" resultid="18964" />
                    <RANKING order="5" place="5" resultid="15257" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1351" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18268" />
                    <RANKING order="2" place="2" resultid="17142" />
                    <RANKING order="3" place="3" resultid="15826" />
                    <RANKING order="4" place="4" resultid="14658" />
                    <RANKING order="5" place="-1" resultid="17055" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1352" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14565" />
                    <RANKING order="2" place="2" resultid="15265" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1353" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14290" />
                    <RANKING order="2" place="2" resultid="14381" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1354" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1355" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1356" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1357" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19413" daytime="12:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19414" daytime="12:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19415" daytime="12:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19416" daytime="12:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19417" daytime="12:55" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19418" daytime="13:00" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1239" daytime="10:00" gender="M" number="13" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1240" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16214" />
                    <RANKING order="2" place="2" resultid="18595" />
                    <RANKING order="3" place="3" resultid="15017" />
                    <RANKING order="4" place="4" resultid="18955" />
                    <RANKING order="5" place="5" resultid="16261" />
                    <RANKING order="6" place="-1" resultid="18569" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1241" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18492" />
                    <RANKING order="2" place="2" resultid="15890" />
                    <RANKING order="3" place="3" resultid="15389" />
                    <RANKING order="4" place="-1" resultid="14268" />
                    <RANKING order="5" place="-1" resultid="14671" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1242" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17304" />
                    <RANKING order="2" place="2" resultid="17085" />
                    <RANKING order="3" place="3" resultid="15444" />
                    <RANKING order="4" place="4" resultid="18125" />
                    <RANKING order="5" place="5" resultid="18002" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1243" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17171" />
                    <RANKING order="2" place="2" resultid="17184" />
                    <RANKING order="3" place="3" resultid="16804" />
                    <RANKING order="4" place="4" resultid="17807" />
                    <RANKING order="5" place="5" resultid="14553" />
                    <RANKING order="6" place="-1" resultid="14883" />
                    <RANKING order="7" place="-1" resultid="15906" />
                    <RANKING order="8" place="-1" resultid="16858" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1244" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18555" />
                    <RANKING order="2" place="2" resultid="18418" />
                    <RANKING order="3" place="3" resultid="16042" />
                    <RANKING order="4" place="4" resultid="16317" />
                    <RANKING order="5" place="5" resultid="14277" />
                    <RANKING order="6" place="6" resultid="17404" />
                    <RANKING order="7" place="7" resultid="17543" />
                    <RANKING order="8" place="8" resultid="17501" />
                    <RANKING order="9" place="-1" resultid="14784" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1245" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14966" />
                    <RANKING order="2" place="2" resultid="16068" />
                    <RANKING order="3" place="3" resultid="16033" />
                    <RANKING order="4" place="4" resultid="14862" />
                    <RANKING order="5" place="5" resultid="14707" />
                    <RANKING order="6" place="6" resultid="18139" />
                    <RANKING order="7" place="7" resultid="17365" />
                    <RANKING order="8" place="-1" resultid="16237" />
                    <RANKING order="9" place="-1" resultid="16396" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1246" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16474" />
                    <RANKING order="2" place="2" resultid="17391" />
                    <RANKING order="3" place="3" resultid="15858" />
                    <RANKING order="4" place="4" resultid="16432" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1247" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18283" />
                    <RANKING order="2" place="2" resultid="18468" />
                    <RANKING order="3" place="3" resultid="17179" />
                    <RANKING order="4" place="4" resultid="15784" />
                    <RANKING order="5" place="5" resultid="18117" />
                    <RANKING order="6" place="6" resultid="16323" />
                    <RANKING order="7" place="-1" resultid="15278" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1248" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14728" />
                    <RANKING order="2" place="2" resultid="15398" />
                    <RANKING order="3" place="3" resultid="15821" />
                    <RANKING order="4" place="4" resultid="16423" />
                    <RANKING order="5" place="-1" resultid="18438" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1249" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17450" />
                    <RANKING order="2" place="2" resultid="15217" />
                    <RANKING order="3" place="3" resultid="14657" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1250" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14359" />
                    <RANKING order="2" place="2" resultid="14413" />
                    <RANKING order="3" place="-1" resultid="17074" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1251" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14474" />
                    <RANKING order="2" place="2" resultid="14289" />
                    <RANKING order="3" place="3" resultid="14928" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1252" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="18299" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1253" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1254" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1255" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19359" daytime="10:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19360" daytime="10:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19361" daytime="10:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19362" daytime="10:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19363" daytime="10:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19364" daytime="10:25" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19365" daytime="10:25" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1381" daytime="13:10" gender="M" number="21" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="16653" agemax="99" agemin="80" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17875" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16654" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16952" />
                    <RANKING order="2" place="2" resultid="16774" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16655" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18402" />
                    <RANKING order="2" place="2" resultid="17242" />
                    <RANKING order="3" place="3" resultid="16888" />
                    <RANKING order="4" place="4" resultid="17514" />
                    <RANKING order="5" place="5" resultid="18230" />
                    <RANKING order="6" place="6" resultid="17120" />
                    <RANKING order="7" place="7" resultid="14954" />
                    <RANKING order="8" place="8" resultid="17873" />
                    <RANKING order="9" place="9" resultid="18016" />
                    <RANKING order="10" place="10" resultid="16889" />
                    <RANKING order="11" place="11" resultid="16890" />
                    <RANKING order="12" place="12" resultid="16776" />
                    <RANKING order="13" place="-1" resultid="16640" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16656" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17515" />
                    <RANKING order="2" place="2" resultid="17654" />
                    <RANKING order="3" place="3" resultid="16091" />
                    <RANKING order="4" place="4" resultid="16484" />
                    <RANKING order="5" place="4" resultid="17874" />
                    <RANKING order="6" place="6" resultid="15997" />
                    <RANKING order="7" place="7" resultid="16092" />
                    <RANKING order="8" place="8" resultid="18232" />
                    <RANKING order="9" place="9" resultid="18018" />
                    <RANKING order="10" place="-1" resultid="15308" />
                    <RANKING order="11" place="-1" resultid="18542" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16657" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17243" />
                    <RANKING order="2" place="2" resultid="18234" />
                    <RANKING order="3" place="3" resultid="16211" />
                    <RANKING order="4" place="-1" resultid="16210" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16658" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15310" />
                    <RANKING order="2" place="2" resultid="15969" />
                    <RANKING order="3" place="3" resultid="14902" />
                    <RANKING order="4" place="4" resultid="16485" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16659" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14535" />
                    <RANKING order="2" place="2" resultid="15830" />
                    <RANKING order="3" place="3" resultid="17115" />
                    <RANKING order="4" place="4" resultid="16486" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19421" daytime="13:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19422" daytime="13:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19423" daytime="13:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19424" daytime="13:20" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1273" daytime="10:50" gender="M" number="15" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1274" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16621" />
                    <RANKING order="2" place="2" resultid="18596" />
                    <RANKING order="3" place="3" resultid="17831" />
                    <RANKING order="4" place="4" resultid="14764" />
                    <RANKING order="5" place="5" resultid="17840" />
                    <RANKING order="6" place="6" resultid="16268" />
                    <RANKING order="7" place="7" resultid="17139" />
                    <RANKING order="8" place="8" resultid="16719" />
                    <RANKING order="9" place="9" resultid="17028" />
                    <RANKING order="10" place="10" resultid="17968" />
                    <RANKING order="11" place="-1" resultid="15049" />
                    <RANKING order="12" place="-1" resultid="18059" />
                    <RANKING order="13" place="-1" resultid="18339" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1275" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17486" />
                    <RANKING order="2" place="2" resultid="15725" />
                    <RANKING order="3" place="3" resultid="15750" />
                    <RANKING order="4" place="4" resultid="15974" />
                    <RANKING order="5" place="5" resultid="14608" />
                    <RANKING order="6" place="6" resultid="14603" />
                    <RANKING order="7" place="7" resultid="17976" />
                    <RANKING order="8" place="8" resultid="16756" />
                    <RANKING order="9" place="9" resultid="17997" />
                    <RANKING order="10" place="10" resultid="15457" />
                    <RANKING order="11" place="-1" resultid="15437" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1276" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16685" />
                    <RANKING order="2" place="2" resultid="14448" />
                    <RANKING order="3" place="3" resultid="18370" />
                    <RANKING order="4" place="4" resultid="17916" />
                    <RANKING order="5" place="5" resultid="18389" />
                    <RANKING order="6" place="6" resultid="18382" />
                    <RANKING order="7" place="7" resultid="17080" />
                    <RANKING order="8" place="8" resultid="17910" />
                    <RANKING order="9" place="9" resultid="17860" />
                    <RANKING order="10" place="10" resultid="16866" />
                    <RANKING order="11" place="11" resultid="18155" />
                    <RANKING order="12" place="12" resultid="16736" />
                    <RANKING order="13" place="13" resultid="14504" />
                    <RANKING order="14" place="14" resultid="14631" />
                    <RANKING order="15" place="15" resultid="17937" />
                    <RANKING order="16" place="16" resultid="17985" />
                    <RANKING order="17" place="-1" resultid="14482" />
                    <RANKING order="18" place="-1" resultid="17697" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1277" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16203" />
                    <RANKING order="2" place="2" resultid="17493" />
                    <RANKING order="3" place="3" resultid="16825" />
                    <RANKING order="4" place="4" resultid="17197" />
                    <RANKING order="5" place="5" resultid="16798" />
                    <RANKING order="6" place="6" resultid="17579" />
                    <RANKING order="7" place="7" resultid="17185" />
                    <RANKING order="8" place="8" resultid="17229" />
                    <RANKING order="9" place="9" resultid="18207" />
                    <RANKING order="10" place="10" resultid="17456" />
                    <RANKING order="11" place="11" resultid="17041" />
                    <RANKING order="12" place="12" resultid="16731" />
                    <RANKING order="13" place="13" resultid="17808" />
                    <RANKING order="14" place="14" resultid="18463" />
                    <RANKING order="15" place="15" resultid="15334" />
                    <RANKING order="16" place="16" resultid="16940" />
                    <RANKING order="17" place="17" resultid="16281" />
                    <RANKING order="18" place="18" resultid="16763" />
                    <RANKING order="19" place="19" resultid="16301" />
                    <RANKING order="20" place="-1" resultid="16172" />
                    <RANKING order="21" place="-1" resultid="16418" />
                    <RANKING order="22" place="-1" resultid="16816" />
                    <RANKING order="23" place="-1" resultid="16852" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1278" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18183" />
                    <RANKING order="2" place="2" resultid="17587" />
                    <RANKING order="3" place="3" resultid="15057" />
                    <RANKING order="4" place="4" resultid="16024" />
                    <RANKING order="5" place="5" resultid="17004" />
                    <RANKING order="6" place="6" resultid="17009" />
                    <RANKING order="7" place="7" resultid="16770" />
                    <RANKING order="8" place="8" resultid="17778" />
                    <RANKING order="9" place="9" resultid="17863" />
                    <RANKING order="10" place="10" resultid="16051" />
                    <RANKING order="11" place="11" resultid="17954" />
                    <RANKING order="12" place="12" resultid="14263" />
                    <RANKING order="13" place="13" resultid="17502" />
                    <RANKING order="14" place="14" resultid="16588" />
                    <RANKING order="15" place="15" resultid="18193" />
                    <RANKING order="16" place="16" resultid="14722" />
                    <RANKING order="17" place="17" resultid="17398" />
                    <RANKING order="18" place="18" resultid="16935" />
                    <RANKING order="19" place="19" resultid="17923" />
                    <RANKING order="20" place="-1" resultid="15344" />
                    <RANKING order="21" place="-1" resultid="15452" />
                    <RANKING order="22" place="-1" resultid="16839" />
                    <RANKING order="23" place="-1" resultid="17971" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1279" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17615" />
                    <RANKING order="2" place="2" resultid="18562" />
                    <RANKING order="3" place="3" resultid="17609" />
                    <RANKING order="4" place="4" resultid="17671" />
                    <RANKING order="5" place="5" resultid="15038" />
                    <RANKING order="6" place="6" resultid="17624" />
                    <RANKING order="7" place="7" resultid="17565" />
                    <RANKING order="8" place="8" resultid="14897" />
                    <RANKING order="9" place="9" resultid="17366" />
                    <RANKING order="10" place="10" resultid="17994" />
                    <RANKING order="11" place="11" resultid="16397" />
                    <RANKING order="12" place="-1" resultid="14863" />
                    <RANKING order="13" place="-1" resultid="16097" />
                    <RANKING order="14" place="-1" resultid="16238" />
                    <RANKING order="15" place="-1" resultid="18007" />
                    <RANKING order="16" place="-1" resultid="16985" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1280" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18457" />
                    <RANKING order="2" place="2" resultid="18536" />
                    <RANKING order="3" place="3" resultid="17680" />
                    <RANKING order="4" place="4" resultid="15925" />
                    <RANKING order="5" place="5" resultid="14909" />
                    <RANKING order="6" place="6" resultid="15211" />
                    <RANKING order="7" place="7" resultid="18277" />
                    <RANKING order="8" place="8" resultid="16126" />
                    <RANKING order="9" place="9" resultid="15759" />
                    <RANKING order="10" place="10" resultid="16475" />
                    <RANKING order="11" place="11" resultid="18112" />
                    <RANKING order="12" place="12" resultid="15193" />
                    <RANKING order="13" place="13" resultid="15943" />
                    <RANKING order="14" place="-1" resultid="18548" />
                    <RANKING order="15" place="-1" resultid="16991" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1281" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17215" />
                    <RANKING order="2" place="2" resultid="14923" />
                    <RANKING order="3" place="3" resultid="15774" />
                    <RANKING order="4" place="4" resultid="14514" />
                    <RANKING order="5" place="5" resultid="15271" />
                    <RANKING order="6" place="6" resultid="17311" />
                    <RANKING order="7" place="7" resultid="15919" />
                    <RANKING order="8" place="-1" resultid="15362" />
                    <RANKING order="9" place="-1" resultid="17318" />
                    <RANKING order="10" place="-1" resultid="18319" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1282" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17411" />
                    <RANKING order="2" place="2" resultid="14274" />
                    <RANKING order="3" place="3" resultid="14440" />
                    <RANKING order="4" place="4" resultid="18635" />
                    <RANKING order="5" place="5" resultid="16184" />
                    <RANKING order="6" place="6" resultid="15256" />
                    <RANKING order="7" place="7" resultid="16254" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1283" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17109" />
                    <RANKING order="2" place="2" resultid="14522" />
                    <RANKING order="3" place="3" resultid="18522" />
                    <RANKING order="4" place="4" resultid="14744" />
                    <RANKING order="5" place="5" resultid="17603" />
                    <RANKING order="6" place="6" resultid="15803" />
                    <RANKING order="7" place="7" resultid="14854" />
                    <RANKING order="8" place="-1" resultid="14701" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1284" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14564" />
                    <RANKING order="2" place="2" resultid="16332" />
                    <RANKING order="3" place="3" resultid="15264" />
                    <RANKING order="4" place="4" resultid="18331" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1285" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16178" />
                    <RANKING order="2" place="2" resultid="17063" />
                    <RANKING order="3" place="3" resultid="16444" />
                    <RANKING order="4" place="4" resultid="14388" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1286" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15764" />
                    <RANKING order="2" place="2" resultid="17069" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1287" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14826" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1288" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1289" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19373" daytime="10:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19374" daytime="10:55" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19375" daytime="10:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19376" daytime="11:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19377" daytime="11:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19378" daytime="11:05" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19379" daytime="11:05" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19380" daytime="11:10" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="19381" daytime="11:10" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="19382" daytime="11:15" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="19383" daytime="11:15" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="19384" daytime="11:15" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="19385" daytime="11:20" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="19386" daytime="11:20" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="19387" daytime="11:25" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="19388" daytime="11:25" number="16" order="16" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1187" daytime="09:00" gender="F" number="10" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1189" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17903" />
                    <RANKING order="2" place="2" resultid="18600" />
                    <RANKING order="3" place="3" resultid="17942" />
                    <RANKING order="4" place="4" resultid="16607" />
                    <RANKING order="5" place="5" resultid="14612" />
                    <RANKING order="6" place="-1" resultid="15406" />
                    <RANKING order="7" place="-1" resultid="16965" />
                    <RANKING order="8" place="-1" resultid="18160" />
                    <RANKING order="9" place="-1" resultid="18577" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1190" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15231" />
                    <RANKING order="2" place="2" resultid="14830" />
                    <RANKING order="3" place="3" resultid="17507" />
                    <RANKING order="4" place="-1" resultid="14583" />
                    <RANKING order="5" place="-1" resultid="18096" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1191" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14999" />
                    <RANKING order="2" place="2" resultid="14870" />
                    <RANKING order="3" place="-1" resultid="18482" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1192" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17014" />
                    <RANKING order="2" place="2" resultid="17929" />
                    <RANKING order="3" place="3" resultid="14715" />
                    <RANKING order="4" place="4" resultid="17000" />
                    <RANKING order="5" place="5" resultid="15875" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1193" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15283" />
                    <RANKING order="2" place="2" resultid="14941" />
                    <RANKING order="3" place="3" resultid="16008" />
                    <RANKING order="4" place="4" resultid="18090" />
                    <RANKING order="5" place="5" resultid="17801" />
                    <RANKING order="6" place="6" resultid="14891" />
                    <RANKING order="7" place="7" resultid="16977" />
                    <RANKING order="8" place="8" resultid="18145" />
                    <RANKING order="9" place="9" resultid="16293" />
                    <RANKING order="10" place="-1" resultid="17633" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1194" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15237" />
                    <RANKING order="2" place="2" resultid="15841" />
                    <RANKING order="3" place="3" resultid="14679" />
                    <RANKING order="4" place="4" resultid="16371" />
                    <RANKING order="5" place="5" resultid="17557" />
                    <RANKING order="6" place="6" resultid="17100" />
                    <RANKING order="7" place="7" resultid="14800" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1195" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16310" />
                    <RANKING order="2" place="2" resultid="17597" />
                    <RANKING order="3" place="3" resultid="17204" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1196" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15224" />
                    <RANKING order="2" place="2" resultid="18622" />
                    <RANKING order="3" place="3" resultid="15780" />
                    <RANKING order="4" place="4" resultid="16149" />
                    <RANKING order="5" place="5" resultid="14509" />
                    <RANKING order="6" place="6" resultid="16350" />
                    <RANKING order="7" place="7" resultid="14519" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1197" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14577" />
                    <RANKING order="2" place="2" resultid="17190" />
                    <RANKING order="3" place="3" resultid="17092" />
                    <RANKING order="4" place="4" resultid="14845" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1198" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15205" />
                    <RANKING order="2" place="2" resultid="17725" />
                    <RANKING order="3" place="3" resultid="17640" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1199" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14458" />
                    <RANKING order="2" place="2" resultid="14404" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1200" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18288" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1201" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18305" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1202" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18311" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1203" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1204" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19336" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19337" daytime="09:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19338" daytime="09:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19339" daytime="09:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19340" daytime="09:05" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19341" daytime="09:10" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1324" daytime="12:20" gender="F" number="18" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1325" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18601" />
                    <RANKING order="2" place="2" resultid="14793" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1326" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="18097" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1327" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18363" />
                    <RANKING order="2" place="2" resultid="17963" />
                    <RANKING order="3" place="3" resultid="17481" />
                    <RANKING order="4" place="-1" resultid="15428" />
                    <RANKING order="5" place="-1" resultid="18483" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1328" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="1329" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15884" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1330" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16381" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1331" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="1332" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15225" />
                    <RANKING order="2" place="2" resultid="14688" />
                    <RANKING order="3" place="3" resultid="16468" />
                    <RANKING order="4" place="4" resultid="18431" />
                    <RANKING order="5" place="-1" resultid="16159" />
                    <RANKING order="6" place="-1" resultid="16351" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1333" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16390" />
                    <RANKING order="2" place="2" resultid="14372" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1334" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1335" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14479" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1336" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1337" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1338" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1339" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1340" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19411" daytime="12:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19412" daytime="12:30" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="14225" daytime="11:25" gender="F" number="16" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="14226" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16581" />
                    <RANKING order="2" place="2" resultid="17235" />
                    <RANKING order="3" place="3" resultid="15731" />
                    <RANKING order="4" place="4" resultid="17943" />
                    <RANKING order="5" place="5" resultid="16608" />
                    <RANKING order="6" place="6" resultid="17904" />
                    <RANKING order="7" place="7" resultid="18161" />
                    <RANKING order="8" place="8" resultid="14878" />
                    <RANKING order="9" place="9" resultid="16541" />
                    <RANKING order="10" place="10" resultid="16594" />
                    <RANKING order="11" place="-1" resultid="15407" />
                    <RANKING order="12" place="-1" resultid="16966" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14227" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14837" />
                    <RANKING order="2" place="2" resultid="16750" />
                    <RANKING order="3" place="3" resultid="17855" />
                    <RANKING order="4" place="4" resultid="17508" />
                    <RANKING order="5" place="5" resultid="14572" />
                    <RANKING order="6" place="-1" resultid="14648" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14228" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17034" />
                    <RANKING order="2" place="2" resultid="15000" />
                    <RANKING order="3" place="3" resultid="17787" />
                    <RANKING order="4" place="4" resultid="16600" />
                    <RANKING order="5" place="5" resultid="14778" />
                    <RANKING order="6" place="6" resultid="17962" />
                    <RANKING order="7" place="7" resultid="17361" />
                    <RANKING order="8" place="8" resultid="17427" />
                    <RANKING order="9" place="9" resultid="17687" />
                    <RANKING order="10" place="10" resultid="17480" />
                    <RANKING order="11" place="-1" resultid="17711" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14229" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17445" />
                    <RANKING order="2" place="2" resultid="14591" />
                    <RANKING order="3" place="3" resultid="14716" />
                    <RANKING order="4" place="4" resultid="17015" />
                    <RANKING order="5" place="5" resultid="17930" />
                    <RANKING order="6" place="6" resultid="15867" />
                    <RANKING order="7" place="7" resultid="17701" />
                    <RANKING order="8" place="8" resultid="15955" />
                    <RANKING order="9" place="9" resultid="15950" />
                    <RANKING order="10" place="-1" resultid="16061" />
                    <RANKING order="11" place="-1" resultid="17645" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14230" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15284" />
                    <RANKING order="2" place="2" resultid="15883" />
                    <RANKING order="3" place="3" resultid="16016" />
                    <RANKING order="4" place="4" resultid="17462" />
                    <RANKING order="5" place="5" resultid="15348" />
                    <RANKING order="6" place="6" resultid="17389" />
                    <RANKING order="7" place="7" resultid="18091" />
                    <RANKING order="8" place="8" resultid="16978" />
                    <RANKING order="9" place="-1" resultid="17634" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14231" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15238" />
                    <RANKING order="2" place="2" resultid="14680" />
                    <RANKING order="3" place="3" resultid="17559" />
                    <RANKING order="4" place="4" resultid="17331" />
                    <RANKING order="5" place="5" resultid="17101" />
                    <RANKING order="6" place="6" resultid="14810" />
                    <RANKING order="7" place="7" resultid="14801" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14232" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16311" />
                    <RANKING order="2" place="2" resultid="17598" />
                    <RANKING order="3" place="3" resultid="16400" />
                    <RANKING order="4" place="4" resultid="15067" />
                    <RANKING order="5" place="5" resultid="16534" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14233" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18623" />
                    <RANKING order="2" place="2" resultid="17551" />
                    <RANKING order="3" place="3" resultid="17815" />
                    <RANKING order="4" place="4" resultid="16150" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14234" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17155" />
                    <RANKING order="2" place="2" resultid="17629" />
                    <RANKING order="3" place="3" resultid="14624" />
                    <RANKING order="4" place="4" resultid="14578" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14235" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17641" />
                    <RANKING order="2" place="2" resultid="16406" />
                    <RANKING order="3" place="3" resultid="15027" />
                    <RANKING order="4" place="-1" resultid="17437" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14236" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14467" />
                    <RANKING order="2" place="2" resultid="16342" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14237" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18289" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14238" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="14239" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="14240" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="14241" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19389" daytime="11:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19390" daytime="11:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19391" daytime="11:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19392" daytime="11:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19393" daytime="11:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19394" daytime="11:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19395" daytime="11:45" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19396" daytime="11:45" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1222" daytime="09:30" gender="F" number="12" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1223" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17234" />
                    <RANKING order="2" place="2" resultid="15846" />
                    <RANKING order="3" place="3" resultid="18578" />
                    <RANKING order="4" place="4" resultid="14792" />
                    <RANKING order="5" place="5" resultid="14877" />
                    <RANKING order="6" place="6" resultid="18201" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1224" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14993" />
                    <RANKING order="2" place="2" resultid="17948" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1225" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17033" />
                    <RANKING order="2" place="2" resultid="18362" />
                    <RANKING order="3" place="3" resultid="17786" />
                    <RANKING order="4" place="4" resultid="17710" />
                    <RANKING order="5" place="5" resultid="15433" />
                    <RANKING order="6" place="6" resultid="18353" />
                    <RANKING order="7" place="7" resultid="14756" />
                    <RANKING order="8" place="-1" resultid="17426" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1226" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16060" />
                    <RANKING order="2" place="2" resultid="17754" />
                    <RANKING order="3" place="3" resultid="16166" />
                    <RANKING order="4" place="4" resultid="15876" />
                    <RANKING order="5" place="5" resultid="16285" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1227" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15960" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1228" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18515" />
                    <RANKING order="2" place="2" resultid="14527" />
                    <RANKING order="3" place="3" resultid="17330" />
                    <RANKING order="4" place="4" resultid="15931" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1229" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17419" />
                    <RANKING order="2" place="2" resultid="15066" />
                    <RANKING order="3" place="3" resultid="18105" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1230" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14687" />
                    <RANKING order="2" place="2" resultid="17550" />
                    <RANKING order="3" place="3" resultid="17814" />
                    <RANKING order="4" place="4" resultid="16158" />
                    <RANKING order="5" place="-1" resultid="16297" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1231" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17154" />
                    <RANKING order="2" place="2" resultid="17605" />
                    <RANKING order="3" place="3" resultid="18170" />
                    <RANKING order="4" place="4" resultid="14371" />
                    <RANKING order="5" place="5" resultid="19743" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1232" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14470" />
                    <RANKING order="2" place="2" resultid="15026" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1233" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1234" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1235" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15791" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1236" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1237" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1238" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19354" daytime="09:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19355" daytime="09:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19356" daytime="09:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19357" daytime="09:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19358" daytime="09:55" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="14243" daytime="11:50" gender="M" number="17" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="14244" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15050" />
                    <RANKING order="2" place="2" resultid="18607" />
                    <RANKING order="3" place="3" resultid="17431" />
                    <RANKING order="4" place="4" resultid="16622" />
                    <RANKING order="5" place="5" resultid="18053" />
                    <RANKING order="6" place="6" resultid="17847" />
                    <RANKING order="7" place="7" resultid="16707" />
                    <RANKING order="8" place="8" resultid="14765" />
                    <RANKING order="9" place="9" resultid="16269" />
                    <RANKING order="10" place="10" resultid="17843" />
                    <RANKING order="11" place="-1" resultid="17280" />
                    <RANKING order="12" place="-1" resultid="18340" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14245" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16713" />
                    <RANKING order="2" place="2" resultid="16743" />
                    <RANKING order="3" place="3" resultid="16726" />
                    <RANKING order="4" place="4" resultid="14269" />
                    <RANKING order="5" place="5" resultid="17487" />
                    <RANKING order="6" place="6" resultid="17825" />
                    <RANKING order="7" place="7" resultid="18167" />
                    <RANKING order="8" place="8" resultid="15975" />
                    <RANKING order="9" place="9" resultid="15751" />
                    <RANKING order="10" place="10" resultid="18518" />
                    <RANKING order="11" place="11" resultid="16632" />
                    <RANKING order="12" place="12" resultid="18493" />
                    <RANKING order="13" place="13" resultid="18348" />
                    <RANKING order="14" place="14" resultid="17977" />
                    <RANKING order="15" place="15" resultid="16757" />
                    <RANKING order="16" place="16" resultid="16277" />
                    <RANKING order="17" place="17" resultid="16142" />
                    <RANKING order="18" place="-1" resultid="16925" />
                    <RANKING order="19" place="-1" resultid="16931" />
                    <RANKING order="20" place="-1" resultid="17295" />
                    <RANKING order="21" place="-1" resultid="15383" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14246" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15898" />
                    <RANKING order="2" place="2" resultid="17917" />
                    <RANKING order="3" place="3" resultid="15445" />
                    <RANKING order="4" place="4" resultid="17355" />
                    <RANKING order="5" place="-1" resultid="16615" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14247" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18375" />
                    <RANKING order="2" place="2" resultid="17475" />
                    <RANKING order="3" place="3" resultid="15295" />
                    <RANKING order="4" place="4" resultid="17021" />
                    <RANKING order="5" place="5" resultid="17372" />
                    <RANKING order="6" place="6" resultid="17494" />
                    <RANKING order="7" place="7" resultid="17198" />
                    <RANKING order="8" place="8" resultid="16419" />
                    <RANKING order="9" place="9" resultid="14991" />
                    <RANKING order="10" place="10" resultid="17580" />
                    <RANKING order="11" place="11" resultid="17049" />
                    <RANKING order="12" place="12" resultid="17274" />
                    <RANKING order="13" place="13" resultid="16192" />
                    <RANKING order="14" place="14" resultid="16810" />
                    <RANKING order="15" place="15" resultid="17714" />
                    <RANKING order="16" place="16" resultid="16847" />
                    <RANKING order="17" place="17" resultid="16732" />
                    <RANKING order="18" place="18" resultid="18464" />
                    <RANKING order="19" place="19" resultid="14554" />
                    <RANKING order="20" place="20" resultid="16764" />
                    <RANKING order="21" place="21" resultid="16358" />
                    <RANKING order="22" place="-1" resultid="14817" />
                    <RANKING order="23" place="-1" resultid="14884" />
                    <RANKING order="24" place="-1" resultid="16870" />
                    <RANKING order="25" place="-1" resultid="16875" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14248" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18556" />
                    <RANKING order="2" place="2" resultid="17821" />
                    <RANKING order="3" place="3" resultid="16025" />
                    <RANKING order="4" place="4" resultid="18047" />
                    <RANKING order="5" place="5" resultid="18184" />
                    <RANKING order="6" place="6" resultid="18529" />
                    <RANKING order="7" place="7" resultid="18419" />
                    <RANKING order="8" place="8" resultid="14949" />
                    <RANKING order="9" place="9" resultid="17468" />
                    <RANKING order="10" place="10" resultid="14972" />
                    <RANKING order="11" place="11" resultid="16043" />
                    <RANKING order="12" place="12" resultid="14423" />
                    <RANKING order="13" place="13" resultid="18176" />
                    <RANKING order="14" place="14" resultid="17760" />
                    <RANKING order="15" place="15" resultid="17955" />
                    <RANKING order="16" place="16" resultid="16690" />
                    <RANKING order="17" place="17" resultid="14264" />
                    <RANKING order="18" place="18" resultid="16589" />
                    <RANKING order="19" place="19" resultid="17924" />
                    <RANKING order="20" place="-1" resultid="17399" />
                    <RANKING order="21" place="-1" resultid="17405" />
                    <RANKING order="22" place="-1" resultid="17779" />
                    <RANKING order="23" place="-1" resultid="17864" />
                    <RANKING order="24" place="-1" resultid="14638" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14249" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14967" />
                    <RANKING order="2" place="2" resultid="18449" />
                    <RANKING order="3" place="3" resultid="14737" />
                    <RANKING order="4" place="4" resultid="17672" />
                    <RANKING order="5" place="5" resultid="16034" />
                    <RANKING order="6" place="6" resultid="17651" />
                    <RANKING order="7" place="7" resultid="14708" />
                    <RANKING order="8" place="8" resultid="17995" />
                    <RANKING order="9" place="-1" resultid="14898" />
                    <RANKING order="10" place="-1" resultid="16085" />
                    <RANKING order="11" place="-1" resultid="16138" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14250" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17340" />
                    <RANKING order="2" place="2" resultid="14299" />
                    <RANKING order="3" place="3" resultid="18458" />
                    <RANKING order="4" place="4" resultid="18509" />
                    <RANKING order="5" place="5" resultid="14910" />
                    <RANKING order="6" place="6" resultid="15010" />
                    <RANKING order="7" place="7" resultid="16127" />
                    <RANKING order="8" place="8" resultid="18549" />
                    <RANKING order="9" place="9" resultid="15194" />
                    <RANKING order="10" place="10" resultid="16945" />
                    <RANKING order="11" place="-1" resultid="18537" />
                    <RANKING order="12" place="-1" resultid="14619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14251" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14924" />
                    <RANKING order="2" place="2" resultid="16364" />
                    <RANKING order="3" place="3" resultid="15785" />
                    <RANKING order="4" place="4" resultid="18118" />
                    <RANKING order="5" place="5" resultid="16324" />
                    <RANKING order="6" place="-1" resultid="17319" />
                    <RANKING order="7" place="-1" resultid="18284" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14252" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15399" />
                    <RANKING order="2" place="2" resultid="14750" />
                    <RANKING order="3" place="3" resultid="17749" />
                    <RANKING order="4" place="4" resultid="15938" />
                    <RANKING order="5" place="5" resultid="18636" />
                    <RANKING order="6" place="6" resultid="16247" />
                    <RANKING order="7" place="-1" resultid="16702" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14253" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17451" />
                    <RANKING order="2" place="2" resultid="17110" />
                    <RANKING order="3" place="3" resultid="14523" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14254" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14360" />
                    <RANKING order="2" place="2" resultid="16333" />
                    <RANKING order="3" place="3" resultid="14414" />
                    <RANKING order="4" place="-1" resultid="16414" />
                    <RANKING order="5" place="-1" resultid="16455" />
                    <RANKING order="6" place="-1" resultid="17286" />
                    <RANKING order="7" place="-1" resultid="17741" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14255" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14560" />
                    <RANKING order="2" place="2" resultid="14454" />
                    <RANKING order="3" place="3" resultid="15810" />
                    <RANKING order="4" place="4" resultid="14929" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14256" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17346" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14257" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="14258" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="14259" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19397" daytime="11:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19398" daytime="11:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19399" daytime="11:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19400" daytime="12:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19401" daytime="12:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19402" daytime="12:05" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19403" daytime="12:05" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19404" daytime="12:05" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="19405" daytime="12:10" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="19406" daytime="12:10" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="19407" daytime="12:15" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="19408" daytime="12:15" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="19409" daytime="12:20" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="19410" daytime="12:20" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1256" daytime="10:30" gender="F" number="14" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1257" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16580" />
                    <RANKING order="2" place="2" resultid="15730" />
                    <RANKING order="3" place="3" resultid="14613" />
                    <RANKING order="4" place="4" resultid="16540" />
                    <RANKING order="5" place="5" resultid="16603" />
                    <RANKING order="6" place="-1" resultid="16637" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1258" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14836" />
                    <RANKING order="2" place="2" resultid="17592" />
                    <RANKING order="3" place="3" resultid="16749" />
                    <RANKING order="4" place="4" resultid="15232" />
                    <RANKING order="5" place="5" resultid="17378" />
                    <RANKING order="6" place="6" resultid="14571" />
                    <RANKING order="7" place="-1" resultid="14647" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1259" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16599" />
                    <RANKING order="2" place="2" resultid="18354" />
                    <RANKING order="3" place="3" resultid="16918" />
                    <RANKING order="4" place="4" resultid="18425" />
                    <RANKING order="5" place="5" resultid="14757" />
                    <RANKING order="6" place="-1" resultid="18396" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1260" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14590" />
                    <RANKING order="2" place="2" resultid="15853" />
                    <RANKING order="3" place="3" resultid="16831" />
                    <RANKING order="4" place="4" resultid="18134" />
                    <RANKING order="5" place="5" resultid="15866" />
                    <RANKING order="6" place="6" resultid="17497" />
                    <RANKING order="7" place="7" resultid="16167" />
                    <RANKING order="8" place="8" resultid="15413" />
                    <RANKING order="9" place="-1" resultid="15418" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1261" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16015" />
                    <RANKING order="2" place="2" resultid="15347" />
                    <RANKING order="3" place="3" resultid="17772" />
                    <RANKING order="4" place="4" resultid="17802" />
                    <RANKING order="5" place="5" resultid="15359" />
                    <RANKING order="6" place="6" resultid="14892" />
                    <RANKING order="7" place="7" resultid="18146" />
                    <RANKING order="8" place="-1" resultid="15423" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1262" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16461" />
                    <RANKING order="2" place="2" resultid="15200" />
                    <RANKING order="3" place="3" resultid="17558" />
                    <RANKING order="4" place="4" resultid="15842" />
                    <RANKING order="5" place="5" resultid="16372" />
                    <RANKING order="6" place="6" resultid="16380" />
                    <RANKING order="7" place="7" resultid="14809" />
                    <RANKING order="8" place="8" resultid="16289" />
                    <RANKING order="9" place="9" resultid="15946" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1263" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15796" />
                    <RANKING order="2" place="2" resultid="18106" />
                    <RANKING order="3" place="3" resultid="17205" />
                    <RANKING order="4" place="4" resultid="16533" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1264" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16467" />
                    <RANKING order="2" place="2" resultid="15243" />
                    <RANKING order="3" place="3" resultid="14488" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1265" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16389" />
                    <RANKING order="2" place="2" resultid="17191" />
                    <RANKING order="3" place="3" resultid="17093" />
                    <RANKING order="4" place="4" resultid="14846" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1266" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15206" />
                    <RANKING order="2" place="2" resultid="17726" />
                    <RANKING order="3" place="3" resultid="14493" />
                    <RANKING order="4" place="4" resultid="17436" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1267" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14459" />
                    <RANKING order="2" place="2" resultid="16341" />
                    <RANKING order="3" place="3" resultid="14405" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1268" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1269" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1270" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18312" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1271" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1272" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19366" daytime="10:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19367" daytime="10:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19368" daytime="10:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19369" daytime="10:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19370" daytime="10:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19371" daytime="10:45" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19372" daytime="10:45" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1358" daytime="13:00" gender="F" number="20" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="16646" agemax="99" agemin="80" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="16638" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16647" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18014" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16648" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17871" />
                    <RANKING order="2" place="2" resultid="17516" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16649" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18228" />
                    <RANKING order="2" place="2" resultid="15967" />
                    <RANKING order="3" place="3" resultid="15368" />
                    <RANKING order="4" place="4" resultid="16303" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16650" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15306" />
                    <RANKING order="2" place="2" resultid="16482" />
                    <RANKING order="3" place="-1" resultid="14901" />
                    <RANKING order="4" place="-1" resultid="17241" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16651" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16483" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16652" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14534" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19419" daytime="13:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19420" daytime="13:05" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1205" daytime="09:10" gender="M" number="11" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1206" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15048" />
                    <RANKING order="2" place="2" resultid="18606" />
                    <RANKING order="3" place="3" resultid="18338" />
                    <RANKING order="4" place="4" resultid="16706" />
                    <RANKING order="5" place="5" resultid="17830" />
                    <RANKING order="6" place="6" resultid="17839" />
                    <RANKING order="7" place="7" resultid="16718" />
                    <RANKING order="8" place="-1" resultid="14772" />
                    <RANKING order="9" place="-1" resultid="15016" />
                    <RANKING order="10" place="-1" resultid="18568" />
                    <RANKING order="11" place="-1" resultid="18614" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1207" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16930" />
                    <RANKING order="2" place="2" resultid="16712" />
                    <RANKING order="3" place="3" resultid="16924" />
                    <RANKING order="4" place="4" resultid="16742" />
                    <RANKING order="5" place="5" resultid="14602" />
                    <RANKING order="6" place="-1" resultid="17294" />
                    <RANKING order="7" place="-1" resultid="18166" />
                    <RANKING order="8" place="-1" resultid="15382" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1208" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16684" />
                    <RANKING order="2" place="2" resultid="16880" />
                    <RANKING order="3" place="3" resultid="18586" />
                    <RANKING order="4" place="4" resultid="18388" />
                    <RANKING order="5" place="5" resultid="17441" />
                    <RANKING order="6" place="6" resultid="18476" />
                    <RANKING order="7" place="7" resultid="16865" />
                    <RANKING order="8" place="8" resultid="17354" />
                    <RANKING order="9" place="9" resultid="14503" />
                    <RANKING order="10" place="10" resultid="17936" />
                    <RANKING order="11" place="-1" resultid="18154" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1209" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18374" />
                    <RANKING order="2" place="2" resultid="17474" />
                    <RANKING order="3" place="3" resultid="17020" />
                    <RANKING order="4" place="4" resultid="17371" />
                    <RANKING order="5" place="5" resultid="17211" />
                    <RANKING order="6" place="6" resultid="15294" />
                    <RANKING order="7" place="7" resultid="17048" />
                    <RANKING order="8" place="8" resultid="18206" />
                    <RANKING order="9" place="9" resultid="17273" />
                    <RANKING order="10" place="10" resultid="17713" />
                    <RANKING order="11" place="11" resultid="16191" />
                    <RANKING order="12" place="12" resultid="16846" />
                    <RANKING order="13" place="13" resultid="17835" />
                    <RANKING order="14" place="14" resultid="16820" />
                    <RANKING order="15" place="15" resultid="16357" />
                    <RANKING order="16" place="-1" resultid="14816" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1210" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17008" />
                    <RANKING order="2" place="2" resultid="18528" />
                    <RANKING order="3" place="3" resultid="14422" />
                    <RANKING order="4" place="4" resultid="17467" />
                    <RANKING order="5" place="5" resultid="17759" />
                    <RANKING order="6" place="6" resultid="18175" />
                    <RANKING order="7" place="7" resultid="14936" />
                    <RANKING order="8" place="8" resultid="17793" />
                    <RANKING order="9" place="9" resultid="16838" />
                    <RANKING order="10" place="10" resultid="16689" />
                    <RANKING order="11" place="11" resultid="16934" />
                    <RANKING order="12" place="12" resultid="18192" />
                    <RANKING order="13" place="-1" resultid="17970" />
                    <RANKING order="14" place="-1" resultid="14637" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1211" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14736" />
                    <RANKING order="2" place="2" resultid="18448" />
                    <RANKING order="3" place="3" resultid="16438" />
                    <RANKING order="4" place="4" resultid="16080" />
                    <RANKING order="5" place="5" resultid="16137" />
                    <RANKING order="6" place="6" resultid="17650" />
                    <RANKING order="7" place="7" resultid="17564" />
                    <RANKING order="8" place="-1" resultid="18006" />
                    <RANKING order="9" place="-1" resultid="16984" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1212" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17339" />
                    <RANKING order="2" place="2" resultid="18508" />
                    <RANKING order="3" place="3" resultid="14298" />
                    <RANKING order="4" place="4" resultid="17222" />
                    <RANKING order="5" place="5" resultid="15009" />
                    <RANKING order="6" place="6" resultid="18276" />
                    <RANKING order="7" place="7" resultid="16431" />
                    <RANKING order="8" place="-1" resultid="15006" />
                    <RANKING order="9" place="-1" resultid="16990" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1213" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15742" />
                    <RANKING order="2" place="2" resultid="18214" />
                    <RANKING order="3" place="3" resultid="16363" />
                    <RANKING order="4" place="4" resultid="14598" />
                    <RANKING order="5" place="5" resultid="16229" />
                    <RANKING order="6" place="6" resultid="14513" />
                    <RANKING order="7" place="7" resultid="17310" />
                    <RANKING order="8" place="-1" resultid="15773" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1214" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17573" />
                    <RANKING order="2" place="2" resultid="15247" />
                    <RANKING order="3" place="3" resultid="14396" />
                    <RANKING order="4" place="4" resultid="14439" />
                    <RANKING order="5" place="5" resultid="17748" />
                    <RANKING order="6" place="6" resultid="18963" />
                    <RANKING order="7" place="7" resultid="16701" />
                    <RANKING order="8" place="8" resultid="16183" />
                    <RANKING order="9" place="9" resultid="15937" />
                    <RANKING order="10" place="10" resultid="16246" />
                    <RANKING order="11" place="11" resultid="16253" />
                    <RANKING order="12" place="12" resultid="16422" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1215" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18267" />
                    <RANKING order="2" place="2" resultid="17734" />
                    <RANKING order="3" place="3" resultid="15216" />
                    <RANKING order="4" place="4" resultid="18521" />
                    <RANKING order="5" place="5" resultid="15287" />
                    <RANKING order="6" place="6" resultid="14853" />
                    <RANKING order="7" place="7" resultid="15802" />
                    <RANKING order="8" place="8" resultid="17054" />
                    <RANKING order="9" place="9" resultid="16385" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1216" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14497" />
                    <RANKING order="2" place="2" resultid="17073" />
                    <RANKING order="3" place="3" resultid="16449" />
                    <RANKING order="4" place="-1" resultid="16454" />
                    <RANKING order="5" place="-1" resultid="17285" />
                    <RANKING order="6" place="-1" resultid="17740" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1217" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15809" />
                    <RANKING order="2" place="2" resultid="14380" />
                    <RANKING order="3" place="3" resultid="17062" />
                    <RANKING order="4" place="4" resultid="14387" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1218" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15763" />
                    <RANKING order="2" place="2" resultid="18298" />
                    <RANKING order="3" place="3" resultid="17345" />
                    <RANKING order="4" place="-1" resultid="15816" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1219" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14825" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1220" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1221" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19342" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19343" daytime="09:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19344" daytime="09:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19345" daytime="09:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19346" daytime="09:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19347" daytime="09:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19348" daytime="09:20" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19349" daytime="09:25" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="19350" daytime="09:25" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="19351" daytime="09:25" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="19352" daytime="09:25" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="19353" daytime="09:30" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2017-11-18" daytime="16:00" endtime="20:21" name="BLOK III" number="3" warmupfrom="15:00">
          <EVENTS>
            <EVENT eventid="1440" daytime="17:05" gender="M" number="25" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1441" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15052" />
                    <RANKING order="2" place="2" resultid="18609" />
                    <RANKING order="3" place="3" resultid="16623" />
                    <RANKING order="4" place="4" resultid="18616" />
                    <RANKING order="5" place="5" resultid="14767" />
                    <RANKING order="6" place="6" resultid="16708" />
                    <RANKING order="7" place="7" resultid="18341" />
                    <RANKING order="8" place="8" resultid="14774" />
                    <RANKING order="9" place="9" resultid="17990" />
                    <RANKING order="10" place="10" resultid="16720" />
                    <RANKING order="11" place="11" resultid="17029" />
                    <RANKING order="12" place="-1" resultid="18061" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1442" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16714" />
                    <RANKING order="2" place="2" resultid="16926" />
                    <RANKING order="3" place="3" resultid="17488" />
                    <RANKING order="4" place="4" resultid="16951" />
                    <RANKING order="5" place="5" resultid="16744" />
                    <RANKING order="6" place="6" resultid="17296" />
                    <RANKING order="7" place="7" resultid="16223" />
                    <RANKING order="8" place="8" resultid="18349" />
                    <RANKING order="9" place="9" resultid="14674" />
                    <RANKING order="10" place="10" resultid="16834" />
                    <RANKING order="11" place="11" resultid="17978" />
                    <RANKING order="12" place="12" resultid="16758" />
                    <RANKING order="13" place="13" resultid="16278" />
                    <RANKING order="14" place="14" resultid="16143" />
                    <RANKING order="15" place="-1" resultid="14609" />
                    <RANKING order="16" place="-1" resultid="15976" />
                    <RANKING order="17" place="-1" resultid="18495" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1443" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14449" />
                    <RANKING order="2" place="2" resultid="15276" />
                    <RANKING order="3" place="3" resultid="18390" />
                    <RANKING order="4" place="4" resultid="18477" />
                    <RANKING order="5" place="5" resultid="18588" />
                    <RANKING order="6" place="6" resultid="17918" />
                    <RANKING order="7" place="7" resultid="15046" />
                    <RANKING order="8" place="8" resultid="16867" />
                    <RANKING order="9" place="8" resultid="17442" />
                    <RANKING order="10" place="10" resultid="18383" />
                    <RANKING order="11" place="11" resultid="17912" />
                    <RANKING order="12" place="12" resultid="17356" />
                    <RANKING order="13" place="13" resultid="17081" />
                    <RANKING order="14" place="14" resultid="18156" />
                    <RANKING order="15" place="-1" resultid="14505" />
                    <RANKING order="16" place="-1" resultid="15446" />
                    <RANKING order="17" place="-1" resultid="15900" />
                    <RANKING order="18" place="-1" resultid="17698" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1444" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18376" />
                    <RANKING order="2" place="2" resultid="17476" />
                    <RANKING order="3" place="3" resultid="17693" />
                    <RANKING order="4" place="4" resultid="16204" />
                    <RANKING order="5" place="5" resultid="17022" />
                    <RANKING order="6" place="6" resultid="17200" />
                    <RANKING order="7" place="7" resultid="16826" />
                    <RANKING order="8" place="8" resultid="15297" />
                    <RANKING order="9" place="9" resultid="16800" />
                    <RANKING order="10" place="10" resultid="16806" />
                    <RANKING order="11" place="11" resultid="17581" />
                    <RANKING order="12" place="12" resultid="16193" />
                    <RANKING order="13" place="13" resultid="16811" />
                    <RANKING order="14" place="14" resultid="17043" />
                    <RANKING order="15" place="15" resultid="16848" />
                    <RANKING order="16" place="16" resultid="18466" />
                    <RANKING order="17" place="17" resultid="16765" />
                    <RANKING order="18" place="-1" resultid="15908" />
                    <RANKING order="19" place="-1" resultid="16853" />
                    <RANKING order="20" place="-1" resultid="17136" />
                    <RANKING order="21" place="-1" resultid="17458" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1445" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18558" />
                    <RANKING order="2" place="2" resultid="17010" />
                    <RANKING order="3" place="3" resultid="15059" />
                    <RANKING order="4" place="4" resultid="17469" />
                    <RANKING order="5" place="5" resultid="16045" />
                    <RANKING order="6" place="6" resultid="14424" />
                    <RANKING order="7" place="7" resultid="16771" />
                    <RANKING order="8" place="8" resultid="17795" />
                    <RANKING order="9" place="9" resultid="14950" />
                    <RANKING order="10" place="10" resultid="16840" />
                    <RANKING order="11" place="11" resultid="17956" />
                    <RANKING order="12" place="12" resultid="17865" />
                    <RANKING order="13" place="13" resultid="18177" />
                    <RANKING order="14" place="14" resultid="14265" />
                    <RANKING order="15" place="15" resultid="16590" />
                    <RANKING order="16" place="16" resultid="18194" />
                    <RANKING order="17" place="-1" resultid="17005" />
                    <RANKING order="18" place="-1" resultid="17400" />
                    <RANKING order="19" place="-1" resultid="17925" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1446" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18415" />
                    <RANKING order="2" place="2" resultid="17611" />
                    <RANKING order="3" place="3" resultid="17616" />
                    <RANKING order="4" place="4" resultid="18450" />
                    <RANKING order="5" place="5" resultid="14969" />
                    <RANKING order="6" place="6" resultid="16439" />
                    <RANKING order="7" place="7" resultid="17673" />
                    <RANKING order="8" place="8" resultid="15040" />
                    <RANKING order="9" place="9" resultid="16076" />
                    <RANKING order="10" place="10" resultid="16036" />
                    <RANKING order="11" place="11" resultid="17625" />
                    <RANKING order="12" place="12" resultid="14899" />
                    <RANKING order="13" place="13" resultid="17566" />
                    <RANKING order="14" place="14" resultid="16086" />
                    <RANKING order="15" place="15" resultid="16095" />
                    <RANKING order="16" place="-1" resultid="16139" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1447" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14300" />
                    <RANKING order="2" place="2" resultid="18538" />
                    <RANKING order="3" place="3" resultid="18510" />
                    <RANKING order="4" place="4" resultid="14911" />
                    <RANKING order="5" place="5" resultid="17681" />
                    <RANKING order="6" place="6" resultid="15011" />
                    <RANKING order="7" place="7" resultid="18294" />
                    <RANKING order="8" place="8" resultid="17148" />
                    <RANKING order="9" place="9" resultid="16477" />
                    <RANKING order="10" place="10" resultid="15195" />
                    <RANKING order="11" place="-1" resultid="16992" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1448" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15744" />
                    <RANKING order="2" place="2" resultid="17216" />
                    <RANKING order="3" place="3" resultid="16365" />
                    <RANKING order="4" place="4" resultid="18320" />
                    <RANKING order="5" place="5" resultid="14515" />
                    <RANKING order="6" place="6" resultid="14351" />
                    <RANKING order="7" place="7" resultid="15920" />
                    <RANKING order="8" place="8" resultid="14979" />
                    <RANKING order="9" place="9" resultid="17312" />
                    <RANKING order="10" place="10" resultid="16326" />
                    <RANKING order="11" place="-1" resultid="15363" />
                    <RANKING order="12" place="-1" resultid="17320" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1449" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17574" />
                    <RANKING order="2" place="2" resultid="15249" />
                    <RANKING order="3" place="3" resultid="14275" />
                    <RANKING order="4" place="4" resultid="15939" />
                    <RANKING order="5" place="5" resultid="16256" />
                    <RANKING order="6" place="-1" resultid="18637" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1450" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18269" />
                    <RANKING order="2" place="2" resultid="14702" />
                    <RANKING order="3" place="3" resultid="17111" />
                    <RANKING order="4" place="4" resultid="14524" />
                    <RANKING order="5" place="5" resultid="15804" />
                    <RANKING order="6" place="6" resultid="14464" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1451" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14566" />
                    <RANKING order="2" place="2" resultid="14361" />
                    <RANKING order="3" place="3" resultid="15266" />
                    <RANKING order="4" place="4" resultid="16456" />
                    <RANKING order="5" place="-1" resultid="14498" />
                    <RANKING order="6" place="-1" resultid="17287" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1452" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14561" />
                    <RANKING order="2" place="2" resultid="14292" />
                    <RANKING order="3" place="3" resultid="16179" />
                    <RANKING order="4" place="4" resultid="15812" />
                    <RANKING order="5" place="5" resultid="14382" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1453" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17348" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1454" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1455" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1456" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19450" daytime="17:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19451" daytime="17:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19452" daytime="17:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19453" daytime="17:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19454" daytime="17:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19455" daytime="17:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19456" daytime="17:15" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19457" daytime="17:15" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="19458" daytime="17:20" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="19459" daytime="17:20" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="19460" daytime="17:20" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="19461" daytime="17:20" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="19462" daytime="17:25" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="19463" daytime="17:25" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="19464" daytime="17:25" number="15" order="15" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1474" daytime="17:40" gender="M" number="27" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1475" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18610" />
                    <RANKING order="2" place="2" resultid="18342" />
                    <RANKING order="3" place="3" resultid="17832" />
                    <RANKING order="4" place="4" resultid="18617" />
                    <RANKING order="5" place="5" resultid="15019" />
                    <RANKING order="6" place="6" resultid="17841" />
                    <RANKING order="7" place="7" resultid="18957" />
                    <RANKING order="8" place="-1" resultid="18571" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1476" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16745" />
                    <RANKING order="2" place="2" resultid="17297" />
                    <RANKING order="3" place="3" resultid="15892" />
                    <RANKING order="4" place="4" resultid="14604" />
                    <RANKING order="5" place="-1" resultid="15384" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1477" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16882" />
                    <RANKING order="2" place="2" resultid="18391" />
                    <RANKING order="3" place="3" resultid="17919" />
                    <RANKING order="4" place="4" resultid="18589" />
                    <RANKING order="5" place="5" resultid="14506" />
                    <RANKING order="6" place="6" resultid="17938" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1478" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18377" />
                    <RANKING order="2" place="2" resultid="17212" />
                    <RANKING order="3" place="3" resultid="17023" />
                    <RANKING order="4" place="4" resultid="17050" />
                    <RANKING order="5" place="5" resultid="17230" />
                    <RANKING order="6" place="6" resultid="17275" />
                    <RANKING order="7" place="7" resultid="17716" />
                    <RANKING order="8" place="8" resultid="17836" />
                    <RANKING order="9" place="9" resultid="16359" />
                    <RANKING order="10" place="10" resultid="15033" />
                    <RANKING order="11" place="-1" resultid="14819" />
                    <RANKING order="12" place="-1" resultid="16173" />
                    <RANKING order="13" place="-1" resultid="16821" />
                    <RANKING order="14" place="-1" resultid="17477" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1479" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17011" />
                    <RANKING order="2" place="2" resultid="18530" />
                    <RANKING order="3" place="3" resultid="14639" />
                    <RANKING order="4" place="4" resultid="14425" />
                    <RANKING order="5" place="5" resultid="17761" />
                    <RANKING order="6" place="6" resultid="14973" />
                    <RANKING order="7" place="7" resultid="18178" />
                    <RANKING order="8" place="8" resultid="16691" />
                    <RANKING order="9" place="9" resultid="16936" />
                    <RANKING order="10" place="-1" resultid="14937" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1480" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14738" />
                    <RANKING order="2" place="2" resultid="18451" />
                    <RANKING order="3" place="3" resultid="14696" />
                    <RANKING order="4" place="4" resultid="16140" />
                    <RANKING order="5" place="5" resultid="17652" />
                    <RANKING order="6" place="6" resultid="18009" />
                    <RANKING order="7" place="-1" resultid="16986" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1481" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17341" />
                    <RANKING order="2" place="2" resultid="17223" />
                    <RANKING order="3" place="3" resultid="15926" />
                    <RANKING order="4" place="4" resultid="14912" />
                    <RANKING order="5" place="5" resultid="18278" />
                    <RANKING order="6" place="6" resultid="16129" />
                    <RANKING order="7" place="-1" resultid="16433" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1482" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15745" />
                    <RANKING order="2" place="2" resultid="16366" />
                    <RANKING order="3" place="3" resultid="15787" />
                    <RANKING order="4" place="4" resultid="14599" />
                    <RANKING order="5" place="5" resultid="14516" />
                    <RANKING order="6" place="6" resultid="14980" />
                    <RANKING order="7" place="-1" resultid="15775" />
                    <RANKING order="8" place="-1" resultid="16231" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1483" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17412" />
                    <RANKING order="2" place="2" resultid="15401" />
                    <RANKING order="3" place="3" resultid="17750" />
                    <RANKING order="4" place="4" resultid="14398" />
                    <RANKING order="5" place="5" resultid="14441" />
                    <RANKING order="6" place="6" resultid="18965" />
                    <RANKING order="7" place="7" resultid="16185" />
                    <RANKING order="8" place="8" resultid="16248" />
                    <RANKING order="9" place="-1" resultid="18440" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1484" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18270" />
                    <RANKING order="2" place="2" resultid="15219" />
                    <RANKING order="3" place="3" resultid="17735" />
                    <RANKING order="4" place="4" resultid="14659" />
                    <RANKING order="5" place="5" resultid="17056" />
                    <RANKING order="6" place="-1" resultid="14855" />
                    <RANKING order="7" place="-1" resultid="15289" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1485" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14499" />
                    <RANKING order="2" place="2" resultid="16450" />
                    <RANKING order="3" place="3" resultid="17076" />
                    <RANKING order="4" place="-1" resultid="17742" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1486" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17064" />
                    <RANKING order="2" place="2" resultid="14389" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1487" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18301" />
                    <RANKING order="2" place="2" resultid="15765" />
                    <RANKING order="3" place="-1" resultid="15818" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1488" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1489" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1490" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19470" daytime="17:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19471" daytime="17:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19472" daytime="17:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19473" daytime="17:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19474" daytime="17:55" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19475" daytime="17:55" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19476" daytime="18:00" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19477" daytime="18:00" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="19478" daytime="18:05" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1548" daytime="19:35" gender="M" number="31" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="16667" agemax="99" agemin="80" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="17877" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16668" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16773" />
                    <RANKING order="2" place="2" resultid="16641" />
                    <RANKING order="3" place="3" resultid="18020" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16669" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18401" />
                    <RANKING order="2" place="2" resultid="17517" />
                    <RANKING order="3" place="3" resultid="17245" />
                    <RANKING order="4" place="4" resultid="16891" />
                    <RANKING order="5" place="5" resultid="17119" />
                    <RANKING order="6" place="6" resultid="18017" />
                    <RANKING order="7" place="7" resultid="14955" />
                    <RANKING order="8" place="8" resultid="17518" />
                    <RANKING order="9" place="9" resultid="16892" />
                    <RANKING order="10" place="10" resultid="16893" />
                    <RANKING order="11" place="-1" resultid="16775" />
                    <RANKING order="12" place="-1" resultid="17719" />
                    <RANKING order="13" place="-1" resultid="18231" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16670" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17655" />
                    <RANKING order="2" place="2" resultid="16089" />
                    <RANKING order="3" place="3" resultid="17876" />
                    <RANKING order="4" place="4" resultid="16090" />
                    <RANKING order="5" place="5" resultid="18019" />
                    <RANKING order="6" place="-1" resultid="14904" />
                    <RANKING order="7" place="-1" resultid="15369" />
                    <RANKING order="8" place="-1" resultid="15996" />
                    <RANKING order="9" place="-1" resultid="18233" />
                    <RANKING order="10" place="-1" resultid="18541" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16671" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18322" />
                    <RANKING order="2" place="2" resultid="17246" />
                    <RANKING order="3" place="3" resultid="18235" />
                    <RANKING order="4" place="4" resultid="15307" />
                    <RANKING order="5" place="5" resultid="15970" />
                    <RANKING order="6" place="-1" resultid="16209" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16672" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16489" />
                    <RANKING order="2" place="2" resultid="15309" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16673" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14537" />
                    <RANKING order="2" place="2" resultid="17116" />
                    <RANKING order="3" place="3" resultid="16490" />
                    <RANKING order="4" place="-1" resultid="15831" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19499" daytime="19:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19500" daytime="19:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19501" daytime="19:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19502" daytime="19:45" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="16953" daytime="16:00" gender="M" number="43" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="16955" agemax="99" agemin="80" calculate="TOTAL" />
                <AGEGROUP agegroupid="16956" agemax="119" agemin="100" calculate="TOTAL" />
                <AGEGROUP agegroupid="16957" agemax="159" agemin="120" calculate="TOTAL" />
                <AGEGROUP agegroupid="16958" agemax="199" agemin="160" calculate="TOTAL" />
                <AGEGROUP agegroupid="16959" agemax="239" agemin="200" calculate="TOTAL" />
                <AGEGROUP agegroupid="16960" agemax="279" agemin="240" calculate="TOTAL" />
                <AGEGROUP agegroupid="16961" agemax="-1" agemin="280" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19425" daytime="16:00" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1578" daytime="20:15" gender="M" number="33" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1579" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17325" />
                    <RANKING order="2" place="2" resultid="16216" />
                    <RANKING order="3" place="3" resultid="16271" />
                    <RANKING order="4" place="4" resultid="16263" />
                    <RANKING order="5" place="-1" resultid="17991" />
                    <RANKING order="6" place="-1" resultid="18055" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1580" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18168" />
                    <RANKING order="2" place="2" resultid="16696" />
                    <RANKING order="3" place="3" resultid="18503" />
                    <RANKING order="4" place="4" resultid="15893" />
                    <RANKING order="5" place="5" resultid="15438" />
                    <RANKING order="6" place="6" resultid="18350" />
                    <RANKING order="7" place="-1" resultid="15392" />
                    <RANKING order="8" place="-1" resultid="15977" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1581" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15901" />
                    <RANKING order="2" place="2" resultid="16546" />
                    <RANKING order="3" place="3" resultid="15447" />
                    <RANKING order="4" place="4" resultid="18128" />
                    <RANKING order="5" place="-1" resultid="16883" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1582" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17174" />
                    <RANKING order="2" place="2" resultid="18209" />
                    <RANKING order="3" place="3" resultid="17582" />
                    <RANKING order="4" place="4" resultid="17276" />
                    <RANKING order="5" place="5" resultid="15909" />
                    <RANKING order="6" place="-1" resultid="16860" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1583" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18186" />
                    <RANKING order="2" place="2" resultid="16529" />
                    <RANKING order="3" place="3" resultid="14640" />
                    <RANKING order="4" place="4" resultid="17796" />
                    <RANKING order="5" place="5" resultid="17762" />
                    <RANKING order="6" place="6" resultid="16054" />
                    <RANKING order="7" place="-1" resultid="14426" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1584" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16070" />
                    <RANKING order="2" place="2" resultid="14697" />
                    <RANKING order="3" place="3" resultid="18223" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1585" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15927" />
                    <RANKING order="2" place="2" resultid="18539" />
                    <RANKING order="3" place="3" resultid="15861" />
                    <RANKING order="4" place="4" resultid="16434" />
                    <RANKING order="5" place="-1" resultid="18460" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1586" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18217" />
                    <RANKING order="2" place="2" resultid="14352" />
                    <RANKING order="3" place="3" resultid="18120" />
                    <RANKING order="4" place="4" resultid="16232" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1587" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14731" />
                    <RANKING order="2" place="2" resultid="17751" />
                    <RANKING order="3" place="3" resultid="18966" />
                    <RANKING order="4" place="4" resultid="15259" />
                    <RANKING order="5" place="-1" resultid="14399" />
                    <RANKING order="6" place="-1" resultid="14668" />
                    <RANKING order="7" place="-1" resultid="15250" />
                    <RANKING order="8" place="-1" resultid="16249" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1588" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17453" />
                    <RANKING order="2" place="2" resultid="15827" />
                    <RANKING order="3" place="3" resultid="14660" />
                    <RANKING order="4" place="4" resultid="17057" />
                    <RANKING order="5" place="-1" resultid="17143" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1589" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14362" />
                    <RANKING order="2" place="2" resultid="16335" />
                    <RANKING order="3" place="-1" resultid="14416" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1590" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14383" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1591" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1592" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1593" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1594" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19506" daytime="20:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19507" daytime="20:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19508" daytime="20:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19509" daytime="20:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19510" daytime="20:55" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19511" daytime="21:00" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19512" daytime="21:10" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1555" daytime="19:50" gender="F" number="32" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1562" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17237" />
                    <RANKING order="2" place="2" resultid="17945" />
                    <RANKING order="3" place="3" resultid="18163" />
                    <RANKING order="4" place="4" resultid="14795" />
                    <RANKING order="5" place="-1" resultid="18604" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1563" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14839" />
                    <RANKING order="2" place="-1" resultid="14650" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1564" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17036" />
                    <RANKING order="2" place="2" resultid="18365" />
                    <RANKING order="3" place="3" resultid="17789" />
                    <RANKING order="4" place="4" resultid="17965" />
                    <RANKING order="5" place="-1" resultid="18485" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1565" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14593" />
                    <RANKING order="2" place="2" resultid="16063" />
                    <RANKING order="3" place="3" resultid="15869" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1566" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="1567" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14529" />
                    <RANKING order="2" place="2" resultid="16374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1568" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16402" />
                    <RANKING order="2" place="2" resultid="18108" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1569" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18625" />
                    <RANKING order="2" place="2" resultid="16470" />
                    <RANKING order="3" place="3" resultid="17817" />
                    <RANKING order="4" place="4" resultid="18433" />
                    <RANKING order="5" place="5" resultid="16161" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1570" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16392" />
                    <RANKING order="2" place="2" resultid="14374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1571" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1572" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1573" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1574" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1575" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1576" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1577" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19503" daytime="19:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19504" daytime="20:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19505" daytime="20:10" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1423" daytime="16:55" gender="F" number="24" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1424" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16582" />
                    <RANKING order="2" place="2" resultid="16609" />
                    <RANKING order="3" place="3" resultid="17944" />
                    <RANKING order="4" place="4" resultid="18162" />
                    <RANKING order="5" place="5" resultid="18202" />
                    <RANKING order="6" place="6" resultid="14614" />
                    <RANKING order="7" place="-1" resultid="17905" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1425" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16752" />
                    <RANKING order="2" place="2" resultid="15736" />
                    <RANKING order="3" place="3" resultid="17856" />
                    <RANKING order="4" place="4" resultid="17509" />
                    <RANKING order="5" place="5" resultid="14573" />
                    <RANKING order="6" place="-1" resultid="15233" />
                    <RANKING order="7" place="-1" resultid="17379" />
                    <RANKING order="8" place="-1" resultid="18098" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1426" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17363" />
                    <RANKING order="2" place="2" resultid="17964" />
                    <RANKING order="3" place="3" resultid="17383" />
                    <RANKING order="4" place="4" resultid="15430" />
                    <RANKING order="5" place="5" resultid="16919" />
                    <RANKING order="6" place="-1" resultid="17482" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1427" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14592" />
                    <RANKING order="2" place="2" resultid="17446" />
                    <RANKING order="3" place="3" resultid="14717" />
                    <RANKING order="4" place="4" resultid="17016" />
                    <RANKING order="5" place="5" resultid="16794" />
                    <RANKING order="6" place="6" resultid="18135" />
                    <RANKING order="7" place="7" resultid="15956" />
                    <RANKING order="8" place="8" resultid="15952" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1428" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16017" />
                    <RANKING order="2" place="2" resultid="15349" />
                    <RANKING order="3" place="-1" resultid="17635" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1429" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16462" />
                    <RANKING order="2" place="2" resultid="15239" />
                    <RANKING order="3" place="3" resultid="16373" />
                    <RANKING order="4" place="4" resultid="15201" />
                    <RANKING order="5" place="5" resultid="17560" />
                    <RANKING order="6" place="6" resultid="16382" />
                    <RANKING order="7" place="7" resultid="15932" />
                    <RANKING order="8" place="8" resultid="14802" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1430" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16312" />
                    <RANKING order="2" place="2" resultid="17599" />
                    <RANKING order="3" place="3" resultid="15069" />
                    <RANKING order="4" place="4" resultid="16535" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1431" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15226" />
                    <RANKING order="2" place="2" resultid="16469" />
                    <RANKING order="3" place="3" resultid="14690" />
                    <RANKING order="4" place="4" resultid="17553" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1432" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14626" />
                    <RANKING order="2" place="2" resultid="16391" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1433" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17727" />
                    <RANKING order="2" place="2" resultid="16408" />
                    <RANKING order="3" place="3" resultid="17642" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1434" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14460" />
                    <RANKING order="2" place="-1" resultid="16344" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1435" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1436" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1437" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1438" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1439" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19444" daytime="16:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19445" daytime="16:55" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19446" daytime="17:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19447" daytime="17:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19448" daytime="17:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19449" daytime="17:00" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1457" daytime="17:30" gender="F" number="26" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1458" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18602" />
                    <RANKING order="2" place="2" resultid="17906" />
                    <RANKING order="3" place="3" resultid="14985" />
                    <RANKING order="4" place="4" resultid="16967" />
                    <RANKING order="5" place="5" resultid="14615" />
                    <RANKING order="6" place="6" resultid="15848" />
                    <RANKING order="7" place="-1" resultid="15408" />
                    <RANKING order="8" place="-1" resultid="18580" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1459" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15234" />
                    <RANKING order="2" place="2" resultid="15737" />
                    <RANKING order="3" place="3" resultid="14831" />
                    <RANKING order="4" place="4" resultid="17510" />
                    <RANKING order="5" place="-1" resultid="14585" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1460" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15001" />
                    <RANKING order="2" place="2" resultid="14871" />
                    <RANKING order="3" place="-1" resultid="18484" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1461" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17017" />
                    <RANKING order="2" place="2" resultid="17931" />
                    <RANKING order="3" place="3" resultid="15878" />
                    <RANKING order="4" place="-1" resultid="17001" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1462" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14942" />
                    <RANKING order="2" place="2" resultid="15885" />
                    <RANKING order="3" place="3" resultid="16009" />
                    <RANKING order="4" place="4" resultid="17803" />
                    <RANKING order="5" place="5" resultid="18092" />
                    <RANKING order="6" place="6" resultid="16294" />
                    <RANKING order="7" place="7" resultid="18148" />
                    <RANKING order="8" place="-1" resultid="17636" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1463" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15240" />
                    <RANKING order="2" place="2" resultid="15843" />
                    <RANKING order="3" place="3" resultid="17102" />
                    <RANKING order="4" place="4" resultid="14803" />
                    <RANKING order="5" place="-1" resultid="14811" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1464" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16313" />
                    <RANKING order="2" place="2" resultid="17206" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1465" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15227" />
                    <RANKING order="2" place="2" resultid="18624" />
                    <RANKING order="3" place="3" resultid="15781" />
                    <RANKING order="4" place="4" resultid="16352" />
                    <RANKING order="5" place="-1" resultid="16151" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1466" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17630" />
                    <RANKING order="2" place="2" resultid="17095" />
                    <RANKING order="3" place="3" resultid="17192" />
                    <RANKING order="4" place="4" resultid="19745" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1467" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15207" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1468" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14406" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1469" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18290" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1470" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1471" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18313" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1472" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1473" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19465" daytime="17:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19466" daytime="17:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19467" daytime="17:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19468" daytime="17:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19469" daytime="17:40" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1406" daytime="16:25" gender="M" number="23" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1407" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17432" />
                    <RANKING order="2" place="2" resultid="17848" />
                    <RANKING order="3" place="3" resultid="18597" />
                    <RANKING order="4" place="4" resultid="16215" />
                    <RANKING order="5" place="5" resultid="14773" />
                    <RANKING order="6" place="6" resultid="14766" />
                    <RANKING order="7" place="7" resultid="15051" />
                    <RANKING order="8" place="8" resultid="18956" />
                    <RANKING order="9" place="9" resultid="17844" />
                    <RANKING order="10" place="10" resultid="16262" />
                    <RANKING order="11" place="-1" resultid="15018" />
                    <RANKING order="12" place="-1" resultid="18570" />
                    <RANKING order="13" place="-1" resultid="18608" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1408" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17826" />
                    <RANKING order="2" place="2" resultid="14270" />
                    <RANKING order="3" place="3" resultid="16727" />
                    <RANKING order="4" place="4" resultid="18494" />
                    <RANKING order="5" place="5" resultid="15391" />
                    <RANKING order="6" place="6" resultid="14673" />
                    <RANKING order="7" place="7" resultid="15458" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1409" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17086" />
                    <RANKING order="2" place="2" resultid="18371" />
                    <RANKING order="3" place="3" resultid="17305" />
                    <RANKING order="4" place="4" resultid="17911" />
                    <RANKING order="5" place="5" resultid="18127" />
                    <RANKING order="6" place="6" resultid="18003" />
                    <RANKING order="7" place="-1" resultid="16616" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1410" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17416" />
                    <RANKING order="2" place="2" resultid="17186" />
                    <RANKING order="3" place="3" resultid="17199" />
                    <RANKING order="4" place="4" resultid="15296" />
                    <RANKING order="5" place="5" resultid="16805" />
                    <RANKING order="6" place="6" resultid="17373" />
                    <RANKING order="7" place="7" resultid="17809" />
                    <RANKING order="8" place="8" resultid="17715" />
                    <RANKING order="9" place="9" resultid="18465" />
                    <RANKING order="10" place="10" resultid="14555" />
                    <RANKING order="11" place="-1" resultid="14818" />
                    <RANKING order="12" place="-1" resultid="14885" />
                    <RANKING order="13" place="-1" resultid="16859" />
                    <RANKING order="14" place="-1" resultid="16871" />
                    <RANKING order="15" place="-1" resultid="16876" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1411" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18557" />
                    <RANKING order="2" place="2" resultid="17822" />
                    <RANKING order="3" place="3" resultid="17588" />
                    <RANKING order="4" place="4" resultid="16026" />
                    <RANKING order="5" place="5" resultid="18420" />
                    <RANKING order="6" place="6" resultid="16044" />
                    <RANKING order="7" place="7" resultid="17406" />
                    <RANKING order="8" place="8" resultid="16318" />
                    <RANKING order="9" place="9" resultid="14278" />
                    <RANKING order="10" place="10" resultid="17780" />
                    <RANKING order="11" place="11" resultid="17544" />
                    <RANKING order="12" place="12" resultid="14723" />
                    <RANKING order="13" place="-1" resultid="14785" />
                    <RANKING order="14" place="-1" resultid="15453" />
                    <RANKING order="15" place="-1" resultid="17503" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1412" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14968" />
                    <RANKING order="2" place="2" resultid="16069" />
                    <RANKING order="3" place="3" resultid="14864" />
                    <RANKING order="4" place="4" resultid="16035" />
                    <RANKING order="5" place="5" resultid="14709" />
                    <RANKING order="6" place="6" resultid="18140" />
                    <RANKING order="7" place="7" resultid="17367" />
                    <RANKING order="8" place="-1" resultid="18008" />
                    <RANKING order="9" place="-1" resultid="16239" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1413" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16128" />
                    <RANKING order="2" place="2" resultid="18550" />
                    <RANKING order="3" place="3" resultid="16476" />
                    <RANKING order="4" place="4" resultid="15760" />
                    <RANKING order="5" place="5" resultid="15860" />
                    <RANKING order="6" place="6" resultid="17393" />
                    <RANKING order="7" place="7" resultid="16946" />
                    <RANKING order="8" place="-1" resultid="14620" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1414" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18469" />
                    <RANKING order="2" place="2" resultid="18285" />
                    <RANKING order="3" place="3" resultid="17180" />
                    <RANKING order="4" place="4" resultid="15786" />
                    <RANKING order="5" place="5" resultid="18119" />
                    <RANKING order="6" place="6" resultid="15279" />
                    <RANKING order="7" place="7" resultid="15272" />
                    <RANKING order="8" place="8" resultid="16325" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1415" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14730" />
                    <RANKING order="2" place="2" resultid="15400" />
                    <RANKING order="3" place="3" resultid="15822" />
                    <RANKING order="4" place="4" resultid="16255" />
                    <RANKING order="5" place="5" resultid="16424" />
                    <RANKING order="6" place="-1" resultid="18439" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1416" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17452" />
                    <RANKING order="2" place="2" resultid="15218" />
                    <RANKING order="3" place="3" resultid="18523" />
                    <RANKING order="4" place="4" resultid="15288" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1417" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15916" />
                    <RANKING order="2" place="2" resultid="17075" />
                    <RANKING order="3" place="3" resultid="14415" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1418" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14475" />
                    <RANKING order="2" place="2" resultid="14291" />
                    <RANKING order="3" place="3" resultid="15811" />
                    <RANKING order="4" place="-1" resultid="14930" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1419" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17347" />
                    <RANKING order="2" place="-1" resultid="18300" />
                    <RANKING order="3" place="-1" resultid="15817" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1420" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14827" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1421" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1422" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19433" daytime="16:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19434" daytime="16:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19435" daytime="16:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19436" daytime="16:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19437" daytime="16:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19438" daytime="16:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19439" daytime="16:45" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19440" daytime="16:45" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="19441" daytime="16:45" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="19442" daytime="16:50" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="19443" daytime="16:50" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1491" daytime="18:05" gender="F" number="28" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1492" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18603" />
                    <RANKING order="2" place="2" resultid="16583" />
                    <RANKING order="3" place="3" resultid="18203" />
                    <RANKING order="4" place="4" resultid="16543" />
                    <RANKING order="5" place="5" resultid="14880" />
                    <RANKING order="6" place="6" resultid="16595" />
                    <RANKING order="7" place="7" resultid="16604" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1493" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14838" />
                    <RANKING order="2" place="2" resultid="17593" />
                    <RANKING order="3" place="3" resultid="17380" />
                    <RANKING order="4" place="4" resultid="14574" />
                    <RANKING order="5" place="-1" resultid="17950" />
                    <RANKING order="6" place="-1" resultid="14649" />
                    <RANKING order="7" place="-1" resultid="18099" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1494" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16601" />
                    <RANKING order="2" place="2" resultid="18364" />
                    <RANKING order="3" place="3" resultid="14872" />
                    <RANKING order="4" place="4" resultid="17384" />
                    <RANKING order="5" place="5" resultid="18356" />
                    <RANKING order="6" place="6" resultid="16920" />
                    <RANKING order="7" place="7" resultid="18426" />
                    <RANKING order="8" place="8" resultid="14759" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1495" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15854" />
                    <RANKING order="2" place="2" resultid="17932" />
                    <RANKING order="3" place="3" resultid="15868" />
                    <RANKING order="4" place="4" resultid="17498" />
                    <RANKING order="5" place="5" resultid="15957" />
                    <RANKING order="6" place="6" resultid="16169" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1496" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16010" />
                    <RANKING order="2" place="2" resultid="16018" />
                    <RANKING order="3" place="3" resultid="15350" />
                    <RANKING order="4" place="4" resultid="17774" />
                    <RANKING order="5" place="5" resultid="14893" />
                    <RANKING order="6" place="6" resultid="16981" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1497" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14682" />
                    <RANKING order="2" place="2" resultid="17333" />
                    <RANKING order="3" place="3" resultid="17103" />
                    <RANKING order="4" place="4" resultid="14812" />
                    <RANKING order="5" place="5" resultid="16290" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1498" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15797" />
                    <RANKING order="2" place="2" resultid="18107" />
                    <RANKING order="3" place="3" resultid="17421" />
                    <RANKING order="4" place="4" resultid="17207" />
                    <RANKING order="5" place="-1" resultid="16536" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1499" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16152" />
                    <RANKING order="2" place="2" resultid="18432" />
                    <RANKING order="3" place="3" resultid="16353" />
                    <RANKING order="4" place="4" resultid="14489" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1500" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17157" />
                    <RANKING order="2" place="2" resultid="14373" />
                    <RANKING order="3" place="3" resultid="14848" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1501" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17728" />
                    <RANKING order="2" place="2" resultid="14494" />
                    <RANKING order="3" place="3" resultid="15029" />
                    <RANKING order="4" place="-1" resultid="17438" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1502" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14407" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1503" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1504" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1505" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="18314" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1506" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1507" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19479" daytime="18:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19480" daytime="18:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19481" daytime="18:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19482" daytime="18:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19483" daytime="18:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19484" daytime="18:30" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1525" daytime="19:30" gender="F" number="30" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="16660" agemax="99" agemin="80" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16639" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16661" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="18015" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16662" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17519" />
                    <RANKING order="2" place="2" resultid="17872" />
                    <RANKING order="3" place="-1" resultid="14903" />
                    <RANKING order="4" place="-1" resultid="15432" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16663" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17656" />
                    <RANKING order="2" place="2" resultid="18229" />
                    <RANKING order="3" place="3" resultid="15968" />
                    <RANKING order="4" place="-1" resultid="15367" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16664" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15305" />
                    <RANKING order="2" place="2" resultid="16487" />
                    <RANKING order="3" place="-1" resultid="17244" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16665" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16488" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16666" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14536" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19497" daytime="19:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19498" daytime="19:30" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1388" daytime="16:05" gender="F" number="22" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1390" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17236" />
                    <RANKING order="2" place="2" resultid="15023" />
                    <RANKING order="3" place="3" resultid="15732" />
                    <RANKING order="4" place="4" resultid="15847" />
                    <RANKING order="5" place="5" resultid="14879" />
                    <RANKING order="6" place="6" resultid="14794" />
                    <RANKING order="7" place="7" resultid="16542" />
                    <RANKING order="8" place="-1" resultid="18579" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1391" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16751" />
                    <RANKING order="2" place="2" resultid="14994" />
                    <RANKING order="3" place="-1" resultid="14584" />
                    <RANKING order="4" place="-1" resultid="17949" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1392" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17035" />
                    <RANKING order="2" place="2" resultid="18397" />
                    <RANKING order="3" place="3" resultid="17428" />
                    <RANKING order="4" place="4" resultid="17788" />
                    <RANKING order="5" place="5" resultid="14779" />
                    <RANKING order="6" place="6" resultid="17688" />
                    <RANKING order="7" place="7" resultid="15429" />
                    <RANKING order="8" place="8" resultid="18355" />
                    <RANKING order="9" place="9" resultid="14758" />
                    <RANKING order="10" place="-1" resultid="17362" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1393" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17702" />
                    <RANKING order="2" place="2" resultid="16062" />
                    <RANKING order="3" place="3" resultid="17646" />
                    <RANKING order="4" place="4" resultid="15951" />
                    <RANKING order="5" place="5" resultid="15877" />
                    <RANKING order="6" place="6" resultid="15414" />
                    <RANKING order="7" place="7" resultid="16168" />
                    <RANKING order="8" place="8" resultid="16286" />
                    <RANKING order="9" place="-1" resultid="15419" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1394" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17463" />
                    <RANKING order="2" place="2" resultid="17773" />
                    <RANKING order="3" place="3" resultid="15961" />
                    <RANKING order="4" place="4" resultid="18147" />
                    <RANKING order="5" place="-1" resultid="16979" />
                    <RANKING order="6" place="-1" resultid="15424" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1395" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18516" />
                    <RANKING order="2" place="2" resultid="14528" />
                    <RANKING order="3" place="3" resultid="14681" />
                    <RANKING order="4" place="4" resultid="17332" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1396" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17420" />
                    <RANKING order="2" place="2" resultid="16401" />
                    <RANKING order="3" place="3" resultid="15068" />
                    <RANKING order="4" place="4" resultid="15353" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1397" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15244" />
                    <RANKING order="2" place="2" resultid="14689" />
                    <RANKING order="3" place="3" resultid="17552" />
                    <RANKING order="4" place="4" resultid="17620" />
                    <RANKING order="5" place="5" resultid="17816" />
                    <RANKING order="6" place="6" resultid="16160" />
                    <RANKING order="7" place="7" resultid="16298" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1398" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17156" />
                    <RANKING order="2" place="2" resultid="14625" />
                    <RANKING order="3" place="3" resultid="14579" />
                    <RANKING order="4" place="4" resultid="17094" />
                    <RANKING order="5" place="5" resultid="14847" />
                    <RANKING order="6" place="6" resultid="18171" />
                    <RANKING order="7" place="-1" resultid="19744" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1399" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14471" />
                    <RANKING order="2" place="2" resultid="16407" />
                    <RANKING order="3" place="3" resultid="15028" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1400" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16343" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1401" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1402" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15792" />
                    <RANKING order="2" place="2" resultid="18306" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1403" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1404" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1405" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19426" daytime="16:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19427" daytime="16:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19428" daytime="16:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19429" daytime="16:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19430" daytime="16:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19431" daytime="16:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19432" daytime="16:25" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1508" daytime="18:35" gender="M" number="29" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1509" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18598" />
                    <RANKING order="2" place="2" resultid="16624" />
                    <RANKING order="3" place="3" resultid="16270" />
                    <RANKING order="4" place="4" resultid="17140" />
                    <RANKING order="5" place="5" resultid="16721" />
                    <RANKING order="6" place="6" resultid="18472" />
                    <RANKING order="7" place="-1" resultid="18054" />
                    <RANKING order="8" place="-1" resultid="18062" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1510" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15726" />
                    <RANKING order="2" place="2" resultid="17489" />
                    <RANKING order="3" place="3" resultid="15752" />
                    <RANKING order="4" place="4" resultid="18502" />
                    <RANKING order="5" place="5" resultid="16695" />
                    <RANKING order="6" place="6" resultid="16633" />
                    <RANKING order="7" place="7" resultid="17979" />
                    <RANKING order="8" place="8" resultid="16224" />
                    <RANKING order="9" place="9" resultid="16759" />
                    <RANKING order="10" place="10" resultid="17998" />
                    <RANKING order="11" place="-1" resultid="14605" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1511" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14946" />
                    <RANKING order="2" place="2" resultid="14450" />
                    <RANKING order="3" place="3" resultid="17087" />
                    <RANKING order="4" place="4" resultid="14483" />
                    <RANKING order="5" place="5" resultid="17357" />
                    <RANKING order="6" place="6" resultid="18157" />
                    <RANKING order="7" place="7" resultid="16737" />
                    <RANKING order="8" place="8" resultid="14632" />
                    <RANKING order="9" place="9" resultid="17986" />
                    <RANKING order="10" place="-1" resultid="17699" />
                    <RANKING order="11" place="-1" resultid="18392" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1512" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17173" />
                    <RANKING order="2" place="2" resultid="16827" />
                    <RANKING order="3" place="3" resultid="17706" />
                    <RANKING order="4" place="4" resultid="18208" />
                    <RANKING order="5" place="5" resultid="15335" />
                    <RANKING order="6" place="6" resultid="16812" />
                    <RANKING order="7" place="7" resultid="16733" />
                    <RANKING order="8" place="8" resultid="14556" />
                    <RANKING order="9" place="9" resultid="17044" />
                    <RANKING order="10" place="10" resultid="16941" />
                    <RANKING order="11" place="11" resultid="16282" />
                    <RANKING order="12" place="12" resultid="16766" />
                    <RANKING order="13" place="13" resultid="16302" />
                    <RANKING order="14" place="14" resultid="15034" />
                    <RANKING order="15" place="-1" resultid="14886" />
                    <RANKING order="16" place="-1" resultid="17810" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1513" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18185" />
                    <RANKING order="2" place="2" resultid="15060" />
                    <RANKING order="3" place="3" resultid="16027" />
                    <RANKING order="4" place="4" resultid="16972" />
                    <RANKING order="5" place="5" resultid="18048" />
                    <RANKING order="6" place="6" resultid="17470" />
                    <RANKING order="7" place="7" resultid="16772" />
                    <RANKING order="8" place="8" resultid="16053" />
                    <RANKING order="9" place="9" resultid="14266" />
                    <RANKING order="10" place="10" resultid="17957" />
                    <RANKING order="11" place="11" resultid="17545" />
                    <RANKING order="12" place="12" resultid="18195" />
                    <RANKING order="13" place="13" resultid="16591" />
                    <RANKING order="14" place="14" resultid="17972" />
                    <RANKING order="15" place="-1" resultid="14786" />
                    <RANKING order="16" place="-1" resultid="16841" />
                    <RANKING order="17" place="-1" resultid="17504" />
                    <RANKING order="18" place="-1" resultid="17781" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1514" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18563" />
                    <RANKING order="2" place="2" resultid="14865" />
                    <RANKING order="3" place="3" resultid="17674" />
                    <RANKING order="4" place="4" resultid="15041" />
                    <RANKING order="5" place="5" resultid="17567" />
                    <RANKING order="6" place="6" resultid="14900" />
                    <RANKING order="7" place="7" resultid="14285" />
                    <RANKING order="8" place="-1" resultid="15991" />
                    <RANKING order="9" place="-1" resultid="16134" />
                    <RANKING order="10" place="-1" resultid="16240" />
                    <RANKING order="11" place="-1" resultid="18141" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1515" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18459" />
                    <RANKING order="2" place="2" resultid="17342" />
                    <RANKING order="3" place="3" resultid="16996" />
                    <RANKING order="4" place="4" resultid="15212" />
                    <RANKING order="5" place="5" resultid="17224" />
                    <RANKING order="6" place="6" resultid="17682" />
                    <RANKING order="7" place="7" resultid="18279" />
                    <RANKING order="8" place="8" resultid="18113" />
                    <RANKING order="9" place="9" resultid="17149" />
                    <RANKING order="10" place="10" resultid="15196" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1516" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17217" />
                    <RANKING order="2" place="2" resultid="18216" />
                    <RANKING order="3" place="3" resultid="15776" />
                    <RANKING order="4" place="4" resultid="17313" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1517" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17413" />
                    <RANKING order="2" place="2" resultid="14751" />
                    <RANKING order="3" place="3" resultid="18638" />
                    <RANKING order="4" place="4" resultid="18630" />
                    <RANKING order="5" place="5" resultid="15258" />
                    <RANKING order="6" place="6" resultid="16425" />
                    <RANKING order="7" place="-1" resultid="16186" />
                    <RANKING order="8" place="-1" resultid="14442" />
                    <RANKING order="9" place="-1" resultid="18441" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1518" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17112" />
                    <RANKING order="2" place="2" resultid="14745" />
                    <RANKING order="3" place="3" resultid="14856" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1519" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14567" />
                    <RANKING order="2" place="2" resultid="16334" />
                    <RANKING order="3" place="-1" resultid="16457" />
                    <RANKING order="4" place="-1" resultid="17288" />
                    <RANKING order="5" place="-1" resultid="18332" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1520" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14455" />
                    <RANKING order="2" place="2" resultid="16180" />
                    <RANKING order="3" place="3" resultid="14931" />
                    <RANKING order="4" place="4" resultid="16445" />
                    <RANKING order="5" place="5" resultid="14390" />
                    <RANKING order="6" place="-1" resultid="17065" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1521" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="15766" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1522" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1523" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1524" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19485" daytime="18:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19486" daytime="18:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19487" daytime="18:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19488" daytime="18:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19489" daytime="19:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19490" daytime="19:05" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19491" daytime="19:10" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19492" daytime="19:10" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="19493" daytime="19:15" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="19494" daytime="19:20" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="19495" daytime="19:20" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="19496" daytime="19:25" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2017-11-19" daytime="09:00" endtime="13:21" name="BLOK IV" number="4" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="1630" daytime="09:35" gender="F" number="36" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1631" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16968" />
                    <RANKING order="2" place="2" resultid="18581" />
                    <RANKING order="3" place="-1" resultid="15409" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1632" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15738" />
                    <RANKING order="2" place="2" resultid="14586" />
                    <RANKING order="3" place="3" resultid="17511" />
                    <RANKING order="4" place="4" resultid="14832" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1633" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15002" />
                    <RANKING order="2" place="2" resultid="14873" />
                    <RANKING order="3" place="3" resultid="18366" />
                    <RANKING order="4" place="4" resultid="18357" />
                    <RANKING order="5" place="-1" resultid="18487" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1634" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17933" />
                    <RANKING order="2" place="2" resultid="18136" />
                    <RANKING order="3" place="3" resultid="15879" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1635" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15285" />
                    <RANKING order="2" place="2" resultid="16011" />
                    <RANKING order="3" place="3" resultid="14943" />
                    <RANKING order="4" place="4" resultid="15886" />
                    <RANKING order="5" place="5" resultid="17804" />
                    <RANKING order="6" place="-1" resultid="18149" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1636" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17104" />
                    <RANKING order="2" place="2" resultid="16376" />
                    <RANKING order="3" place="3" resultid="14804" />
                    <RANKING order="4" place="-1" resultid="15844" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1637" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15798" />
                    <RANKING order="2" place="2" resultid="17208" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1638" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18626" />
                    <RANKING order="2" place="2" resultid="15782" />
                    <RANKING order="3" place="3" resultid="17818" />
                    <RANKING order="4" place="4" resultid="16153" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1639" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14375" />
                    <RANKING order="2" place="2" resultid="17193" />
                    <RANKING order="3" place="3" resultid="17096" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1640" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15208" />
                    <RANKING order="2" place="2" resultid="14495" />
                    <RANKING order="3" place="3" resultid="15030" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1641" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14408" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1642" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18291" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1643" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1644" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18315" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1645" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1646" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19526" daytime="09:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19527" daytime="09:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19528" daytime="09:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19529" daytime="09:50" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1721" daytime="11:40" gender="F" number="41" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="19709" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14797" />
                    <RANKING order="2" place="2" resultid="16605" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19710" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14841" />
                    <RANKING order="2" place="2" resultid="17594" />
                    <RANKING order="3" place="3" resultid="17381" />
                    <RANKING order="4" place="-1" resultid="14652" />
                    <RANKING order="5" place="-1" resultid="18101" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19711" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17038" />
                    <RANKING order="2" place="2" resultid="18367" />
                    <RANKING order="3" place="3" resultid="17386" />
                    <RANKING order="4" place="4" resultid="18427" />
                    <RANKING order="5" place="-1" resultid="14874" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19712" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15855" />
                    <RANKING order="2" place="2" resultid="15871" />
                    <RANKING order="3" place="3" resultid="17499" />
                    <RANKING order="4" place="4" resultid="15958" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19713" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16012" />
                    <RANKING order="2" place="2" resultid="15887" />
                    <RANKING order="3" place="3" resultid="15341" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19714" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14531" />
                    <RANKING order="2" place="2" resultid="17335" />
                    <RANKING order="3" place="3" resultid="15339" />
                    <RANKING order="4" place="4" resultid="17105" />
                    <RANKING order="5" place="5" resultid="14814" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19715" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15799" />
                    <RANKING order="2" place="2" resultid="18109" />
                    <RANKING order="3" place="3" resultid="17423" />
                    <RANKING order="4" place="-1" resultid="17209" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19716" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16472" />
                    <RANKING order="2" place="2" resultid="18627" />
                    <RANKING order="3" place="3" resultid="17819" />
                    <RANKING order="4" place="4" resultid="14510" />
                    <RANKING order="5" place="5" resultid="18435" />
                    <RANKING order="6" place="6" resultid="16355" />
                    <RANKING order="7" place="7" resultid="14490" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19717" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16394" />
                    <RANKING order="2" place="2" resultid="14376" />
                    <RANKING order="3" place="3" resultid="14849" />
                    <RANKING order="4" place="4" resultid="17194" />
                    <RANKING order="5" place="5" resultid="19747" />
                    <RANKING order="6" place="6" resultid="18172" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19718" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17730" />
                    <RANKING order="2" place="2" resultid="17439" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19719" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14409" />
                    <RANKING order="2" place="-1" resultid="14461" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19720" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="19721" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="19722" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18316" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19723" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="19724" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19694" daytime="11:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19695" daytime="11:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19696" daytime="12:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19697" daytime="12:10" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="19692" daytime="12:20" gender="M" number="42" order="10" round="FHT" preveventid="1744">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="19708" daytime="12:20" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1647" daytime="09:55" gender="M" number="37" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1648" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17326" />
                    <RANKING order="2" place="2" resultid="18958" />
                    <RANKING order="3" place="3" resultid="18572" />
                    <RANKING order="4" place="-1" resultid="15020" />
                    <RANKING order="5" place="-1" resultid="18618" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1649" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17298" />
                    <RANKING order="2" place="2" resultid="15894" />
                    <RANKING order="3" place="3" resultid="15393" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1650" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18544" />
                    <RANKING order="2" place="2" resultid="16884" />
                    <RANKING order="3" place="3" resultid="15680" />
                    <RANKING order="4" place="4" resultid="17939" />
                    <RANKING order="5" place="-1" resultid="18591" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1651" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17024" />
                    <RANKING order="2" place="2" resultid="17213" />
                    <RANKING order="3" place="3" resultid="17374" />
                    <RANKING order="4" place="4" resultid="17277" />
                    <RANKING order="5" place="5" resultid="17051" />
                    <RANKING order="6" place="6" resultid="16174" />
                    <RANKING order="7" place="7" resultid="15035" />
                    <RANKING order="8" place="-1" resultid="16861" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1652" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17012" />
                    <RANKING order="2" place="2" resultid="14641" />
                    <RANKING order="3" place="3" resultid="17763" />
                    <RANKING order="4" place="4" resultid="18179" />
                    <RANKING order="5" place="5" resultid="16055" />
                    <RANKING order="6" place="-1" resultid="18531" />
                    <RANKING order="7" place="-1" resultid="16842" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1653" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14739" />
                    <RANKING order="2" place="2" resultid="14698" />
                    <RANKING order="3" place="-1" resultid="18453" />
                    <RANKING order="4" place="-1" resultid="16987" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1654" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17343" />
                    <RANKING order="2" place="2" resultid="15928" />
                    <RANKING order="3" place="3" resultid="17225" />
                    <RANKING order="4" place="4" resultid="14914" />
                    <RANKING order="5" place="5" resultid="18280" />
                    <RANKING order="6" place="6" resultid="15862" />
                    <RANKING order="7" place="7" resultid="16436" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1655" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15746" />
                    <RANKING order="2" place="2" resultid="14600" />
                    <RANKING order="3" place="3" resultid="14981" />
                    <RANKING order="4" place="4" resultid="15777" />
                    <RANKING order="5" place="5" resultid="14517" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1656" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17414" />
                    <RANKING order="2" place="2" resultid="17752" />
                    <RANKING order="3" place="3" resultid="14401" />
                    <RANKING order="4" place="4" resultid="18967" />
                    <RANKING order="5" place="5" resultid="16250" />
                    <RANKING order="6" place="6" resultid="15940" />
                    <RANKING order="7" place="7" resultid="15261" />
                    <RANKING order="8" place="8" resultid="16426" />
                    <RANKING order="9" place="-1" resultid="14443" />
                    <RANKING order="10" place="-1" resultid="16187" />
                    <RANKING order="11" place="-1" resultid="18442" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1657" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18272" />
                    <RANKING order="2" place="2" resultid="17736" />
                    <RANKING order="3" place="3" resultid="14662" />
                    <RANKING order="4" place="4" resultid="14857" />
                    <RANKING order="5" place="5" resultid="17059" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1658" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14500" />
                    <RANKING order="2" place="2" resultid="17743" />
                    <RANKING order="3" place="3" resultid="16451" />
                    <RANKING order="4" place="4" resultid="14417" />
                    <RANKING order="5" place="-1" resultid="16458" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1659" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14385" />
                    <RANKING order="2" place="2" resultid="14932" />
                    <RANKING order="3" place="3" resultid="17066" />
                    <RANKING order="4" place="4" resultid="14391" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1660" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18302" />
                    <RANKING order="2" place="2" resultid="15767" />
                    <RANKING order="3" place="3" resultid="17349" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1661" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1662" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1663" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19530" daytime="09:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19531" daytime="10:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19532" daytime="10:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19533" daytime="10:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19534" daytime="10:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19535" daytime="10:25" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19536" daytime="10:30" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19537" daytime="10:35" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1595" daytime="09:00" gender="F" number="34" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1597" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17946" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1598" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14575" />
                    <RANKING order="2" place="-1" resultid="14651" />
                    <RANKING order="3" place="-1" resultid="18100" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1599" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17966" />
                    <RANKING order="2" place="2" resultid="17385" />
                    <RANKING order="3" place="3" resultid="16921" />
                    <RANKING order="4" place="-1" resultid="17483" />
                    <RANKING order="5" place="-1" resultid="18486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1600" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17447" />
                    <RANKING order="2" place="2" resultid="14594" />
                    <RANKING order="3" place="3" resultid="16795" />
                    <RANKING order="4" place="4" resultid="15870" />
                    <RANKING order="5" place="5" resultid="16064" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1601" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16019" />
                    <RANKING order="2" place="2" resultid="15964" />
                    <RANKING order="3" place="-1" resultid="17637" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1602" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15241" />
                    <RANKING order="2" place="2" resultid="16463" />
                    <RANKING order="3" place="3" resultid="16375" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1603" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17600" />
                    <RANKING order="2" place="2" resultid="16403" />
                    <RANKING order="3" place="3" resultid="15070" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1604" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15228" />
                    <RANKING order="2" place="2" resultid="14691" />
                    <RANKING order="3" place="3" resultid="16471" />
                    <RANKING order="4" place="4" resultid="18434" />
                    <RANKING order="5" place="5" resultid="16162" />
                    <RANKING order="6" place="-1" resultid="16354" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1605" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16393" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1606" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1607" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16345" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1608" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1609" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1610" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1611" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1612" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19513" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19514" daytime="09:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19515" daytime="09:05" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1744" daytime="12:25" gender="M" number="42" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="19725" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16218" />
                    <RANKING order="2" place="2" resultid="14769" />
                    <RANKING order="3" place="3" resultid="18343" />
                    <RANKING order="4" place="-1" resultid="16273" />
                    <RANKING order="5" place="-1" resultid="16626" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19726" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16698" />
                    <RANKING order="2" place="2" resultid="18505" />
                    <RANKING order="3" place="3" resultid="15727" />
                    <RANKING order="4" place="4" resultid="17981" />
                    <RANKING order="5" place="5" resultid="16760" />
                    <RANKING order="6" place="-1" resultid="15439" />
                    <RANKING order="7" place="-1" resultid="16634" />
                    <RANKING order="8" place="-1" resultid="17299" />
                    <RANKING order="9" place="-1" resultid="17999" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19727" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14947" />
                    <RANKING order="2" place="2" resultid="17089" />
                    <RANKING order="3" place="3" resultid="14484" />
                    <RANKING order="4" place="4" resultid="17359" />
                    <RANKING order="5" place="5" resultid="15449" />
                    <RANKING order="6" place="6" resultid="16738" />
                    <RANKING order="7" place="7" resultid="15681" />
                    <RANKING order="8" place="8" resultid="14633" />
                    <RANKING order="9" place="9" resultid="17987" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19728" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17176" />
                    <RANKING order="2" place="2" resultid="18210" />
                    <RANKING order="3" place="3" resultid="17584" />
                    <RANKING order="4" place="4" resultid="17495" />
                    <RANKING order="5" place="5" resultid="15336" />
                    <RANKING order="6" place="6" resultid="16734" />
                    <RANKING order="7" place="7" resultid="17046" />
                    <RANKING order="8" place="8" resultid="16175" />
                    <RANKING order="9" place="9" resultid="16767" />
                    <RANKING order="10" place="-1" resultid="16828" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19729" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18188" />
                    <RANKING order="2" place="2" resultid="15062" />
                    <RANKING order="3" place="3" resultid="16974" />
                    <RANKING order="4" place="4" resultid="17471" />
                    <RANKING order="5" place="5" resultid="14642" />
                    <RANKING order="6" place="6" resultid="17764" />
                    <RANKING order="7" place="7" resultid="16056" />
                    <RANKING order="8" place="8" resultid="14951" />
                    <RANKING order="9" place="9" resultid="17959" />
                    <RANKING order="10" place="10" resultid="18197" />
                    <RANKING order="11" place="-1" resultid="14788" />
                    <RANKING order="12" place="-1" resultid="16843" />
                    <RANKING order="13" place="-1" resultid="16937" />
                    <RANKING order="14" place="-1" resultid="17783" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19730" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18564" />
                    <RANKING order="2" place="2" resultid="16135" />
                    <RANKING order="3" place="3" resultid="14867" />
                    <RANKING order="4" place="4" resultid="17569" />
                    <RANKING order="5" place="5" resultid="14711" />
                    <RANKING order="6" place="6" resultid="18142" />
                    <RANKING order="7" place="7" resultid="14286" />
                    <RANKING order="8" place="-1" resultid="15992" />
                    <RANKING order="9" place="-1" resultid="16242" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19731" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18461" />
                    <RANKING order="2" place="2" resultid="16997" />
                    <RANKING order="3" place="3" resultid="17226" />
                    <RANKING order="4" place="4" resultid="18281" />
                    <RANKING order="5" place="5" resultid="16131" />
                    <RANKING order="6" place="6" resultid="18114" />
                    <RANKING order="7" place="-1" resultid="17151" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19732" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17218" />
                    <RANKING order="2" place="2" resultid="18219" />
                    <RANKING order="3" place="3" resultid="18122" />
                    <RANKING order="4" place="4" resultid="16328" />
                    <RANKING order="5" place="-1" resultid="14354" />
                    <RANKING order="6" place="-1" resultid="15778" />
                    <RANKING order="7" place="-1" resultid="16234" />
                    <RANKING order="8" place="-1" resultid="17315" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19733" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14752" />
                    <RANKING order="2" place="2" resultid="14444" />
                    <RANKING order="3" place="3" resultid="18639" />
                    <RANKING order="4" place="4" resultid="18631" />
                    <RANKING order="5" place="5" resultid="16188" />
                    <RANKING order="6" place="6" resultid="18968" />
                    <RANKING order="7" place="7" resultid="14434" />
                    <RANKING order="8" place="-1" resultid="14669" />
                    <RANKING order="9" place="-1" resultid="15252" />
                    <RANKING order="10" place="-1" resultid="17753" />
                    <RANKING order="11" place="-1" resultid="18443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19734" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17114" />
                    <RANKING order="2" place="2" resultid="17737" />
                    <RANKING order="3" place="3" resultid="15221" />
                    <RANKING order="4" place="4" resultid="14746" />
                    <RANKING order="5" place="5" resultid="14858" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19735" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16337" />
                    <RANKING order="2" place="2" resultid="15268" />
                    <RANKING order="3" place="3" resultid="18334" />
                    <RANKING order="4" place="-1" resultid="14569" />
                    <RANKING order="5" place="-1" resultid="17290" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19736" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14933" />
                    <RANKING order="2" place="2" resultid="16447" />
                    <RANKING order="3" place="3" resultid="14392" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19737" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="19738" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="19739" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="19740" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19699" daytime="12:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19700" daytime="12:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19701" daytime="12:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19702" daytime="12:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19703" daytime="13:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19704" daytime="13:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19705" daytime="13:15" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19706" daytime="13:20" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="19707" daytime="13:30" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1681" daytime="10:55" gender="M" number="39" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1682" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14768" />
                    <RANKING order="2" place="2" resultid="17433" />
                    <RANKING order="3" place="3" resultid="14775" />
                    <RANKING order="4" place="4" resultid="17849" />
                    <RANKING order="5" place="5" resultid="16217" />
                    <RANKING order="6" place="6" resultid="18959" />
                    <RANKING order="7" place="7" resultid="17845" />
                    <RANKING order="8" place="8" resultid="18573" />
                    <RANKING order="9" place="9" resultid="16264" />
                    <RANKING order="10" place="10" resultid="16723" />
                    <RANKING order="11" place="-1" resultid="15021" />
                    <RANKING order="12" place="-1" resultid="17281" />
                    <RANKING order="13" place="-1" resultid="18056" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1683" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16927" />
                    <RANKING order="2" place="2" resultid="16728" />
                    <RANKING order="3" place="3" resultid="17827" />
                    <RANKING order="4" place="4" resultid="18496" />
                    <RANKING order="5" place="5" resultid="14271" />
                    <RANKING order="6" place="6" resultid="15394" />
                    <RANKING order="7" place="7" resultid="15754" />
                    <RANKING order="8" place="8" resultid="14676" />
                    <RANKING order="9" place="9" resultid="17980" />
                    <RANKING order="10" place="10" resultid="15459" />
                    <RANKING order="11" place="11" resultid="16144" />
                    <RANKING order="12" place="-1" resultid="15385" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1684" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18372" />
                    <RANKING order="2" place="2" resultid="15903" />
                    <RANKING order="3" place="3" resultid="17088" />
                    <RANKING order="4" place="4" resultid="18394" />
                    <RANKING order="5" place="5" resultid="17306" />
                    <RANKING order="6" place="6" resultid="17913" />
                    <RANKING order="7" place="7" resultid="17921" />
                    <RANKING order="8" place="8" resultid="17443" />
                    <RANKING order="9" place="9" resultid="18384" />
                    <RANKING order="10" place="10" resultid="17082" />
                    <RANKING order="11" place="-1" resultid="16617" />
                    <RANKING order="12" place="-1" resultid="16885" />
                    <RANKING order="13" place="-1" resultid="18004" />
                    <RANKING order="14" place="-1" resultid="18130" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1685" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17694" />
                    <RANKING order="2" place="2" resultid="17201" />
                    <RANKING order="3" place="3" resultid="17417" />
                    <RANKING order="4" place="4" resultid="15299" />
                    <RANKING order="5" place="5" resultid="17175" />
                    <RANKING order="6" place="6" resultid="16807" />
                    <RANKING order="7" place="7" resultid="17187" />
                    <RANKING order="8" place="8" resultid="18379" />
                    <RANKING order="9" place="9" resultid="17375" />
                    <RANKING order="10" place="10" resultid="17811" />
                    <RANKING order="11" place="11" resultid="16862" />
                    <RANKING order="12" place="12" resultid="16817" />
                    <RANKING order="13" place="13" resultid="16813" />
                    <RANKING order="14" place="14" resultid="16877" />
                    <RANKING order="15" place="15" resultid="16849" />
                    <RANKING order="16" place="16" resultid="16942" />
                    <RANKING order="17" place="17" resultid="15036" />
                    <RANKING order="18" place="-1" resultid="14558" />
                    <RANKING order="19" place="-1" resultid="14821" />
                    <RANKING order="20" place="-1" resultid="14887" />
                    <RANKING order="21" place="-1" resultid="15911" />
                    <RANKING order="22" place="-1" resultid="16360" />
                    <RANKING order="23" place="-1" resultid="16854" />
                    <RANKING order="24" place="-1" resultid="16872" />
                    <RANKING order="25" place="-1" resultid="17137" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1686" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18559" />
                    <RANKING order="2" place="2" resultid="17823" />
                    <RANKING order="3" place="3" resultid="17589" />
                    <RANKING order="4" place="4" resultid="16029" />
                    <RANKING order="5" place="5" resultid="17407" />
                    <RANKING order="6" place="6" resultid="16047" />
                    <RANKING order="7" place="7" resultid="14279" />
                    <RANKING order="8" place="8" resultid="17782" />
                    <RANKING order="9" place="9" resultid="17798" />
                    <RANKING order="10" place="10" resultid="17958" />
                    <RANKING order="11" place="11" resultid="14938" />
                    <RANKING order="12" place="12" resultid="14724" />
                    <RANKING order="13" place="-1" resultid="14787" />
                    <RANKING order="14" place="-1" resultid="15357" />
                    <RANKING order="15" place="-1" resultid="15454" />
                    <RANKING order="16" place="-1" resultid="16319" />
                    <RANKING order="17" place="-1" resultid="17401" />
                    <RANKING order="18" place="-1" resultid="17546" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1687" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17617" />
                    <RANKING order="2" place="2" resultid="14970" />
                    <RANKING order="3" place="3" resultid="16072" />
                    <RANKING order="4" place="4" resultid="14866" />
                    <RANKING order="5" place="5" resultid="16038" />
                    <RANKING order="6" place="6" resultid="16440" />
                    <RANKING order="7" place="7" resultid="14710" />
                    <RANKING order="8" place="8" resultid="16081" />
                    <RANKING order="9" place="-1" resultid="16241" />
                    <RANKING order="10" place="-1" resultid="17676" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1688" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14302" />
                    <RANKING order="2" place="2" resultid="18540" />
                    <RANKING order="3" place="3" resultid="18512" />
                    <RANKING order="4" place="4" resultid="15012" />
                    <RANKING order="5" place="5" resultid="18295" />
                    <RANKING order="6" place="6" resultid="16130" />
                    <RANKING order="7" place="7" resultid="16478" />
                    <RANKING order="8" place="8" resultid="17395" />
                    <RANKING order="9" place="9" resultid="15863" />
                    <RANKING order="10" place="10" resultid="16947" />
                    <RANKING order="11" place="-1" resultid="14621" />
                    <RANKING order="12" place="-1" resultid="18551" />
                    <RANKING order="13" place="-1" resultid="16993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1689" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18286" />
                    <RANKING order="2" place="2" resultid="16368" />
                    <RANKING order="3" place="3" resultid="17181" />
                    <RANKING order="4" place="4" resultid="15789" />
                    <RANKING order="5" place="5" resultid="15280" />
                    <RANKING order="6" place="6" resultid="15273" />
                    <RANKING order="7" place="7" resultid="16327" />
                    <RANKING order="8" place="-1" resultid="17321" />
                    <RANKING order="9" place="-1" resultid="18470" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1690" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14733" />
                    <RANKING order="2" place="2" resultid="15403" />
                    <RANKING order="3" place="3" resultid="15823" />
                    <RANKING order="4" place="4" resultid="16258" />
                    <RANKING order="5" place="5" resultid="16427" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1691" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17454" />
                    <RANKING order="2" place="2" resultid="15220" />
                    <RANKING order="3" place="3" resultid="14703" />
                    <RANKING order="4" place="4" resultid="18524" />
                    <RANKING order="5" place="5" resultid="15829" />
                    <RANKING order="6" place="6" resultid="15290" />
                    <RANKING order="7" place="7" resultid="15805" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1692" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14364" />
                    <RANKING order="2" place="2" resultid="18333" />
                    <RANKING order="3" place="3" resultid="17744" />
                    <RANKING order="4" place="4" resultid="15917" />
                    <RANKING order="5" place="5" resultid="16415" />
                    <RANKING order="6" place="6" resultid="14418" />
                    <RANKING order="7" place="-1" resultid="17077" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1693" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14562" />
                    <RANKING order="2" place="2" resultid="14476" />
                    <RANKING order="3" place="3" resultid="14294" />
                    <RANKING order="4" place="4" resultid="15814" />
                    <RANKING order="5" place="5" resultid="16446" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1694" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17350" />
                    <RANKING order="2" place="2" resultid="15768" />
                    <RANKING order="3" place="3" resultid="18303" />
                    <RANKING order="4" place="-1" resultid="15819" />
                    <RANKING order="5" place="-1" resultid="17070" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1695" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14828" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1696" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1697" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19546" daytime="10:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19547" daytime="10:55" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19548" daytime="11:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19549" daytime="11:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19550" daytime="11:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19551" daytime="11:05" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19552" daytime="11:05" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19553" daytime="11:05" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="19554" daytime="11:10" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="19555" daytime="11:10" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="19556" daytime="11:10" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="19557" daytime="11:15" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="19558" daytime="11:15" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="19559" daytime="11:15" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="19560" daytime="11:20" number="15" order="15" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1664" daytime="10:35" gender="F" number="38" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1665" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15024" />
                    <RANKING order="2" place="2" resultid="17238" />
                    <RANKING order="3" place="3" resultid="15733" />
                    <RANKING order="4" place="4" resultid="16610" />
                    <RANKING order="5" place="5" resultid="18582" />
                    <RANKING order="6" place="6" resultid="14881" />
                    <RANKING order="7" place="7" resultid="17907" />
                    <RANKING order="8" place="8" resultid="16544" />
                    <RANKING order="9" place="9" resultid="14796" />
                    <RANKING order="10" place="10" resultid="16596" />
                    <RANKING order="11" place="-1" resultid="15849" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1666" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14840" />
                    <RANKING order="2" place="2" resultid="16753" />
                    <RANKING order="3" place="3" resultid="17857" />
                    <RANKING order="4" place="4" resultid="14995" />
                    <RANKING order="5" place="-1" resultid="17951" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1667" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18398" />
                    <RANKING order="2" place="2" resultid="15301" />
                    <RANKING order="3" place="3" resultid="15003" />
                    <RANKING order="4" place="4" resultid="17037" />
                    <RANKING order="5" place="5" resultid="17790" />
                    <RANKING order="6" place="6" resultid="17429" />
                    <RANKING order="7" place="7" resultid="14780" />
                    <RANKING order="8" place="8" resultid="17689" />
                    <RANKING order="9" place="9" resultid="15431" />
                    <RANKING order="10" place="10" resultid="18358" />
                    <RANKING order="11" place="-1" resultid="14760" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1668" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14595" />
                    <RANKING order="2" place="2" resultid="17647" />
                    <RANKING order="3" place="3" resultid="17703" />
                    <RANKING order="4" place="4" resultid="16065" />
                    <RANKING order="5" place="5" resultid="15953" />
                    <RANKING order="6" place="6" resultid="15880" />
                    <RANKING order="7" place="7" resultid="15415" />
                    <RANKING order="8" place="8" resultid="17852" />
                    <RANKING order="9" place="9" resultid="16170" />
                    <RANKING order="10" place="-1" resultid="15420" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1669" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17464" />
                    <RANKING order="2" place="2" resultid="15351" />
                    <RANKING order="3" place="3" resultid="16020" />
                    <RANKING order="4" place="4" resultid="17775" />
                    <RANKING order="5" place="5" resultid="16980" />
                    <RANKING order="6" place="6" resultid="15962" />
                    <RANKING order="7" place="-1" resultid="18150" />
                    <RANKING order="8" place="-1" resultid="15425" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1670" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18517" />
                    <RANKING order="2" place="2" resultid="14683" />
                    <RANKING order="3" place="3" resultid="17334" />
                    <RANKING order="4" place="4" resultid="15202" />
                    <RANKING order="5" place="5" resultid="15933" />
                    <RANKING order="6" place="6" resultid="14805" />
                    <RANKING order="7" place="7" resultid="15947" />
                    <RANKING order="8" place="-1" resultid="14530" />
                    <RANKING order="9" place="-1" resultid="14813" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1671" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16314" />
                    <RANKING order="2" place="2" resultid="17422" />
                    <RANKING order="3" place="3" resultid="15071" />
                    <RANKING order="4" place="4" resultid="15354" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1672" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15245" />
                    <RANKING order="2" place="2" resultid="14692" />
                    <RANKING order="3" place="3" resultid="17554" />
                    <RANKING order="4" place="4" resultid="16154" />
                    <RANKING order="5" place="5" resultid="16163" />
                    <RANKING order="6" place="-1" resultid="17621" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1673" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17158" />
                    <RANKING order="2" place="2" resultid="14627" />
                    <RANKING order="3" place="3" resultid="17606" />
                    <RANKING order="4" place="4" resultid="14580" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1674" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17729" />
                    <RANKING order="2" place="2" resultid="14472" />
                    <RANKING order="3" place="3" resultid="16409" />
                    <RANKING order="4" place="4" resultid="15031" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1675" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14468" />
                    <RANKING order="2" place="2" resultid="16346" />
                    <RANKING order="3" place="-1" resultid="14664" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1676" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1677" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15793" />
                    <RANKING order="2" place="2" resultid="18307" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1678" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1679" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1680" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19538" daytime="10:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19539" daytime="10:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19540" daytime="10:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19541" daytime="10:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19542" daytime="10:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19543" daytime="10:50" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19544" daytime="10:50" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19545" daytime="10:55" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="19690" daytime="11:35" gender="F" number="41" order="8" round="FHT" preveventid="1721">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="19698" daytime="11:35" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1698" daytime="11:20" gender="X" number="40" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="16674" agemax="99" agemin="80" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16645" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16675" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="18013" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16676" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17520" />
                    <RANKING order="2" place="2" resultid="18011" />
                    <RANKING order="3" place="3" resultid="16887" />
                    <RANKING order="4" place="4" resultid="18400" />
                    <RANKING order="5" place="5" resultid="17878" />
                    <RANKING order="6" place="6" resultid="17118" />
                    <RANKING order="7" place="7" resultid="15913" />
                    <RANKING order="8" place="8" resultid="18227" />
                    <RANKING order="9" place="-1" resultid="14905" />
                    <RANKING order="10" place="-1" resultid="16643" />
                    <RANKING order="11" place="-1" resultid="17718" />
                    <RANKING order="12" place="-1" resultid="17870" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16677" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16491" />
                    <RANKING order="2" place="2" resultid="15311" />
                    <RANKING order="3" place="3" resultid="17868" />
                    <RANKING order="4" place="4" resultid="17521" />
                    <RANKING order="5" place="5" resultid="16088" />
                    <RANKING order="6" place="6" resultid="17247" />
                    <RANKING order="7" place="7" resultid="17522" />
                    <RANKING order="8" place="8" resultid="15966" />
                    <RANKING order="9" place="-1" resultid="15365" />
                    <RANKING order="10" place="-1" resultid="18224" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16678" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17657" />
                    <RANKING order="2" place="2" resultid="14719" />
                    <RANKING order="3" place="3" resultid="15971" />
                    <RANKING order="4" place="4" resultid="16207" />
                    <RANKING order="5" place="-1" resultid="17248" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16679" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15304" />
                    <RANKING order="2" place="2" resultid="16492" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16680" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14538" />
                    <RANKING order="2" place="2" resultid="16493" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19561" daytime="11:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19562" daytime="11:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19563" daytime="11:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19564" daytime="11:30" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1613" daytime="09:10" gender="M" number="35" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1614" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16625" />
                    <RANKING order="2" place="2" resultid="16709" />
                    <RANKING order="3" place="3" resultid="16272" />
                    <RANKING order="4" place="4" resultid="17992" />
                    <RANKING order="5" place="5" resultid="18473" />
                    <RANKING order="6" place="-1" resultid="16722" />
                    <RANKING order="7" place="-1" resultid="18063" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1615" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="16715" />
                    <RANKING order="2" place="2" resultid="16746" />
                    <RANKING order="3" place="3" resultid="18504" />
                    <RANKING order="4" place="4" resultid="15753" />
                    <RANKING order="5" place="-1" resultid="14675" />
                    <RANKING order="6" place="-1" resultid="15978" />
                    <RANKING order="7" place="-1" resultid="16697" />
                    <RANKING order="8" place="-1" resultid="17490" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1616" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18478" />
                    <RANKING order="2" place="2" resultid="15902" />
                    <RANKING order="3" place="3" resultid="18393" />
                    <RANKING order="4" place="4" resultid="17920" />
                    <RANKING order="5" place="5" resultid="16547" />
                    <RANKING order="6" place="6" resultid="17358" />
                    <RANKING order="7" place="-1" resultid="15448" />
                    <RANKING order="8" place="-1" resultid="18129" />
                    <RANKING order="9" place="-1" resultid="18590" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1617" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18378" />
                    <RANKING order="2" place="2" resultid="16205" />
                    <RANKING order="3" place="3" resultid="16801" />
                    <RANKING order="4" place="4" resultid="15298" />
                    <RANKING order="5" place="5" resultid="17459" />
                    <RANKING order="6" place="6" resultid="17231" />
                    <RANKING order="7" place="7" resultid="17045" />
                    <RANKING order="8" place="8" resultid="14557" />
                    <RANKING order="9" place="-1" resultid="14820" />
                    <RANKING order="10" place="-1" resultid="15910" />
                    <RANKING order="11" place="-1" resultid="17583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1618" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15061" />
                    <RANKING order="2" place="2" resultid="16973" />
                    <RANKING order="3" place="3" resultid="18187" />
                    <RANKING order="4" place="4" resultid="16028" />
                    <RANKING order="5" place="5" resultid="18049" />
                    <RANKING order="6" place="6" resultid="17797" />
                    <RANKING order="7" place="7" resultid="18196" />
                    <RANKING order="8" place="-1" resultid="14427" />
                    <RANKING order="9" place="-1" resultid="14974" />
                    <RANKING order="10" place="-1" resultid="16046" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1619" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="17612" />
                    <RANKING order="2" place="2" resultid="18452" />
                    <RANKING order="3" place="3" resultid="17675" />
                    <RANKING order="4" place="4" resultid="16071" />
                    <RANKING order="5" place="5" resultid="15042" />
                    <RANKING order="6" place="6" resultid="16077" />
                    <RANKING order="7" place="7" resultid="17626" />
                    <RANKING order="8" place="8" resultid="16096" />
                    <RANKING order="9" place="-1" resultid="16037" />
                    <RANKING order="10" place="-1" resultid="17568" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1620" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18511" />
                    <RANKING order="2" place="2" resultid="14301" />
                    <RANKING order="3" place="3" resultid="14913" />
                    <RANKING order="4" place="4" resultid="17683" />
                    <RANKING order="5" place="5" resultid="15213" />
                    <RANKING order="6" place="6" resultid="17150" />
                    <RANKING order="7" place="7" resultid="17394" />
                    <RANKING order="8" place="-1" resultid="16435" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1621" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18218" />
                    <RANKING order="2" place="2" resultid="16367" />
                    <RANKING order="3" place="3" resultid="18321" />
                    <RANKING order="4" place="4" resultid="15788" />
                    <RANKING order="5" place="5" resultid="18121" />
                    <RANKING order="6" place="6" resultid="16233" />
                    <RANKING order="7" place="7" resultid="17314" />
                    <RANKING order="8" place="-1" resultid="15921" />
                    <RANKING order="9" place="-1" resultid="14353" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1622" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15251" />
                    <RANKING order="2" place="2" resultid="15402" />
                    <RANKING order="3" place="3" resultid="14732" />
                    <RANKING order="4" place="4" resultid="14400" />
                    <RANKING order="5" place="5" resultid="15260" />
                    <RANKING order="6" place="-1" resultid="16257" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1623" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="18271" />
                    <RANKING order="2" place="2" resultid="17113" />
                    <RANKING order="3" place="3" resultid="14661" />
                    <RANKING order="4" place="4" resultid="17058" />
                    <RANKING order="5" place="-1" resultid="14465" />
                    <RANKING order="6" place="-1" resultid="15828" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1624" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14568" />
                    <RANKING order="2" place="2" resultid="14363" />
                    <RANKING order="3" place="3" resultid="15267" />
                    <RANKING order="4" place="4" resultid="16336" />
                    <RANKING order="5" place="-1" resultid="17289" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1625" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14293" />
                    <RANKING order="2" place="2" resultid="15813" />
                    <RANKING order="3" place="3" resultid="14384" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1626" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1627" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1628" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1629" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="19516" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="19517" daytime="09:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="19518" daytime="09:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="19519" daytime="09:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="19520" daytime="09:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="19521" daytime="09:25" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="19522" daytime="09:25" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="19523" daytime="09:25" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="19524" daytime="09:30" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="19525" daytime="09:30" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" nation="POL" clubid="18087" name="AQUASFERA Masters Olsztyn">
          <CONTACT email="annamariaaneczka@uwm.edu.pl" name="Goździejewska Anna" />
          <ATHLETES>
            <ATHLETE birthdate="1974-04-01" firstname="Paweł" gender="M" lastname="Dąbrowski" nation="POL" athleteid="18173">
              <RESULTS>
                <RESULT eventid="1079" points="335" reactiontime="+83" swimtime="00:00:29.16" resultid="18174" heatid="19294" lane="8" entrytime="00:00:29.50" />
                <RESULT eventid="1205" points="251" reactiontime="+81" swimtime="00:00:35.18" resultid="18175" heatid="19348" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="14243" points="297" reactiontime="+83" swimtime="00:01:15.37" resultid="18176" heatid="19403" lane="8" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="279" reactiontime="+85" swimtime="00:00:33.36" resultid="18177" heatid="19450" lane="8" />
                <RESULT eventid="1474" points="239" reactiontime="+82" swimtime="00:01:18.77" resultid="18178" heatid="19474" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="224" reactiontime="+83" swimtime="00:02:53.88" resultid="18179" heatid="19535" lane="0" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.48" />
                    <SPLIT distance="100" swimtime="00:01:24.35" />
                    <SPLIT distance="150" swimtime="00:02:08.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-03-18" firstname="Anna" gender="F" lastname="Goździejewska" nation="POL" athleteid="18102">
              <RESULTS>
                <RESULT eventid="1062" points="295" reactiontime="+86" swimtime="00:00:34.91" resultid="18103" heatid="19280" lane="8" entrytime="00:00:33.80" />
                <RESULT eventid="1165" points="342" reactiontime="+101" swimtime="00:21:54.74" resultid="18104" heatid="19624" lane="5" entrytime="00:23:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.91" />
                    <SPLIT distance="100" swimtime="00:01:24.84" />
                    <SPLIT distance="150" swimtime="00:02:09.32" />
                    <SPLIT distance="200" swimtime="00:02:53.90" />
                    <SPLIT distance="250" swimtime="00:03:38.27" />
                    <SPLIT distance="300" swimtime="00:04:22.69" />
                    <SPLIT distance="350" swimtime="00:05:07.01" />
                    <SPLIT distance="400" swimtime="00:05:51.57" />
                    <SPLIT distance="450" swimtime="00:06:35.87" />
                    <SPLIT distance="500" swimtime="00:07:20.03" />
                    <SPLIT distance="550" swimtime="00:08:04.17" />
                    <SPLIT distance="600" swimtime="00:08:48.31" />
                    <SPLIT distance="650" swimtime="00:09:32.36" />
                    <SPLIT distance="700" swimtime="00:10:16.52" />
                    <SPLIT distance="750" swimtime="00:11:00.48" />
                    <SPLIT distance="800" swimtime="00:11:44.32" />
                    <SPLIT distance="850" swimtime="00:12:28.07" />
                    <SPLIT distance="900" swimtime="00:13:11.79" />
                    <SPLIT distance="950" swimtime="00:13:55.43" />
                    <SPLIT distance="1000" swimtime="00:14:39.14" />
                    <SPLIT distance="1050" swimtime="00:15:22.58" />
                    <SPLIT distance="1100" swimtime="00:16:06.01" />
                    <SPLIT distance="1150" swimtime="00:16:49.94" />
                    <SPLIT distance="1200" swimtime="00:17:33.48" />
                    <SPLIT distance="1250" swimtime="00:18:17.18" />
                    <SPLIT distance="1300" swimtime="00:19:01.12" />
                    <SPLIT distance="1350" swimtime="00:19:44.91" />
                    <SPLIT distance="1400" swimtime="00:20:29.08" />
                    <SPLIT distance="1450" swimtime="00:21:12.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="246" reactiontime="+91" swimtime="00:03:34.73" resultid="18105" heatid="19357" lane="8" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.28" />
                    <SPLIT distance="100" swimtime="00:01:46.48" />
                    <SPLIT distance="150" swimtime="00:02:41.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="303" reactiontime="+88" swimtime="00:01:15.73" resultid="18106" heatid="19370" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="314" reactiontime="+89" swimtime="00:02:42.87" resultid="18107" heatid="19480" lane="5" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.59" />
                    <SPLIT distance="100" swimtime="00:01:20.51" />
                    <SPLIT distance="150" swimtime="00:02:02.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="249" reactiontime="+92" swimtime="00:06:52.26" resultid="18108" heatid="19504" lane="8" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.64" />
                    <SPLIT distance="100" swimtime="00:01:43.84" />
                    <SPLIT distance="150" swimtime="00:02:37.31" />
                    <SPLIT distance="200" swimtime="00:03:30.49" />
                    <SPLIT distance="250" swimtime="00:04:27.23" />
                    <SPLIT distance="300" swimtime="00:05:24.14" />
                    <SPLIT distance="350" swimtime="00:06:08.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="342" reactiontime="+87" swimtime="00:05:35.15" resultid="18109" heatid="19697" lane="4" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.17" />
                    <SPLIT distance="100" swimtime="00:01:21.16" />
                    <SPLIT distance="150" swimtime="00:02:03.83" />
                    <SPLIT distance="200" swimtime="00:02:46.72" />
                    <SPLIT distance="250" swimtime="00:03:29.69" />
                    <SPLIT distance="300" swimtime="00:04:12.30" />
                    <SPLIT distance="350" swimtime="00:04:54.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-09-01" firstname="Grzegorz" gender="M" lastname="Mówiński" nation="POL" athleteid="18220">
              <RESULTS>
                <RESULT eventid="14189" points="225" reactiontime="+105" swimtime="00:12:08.33" resultid="18221" heatid="19616" lane="1" entrytime="00:12:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.43" />
                    <SPLIT distance="100" swimtime="00:01:23.23" />
                    <SPLIT distance="150" swimtime="00:02:08.44" />
                    <SPLIT distance="200" swimtime="00:02:53.88" />
                    <SPLIT distance="250" swimtime="00:03:40.25" />
                    <SPLIT distance="300" swimtime="00:04:26.75" />
                    <SPLIT distance="350" swimtime="00:05:13.09" />
                    <SPLIT distance="400" swimtime="00:05:59.85" />
                    <SPLIT distance="450" swimtime="00:06:46.89" />
                    <SPLIT distance="500" swimtime="00:07:33.64" />
                    <SPLIT distance="550" swimtime="00:08:20.65" />
                    <SPLIT distance="600" swimtime="00:09:07.62" />
                    <SPLIT distance="650" swimtime="00:09:54.35" />
                    <SPLIT distance="700" swimtime="00:10:40.75" />
                    <SPLIT distance="750" swimtime="00:11:25.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="205" reactiontime="+93" swimtime="00:03:03.97" resultid="18222" heatid="19415" lane="3" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.06" />
                    <SPLIT distance="100" swimtime="00:01:27.90" />
                    <SPLIT distance="150" swimtime="00:02:16.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="206" reactiontime="+90" swimtime="00:06:38.38" resultid="18223" heatid="19508" lane="2" entrytime="00:07:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.97" />
                    <SPLIT distance="100" swimtime="00:01:30.49" />
                    <SPLIT distance="150" swimtime="00:02:28.04" />
                    <SPLIT distance="200" swimtime="00:03:23.04" />
                    <SPLIT distance="250" swimtime="00:04:18.63" />
                    <SPLIT distance="300" swimtime="00:05:13.16" />
                    <SPLIT distance="350" swimtime="00:05:58.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-08-31" firstname="Iwona" gender="F" lastname="Bardzicka" nation="POL" athleteid="18169">
              <RESULTS>
                <RESULT eventid="1222" points="102" swimtime="00:04:47.73" resultid="18170" heatid="19354" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.61" />
                    <SPLIT distance="100" swimtime="00:02:16.16" />
                    <SPLIT distance="150" swimtime="00:03:31.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="96" swimtime="00:02:16.08" resultid="18171" heatid="19427" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="48" swimtime="00:10:41.50" resultid="18172" heatid="19694" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.44" />
                    <SPLIT distance="100" swimtime="00:02:30.58" />
                    <SPLIT distance="150" swimtime="00:03:53.03" />
                    <SPLIT distance="200" swimtime="00:05:13.40" />
                    <SPLIT distance="250" swimtime="00:06:38.65" />
                    <SPLIT distance="300" swimtime="00:07:58.30" />
                    <SPLIT distance="350" swimtime="00:09:23.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-06-25" firstname="Adam" gender="M" lastname="Matusiak vel Matuszewski" nation="POL" athleteid="18189">
              <RESULTS>
                <RESULT eventid="1079" points="213" reactiontime="+88" swimtime="00:00:33.92" resultid="18190" heatid="19288" lane="0" entrytime="00:00:35.12" />
                <RESULT eventid="14207" reactiontime="+92" status="OTL" swimtime="00:23:51.45" resultid="18191" heatid="19622" lane="9" entrytime="00:23:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.19" />
                    <SPLIT distance="100" swimtime="00:01:26.30" />
                    <SPLIT distance="150" swimtime="00:02:13.37" />
                    <SPLIT distance="200" swimtime="00:03:01.79" />
                    <SPLIT distance="250" swimtime="00:03:51.72" />
                    <SPLIT distance="300" swimtime="00:04:41.56" />
                    <SPLIT distance="350" swimtime="00:05:31.41" />
                    <SPLIT distance="400" swimtime="00:06:20.65" />
                    <SPLIT distance="450" swimtime="00:07:10.56" />
                    <SPLIT distance="500" swimtime="00:08:00.32" />
                    <SPLIT distance="550" swimtime="00:08:49.33" />
                    <SPLIT distance="600" swimtime="00:09:38.98" />
                    <SPLIT distance="650" swimtime="00:10:29.22" />
                    <SPLIT distance="700" swimtime="00:11:19.52" />
                    <SPLIT distance="750" swimtime="00:12:10.25" />
                    <SPLIT distance="800" swimtime="00:13:00.79" />
                    <SPLIT distance="850" swimtime="00:13:52.13" />
                    <SPLIT distance="900" swimtime="00:14:43.20" />
                    <SPLIT distance="950" swimtime="00:15:34.54" />
                    <SPLIT distance="1000" swimtime="00:16:25.36" />
                    <SPLIT distance="1050" swimtime="00:17:16.09" />
                    <SPLIT distance="1100" swimtime="00:18:06.74" />
                    <SPLIT distance="1150" swimtime="00:18:57.54" />
                    <SPLIT distance="1200" swimtime="00:19:48.19" />
                    <SPLIT distance="1250" swimtime="00:20:38.60" />
                    <SPLIT distance="1300" swimtime="00:21:28.76" />
                    <SPLIT distance="1350" swimtime="00:22:18.61" />
                    <SPLIT distance="1400" swimtime="00:23:09.46" />
                    <SPLIT distance="1450" swimtime="00:23:10.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="107" reactiontime="+76" swimtime="00:00:46.68" resultid="18192" heatid="19342" lane="6" />
                <RESULT eventid="1273" points="212" reactiontime="+90" swimtime="00:01:15.36" resultid="18193" heatid="19377" lane="5" entrytime="00:01:19.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="140" reactiontime="+85" swimtime="00:00:41.90" resultid="18194" heatid="19452" lane="7" entrytime="00:00:42.87" />
                <RESULT eventid="1508" points="185" reactiontime="+102" swimtime="00:02:54.35" resultid="18195" heatid="19489" lane="1" entrytime="00:02:54.08">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="90" reactiontime="+102" swimtime="00:01:47.17" resultid="18196" heatid="19516" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="176" reactiontime="+91" swimtime="00:06:18.53" resultid="18197" heatid="19702" lane="7" entrytime="00:06:17.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.92" />
                    <SPLIT distance="100" swimtime="00:01:30.43" />
                    <SPLIT distance="150" swimtime="00:02:19.94" />
                    <SPLIT distance="200" swimtime="00:03:09.71" />
                    <SPLIT distance="250" swimtime="00:03:59.82" />
                    <SPLIT distance="300" swimtime="00:04:49.52" />
                    <SPLIT distance="350" swimtime="00:05:36.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-02-15" firstname="Jowita" gender="F" lastname="Kucharska" nation="POL" athleteid="18131">
              <RESULTS>
                <RESULT eventid="1062" points="359" reactiontime="+86" swimtime="00:00:32.67" resultid="18132" heatid="19281" lane="8" entrytime="00:00:32.50" />
                <RESULT eventid="1096" points="292" reactiontime="+86" swimtime="00:03:03.60" resultid="18133" heatid="19307" lane="6" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.59" />
                    <SPLIT distance="100" swimtime="00:01:27.76" />
                    <SPLIT distance="150" swimtime="00:02:24.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="353" reactiontime="+84" swimtime="00:01:12.01" resultid="18134" heatid="19370" lane="3" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="315" reactiontime="+84" swimtime="00:00:35.82" resultid="18135" heatid="19447" lane="5" entrytime="00:00:36.00" />
                <RESULT eventid="1630" points="261" swimtime="00:03:06.49" resultid="18136" heatid="19528" lane="7" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.91" />
                    <SPLIT distance="100" swimtime="00:01:31.08" />
                    <SPLIT distance="150" swimtime="00:02:19.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-02-09" firstname="Aleksandra" gender="F" lastname="Milewska" nation="POL" athleteid="18198">
              <RESULTS>
                <RESULT eventid="1062" points="391" reactiontime="+85" swimtime="00:00:31.78" resultid="18199" heatid="19281" lane="7" entrytime="00:00:32.30" />
                <RESULT eventid="1147" reactiontime="+81" status="OTL" swimtime="00:12:03.48" resultid="18200" heatid="19596" lane="8" entrytime="00:11:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                    <SPLIT distance="100" swimtime="00:01:18.06" />
                    <SPLIT distance="150" swimtime="00:02:00.36" />
                    <SPLIT distance="200" swimtime="00:02:44.80" />
                    <SPLIT distance="250" swimtime="00:03:29.93" />
                    <SPLIT distance="300" swimtime="00:04:16.32" />
                    <SPLIT distance="350" swimtime="00:05:02.51" />
                    <SPLIT distance="400" swimtime="00:05:48.51" />
                    <SPLIT distance="450" swimtime="00:06:35.36" />
                    <SPLIT distance="500" swimtime="00:07:21.89" />
                    <SPLIT distance="550" swimtime="00:08:08.73" />
                    <SPLIT distance="600" swimtime="00:08:55.51" />
                    <SPLIT distance="650" swimtime="00:09:42.89" />
                    <SPLIT distance="700" swimtime="00:10:30.04" />
                    <SPLIT distance="750" swimtime="00:11:16.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="299" reactiontime="+90" swimtime="00:03:21.13" resultid="18201" heatid="19357" lane="5" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.63" />
                    <SPLIT distance="100" swimtime="00:01:37.93" />
                    <SPLIT distance="150" swimtime="00:02:29.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="369" reactiontime="+89" swimtime="00:00:33.99" resultid="18202" heatid="19448" lane="1" entrytime="00:00:33.80" />
                <RESULT eventid="1491" points="348" reactiontime="+89" swimtime="00:02:37.49" resultid="18203" heatid="19483" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.38" />
                    <SPLIT distance="100" swimtime="00:01:16.30" />
                    <SPLIT distance="150" swimtime="00:01:57.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-02-18" firstname="Bogdan" gender="M" lastname="Milewski" nation="POL" athleteid="18137">
              <RESULTS>
                <RESULT eventid="1079" points="255" reactiontime="+89" swimtime="00:00:31.92" resultid="18138" heatid="19291" lane="3" entrytime="00:00:31.25" />
                <RESULT eventid="1239" points="217" reactiontime="+85" swimtime="00:03:20.35" resultid="18139" heatid="19362" lane="0" entrytime="00:03:15.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.10" />
                    <SPLIT distance="100" swimtime="00:01:34.29" />
                    <SPLIT distance="150" swimtime="00:02:27.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="249" reactiontime="+98" swimtime="00:01:28.29" resultid="18140" heatid="19438" lane="1" entrytime="00:01:27.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="18141" heatid="19490" lane="1" entrytime="00:02:45.00" />
                <RESULT eventid="1744" points="176" reactiontime="+89" swimtime="00:06:18.22" resultid="18142" heatid="19703" lane="9" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.59" />
                    <SPLIT distance="100" swimtime="00:01:27.39" />
                    <SPLIT distance="150" swimtime="00:02:13.75" />
                    <SPLIT distance="200" swimtime="00:03:02.51" />
                    <SPLIT distance="250" swimtime="00:03:52.60" />
                    <SPLIT distance="300" swimtime="00:04:41.25" />
                    <SPLIT distance="350" swimtime="00:05:30.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-30" firstname="Paweł" gender="M" lastname="Gregorowicz" nation="POL" athleteid="18180">
              <RESULTS>
                <RESULT eventid="1079" points="473" reactiontime="+75" swimtime="00:00:26.00" resultid="18181" heatid="19299" lane="0" entrytime="00:00:27.20" />
                <RESULT eventid="14189" points="491" reactiontime="+83" swimtime="00:09:22.06" resultid="18182" heatid="19618" lane="6" entrytime="00:09:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.41" />
                    <SPLIT distance="100" swimtime="00:01:05.98" />
                    <SPLIT distance="150" swimtime="00:01:41.15" />
                    <SPLIT distance="200" swimtime="00:02:16.70" />
                    <SPLIT distance="250" swimtime="00:02:52.11" />
                    <SPLIT distance="300" swimtime="00:03:27.56" />
                    <SPLIT distance="350" swimtime="00:04:03.03" />
                    <SPLIT distance="400" swimtime="00:04:38.67" />
                    <SPLIT distance="450" swimtime="00:05:14.19" />
                    <SPLIT distance="500" swimtime="00:05:49.74" />
                    <SPLIT distance="550" swimtime="00:06:25.36" />
                    <SPLIT distance="600" swimtime="00:07:01.00" />
                    <SPLIT distance="650" swimtime="00:07:36.40" />
                    <SPLIT distance="700" swimtime="00:08:12.00" />
                    <SPLIT distance="750" swimtime="00:08:47.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="496" reactiontime="+78" swimtime="00:00:56.76" resultid="18183" heatid="19386" lane="4" entrytime="00:00:57.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="421" reactiontime="+72" swimtime="00:01:07.10" resultid="18184" heatid="19407" lane="9" entrytime="00:01:08.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="499" reactiontime="+78" swimtime="00:02:05.21" resultid="18185" heatid="19495" lane="5" entrytime="00:02:05.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.56" />
                    <SPLIT distance="100" swimtime="00:01:01.36" />
                    <SPLIT distance="150" swimtime="00:01:33.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="412" reactiontime="+80" swimtime="00:05:16.34" resultid="18186" heatid="19511" lane="5" entrytime="00:05:28.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                    <SPLIT distance="100" swimtime="00:01:09.06" />
                    <SPLIT distance="150" swimtime="00:01:53.34" />
                    <SPLIT distance="200" swimtime="00:02:35.10" />
                    <SPLIT distance="250" swimtime="00:03:20.52" />
                    <SPLIT distance="300" swimtime="00:04:06.00" />
                    <SPLIT distance="350" swimtime="00:04:42.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="440" reactiontime="+78" swimtime="00:01:03.21" resultid="18187" heatid="19523" lane="3" entrytime="00:01:05.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="486" reactiontime="+82" swimtime="00:04:29.80" resultid="18188" heatid="19708" lane="6" entrytime="00:04:29.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.96" />
                    <SPLIT distance="100" swimtime="00:01:04.24" />
                    <SPLIT distance="150" swimtime="00:01:37.95" />
                    <SPLIT distance="200" swimtime="00:02:12.21" />
                    <SPLIT distance="250" swimtime="00:02:46.57" />
                    <SPLIT distance="300" swimtime="00:03:21.37" />
                    <SPLIT distance="350" swimtime="00:03:55.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-04-01" firstname="Piotr" gender="M" lastname="Konopacki" nation="POL" athleteid="18204">
              <RESULTS>
                <RESULT eventid="14189" points="378" reactiontime="+78" swimtime="00:10:12.92" resultid="18205" heatid="19617" lane="9" entrytime="00:10:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.66" />
                    <SPLIT distance="100" swimtime="00:01:09.66" />
                    <SPLIT distance="150" swimtime="00:01:48.04" />
                    <SPLIT distance="200" swimtime="00:02:27.39" />
                    <SPLIT distance="250" swimtime="00:03:07.03" />
                    <SPLIT distance="300" swimtime="00:03:46.35" />
                    <SPLIT distance="350" swimtime="00:04:25.77" />
                    <SPLIT distance="400" swimtime="00:05:05.07" />
                    <SPLIT distance="450" swimtime="00:05:44.47" />
                    <SPLIT distance="500" swimtime="00:06:23.35" />
                    <SPLIT distance="550" swimtime="00:07:02.41" />
                    <SPLIT distance="600" swimtime="00:07:41.13" />
                    <SPLIT distance="650" swimtime="00:08:20.32" />
                    <SPLIT distance="700" swimtime="00:08:59.00" />
                    <SPLIT distance="750" swimtime="00:09:37.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="312" swimtime="00:00:32.75" resultid="18206" heatid="19350" lane="8" entrytime="00:00:32.60" />
                <RESULT eventid="1273" points="378" reactiontime="+82" swimtime="00:01:02.15" resultid="18207" heatid="19384" lane="1" entrytime="00:01:01.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="376" reactiontime="+81" swimtime="00:02:17.59" resultid="18208" heatid="19485" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                    <SPLIT distance="100" swimtime="00:01:04.80" />
                    <SPLIT distance="150" swimtime="00:01:41.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="332" reactiontime="+67" swimtime="00:05:40.05" resultid="18209" heatid="19510" lane="0" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                    <SPLIT distance="100" swimtime="00:01:17.53" />
                    <SPLIT distance="150" swimtime="00:02:03.23" />
                    <SPLIT distance="200" swimtime="00:02:47.79" />
                    <SPLIT distance="250" swimtime="00:03:38.27" />
                    <SPLIT distance="300" swimtime="00:04:27.20" />
                    <SPLIT distance="350" swimtime="00:05:05.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="395" reactiontime="+75" swimtime="00:04:49.18" resultid="18210" heatid="19706" lane="5" entrytime="00:04:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                    <SPLIT distance="100" swimtime="00:01:07.53" />
                    <SPLIT distance="150" swimtime="00:01:44.90" />
                    <SPLIT distance="200" swimtime="00:02:23.37" />
                    <SPLIT distance="250" swimtime="00:03:01.01" />
                    <SPLIT distance="300" swimtime="00:03:38.49" />
                    <SPLIT distance="350" swimtime="00:04:15.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-06-13" firstname="Michał" gender="M" lastname="Kieres" nation="POL" athleteid="18123">
              <RESULTS>
                <RESULT eventid="1113" points="293" reactiontime="+76" swimtime="00:02:45.01" resultid="18124" heatid="19316" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                    <SPLIT distance="100" swimtime="00:01:18.77" />
                    <SPLIT distance="150" swimtime="00:02:05.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="319" reactiontime="+72" swimtime="00:02:56.09" resultid="18125" heatid="19364" lane="7" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                    <SPLIT distance="100" swimtime="00:01:22.71" />
                    <SPLIT distance="150" swimtime="00:02:09.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="297" reactiontime="+71" swimtime="00:02:42.60" resultid="18126" heatid="19417" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                    <SPLIT distance="100" swimtime="00:01:13.11" />
                    <SPLIT distance="150" swimtime="00:01:56.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="355" reactiontime="+68" swimtime="00:01:18.51" resultid="18127" heatid="19441" lane="8" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="303" reactiontime="+68" swimtime="00:05:50.38" resultid="18128" heatid="19511" lane="0" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="100" swimtime="00:01:16.64" />
                    <SPLIT distance="150" swimtime="00:02:05.00" />
                    <SPLIT distance="200" swimtime="00:02:52.78" />
                    <SPLIT distance="250" swimtime="00:03:41.05" />
                    <SPLIT distance="300" swimtime="00:04:30.14" />
                    <SPLIT distance="350" swimtime="00:05:10.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="18129" heatid="19523" lane="7" entrytime="00:01:08.00" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="18130" heatid="19557" lane="8" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-06-26" firstname="Monika" gender="F" lastname="Piwońska" nation="POL" athleteid="18158">
              <RESULTS>
                <RESULT eventid="1096" points="364" reactiontime="+86" swimtime="00:02:50.57" resultid="18159" heatid="19307" lane="5" entrytime="00:03:01.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                    <SPLIT distance="100" swimtime="00:01:18.12" />
                    <SPLIT distance="150" swimtime="00:02:08.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="18160" heatid="19336" lane="8" />
                <RESULT eventid="14225" points="394" reactiontime="+86" swimtime="00:01:17.25" resultid="18161" heatid="19394" lane="2" entrytime="00:01:17.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="433" reactiontime="+83" swimtime="00:00:32.22" resultid="18162" heatid="19448" lane="2" entrytime="00:00:33.33" />
                <RESULT eventid="1555" points="380" reactiontime="+85" swimtime="00:05:58.10" resultid="18163" heatid="19505" lane="8" entrytime="00:06:07.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.96" />
                    <SPLIT distance="100" swimtime="00:01:17.67" />
                    <SPLIT distance="150" swimtime="00:02:03.65" />
                    <SPLIT distance="200" swimtime="00:02:50.18" />
                    <SPLIT distance="250" swimtime="00:03:39.85" />
                    <SPLIT distance="300" swimtime="00:04:31.95" />
                    <SPLIT distance="350" swimtime="00:05:14.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-09-09" firstname="Marek" gender="M" lastname="Koźlikowski" nation="POL" athleteid="18115">
              <RESULTS>
                <RESULT eventid="14207" points="220" reactiontime="+98" swimtime="00:23:24.05" resultid="18116" heatid="19621" lane="9" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.88" />
                    <SPLIT distance="100" swimtime="00:01:29.29" />
                    <SPLIT distance="150" swimtime="00:02:15.89" />
                    <SPLIT distance="200" swimtime="00:03:03.16" />
                    <SPLIT distance="250" swimtime="00:03:50.44" />
                    <SPLIT distance="300" swimtime="00:04:37.90" />
                    <SPLIT distance="350" swimtime="00:05:25.76" />
                    <SPLIT distance="400" swimtime="00:06:13.55" />
                    <SPLIT distance="450" swimtime="00:07:00.79" />
                    <SPLIT distance="500" swimtime="00:07:48.18" />
                    <SPLIT distance="550" swimtime="00:08:35.02" />
                    <SPLIT distance="600" swimtime="00:09:22.17" />
                    <SPLIT distance="650" swimtime="00:10:09.21" />
                    <SPLIT distance="700" swimtime="00:10:55.93" />
                    <SPLIT distance="750" swimtime="00:11:43.27" />
                    <SPLIT distance="800" swimtime="00:12:30.11" />
                    <SPLIT distance="850" swimtime="00:13:17.22" />
                    <SPLIT distance="900" swimtime="00:14:04.22" />
                    <SPLIT distance="950" swimtime="00:14:51.15" />
                    <SPLIT distance="1000" swimtime="00:15:37.52" />
                    <SPLIT distance="1050" swimtime="00:16:23.82" />
                    <SPLIT distance="1100" swimtime="00:17:10.73" />
                    <SPLIT distance="1150" swimtime="00:17:57.52" />
                    <SPLIT distance="1200" swimtime="00:18:44.53" />
                    <SPLIT distance="1250" swimtime="00:19:31.78" />
                    <SPLIT distance="1300" swimtime="00:20:19.51" />
                    <SPLIT distance="1350" swimtime="00:21:06.91" />
                    <SPLIT distance="1400" swimtime="00:21:54.43" />
                    <SPLIT distance="1450" swimtime="00:22:41.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="229" reactiontime="+86" swimtime="00:03:16.85" resultid="18117" heatid="19361" lane="0" entrytime="00:03:30.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.09" />
                    <SPLIT distance="100" swimtime="00:01:35.30" />
                    <SPLIT distance="150" swimtime="00:02:26.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="230" reactiontime="+99" swimtime="00:01:22.00" resultid="18118" heatid="19399" lane="3" entrytime="00:01:37.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="228" reactiontime="+102" swimtime="00:01:30.97" resultid="18119" heatid="19435" lane="4" entrytime="00:01:44.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="199" reactiontime="+99" swimtime="00:06:42.72" resultid="18120" heatid="19508" lane="6" entrytime="00:07:00.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.12" />
                    <SPLIT distance="100" swimtime="00:01:39.54" />
                    <SPLIT distance="150" swimtime="00:02:34.70" />
                    <SPLIT distance="200" swimtime="00:03:29.22" />
                    <SPLIT distance="250" swimtime="00:04:22.49" />
                    <SPLIT distance="300" swimtime="00:05:15.66" />
                    <SPLIT distance="350" swimtime="00:06:00.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="156" reactiontime="+107" swimtime="00:01:29.18" resultid="18121" heatid="19518" lane="4" entrytime="00:01:34.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="222" reactiontime="+97" swimtime="00:05:50.50" resultid="18122" heatid="19702" lane="5" entrytime="00:06:03.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.95" />
                    <SPLIT distance="100" swimtime="00:01:24.94" />
                    <SPLIT distance="150" swimtime="00:02:10.35" />
                    <SPLIT distance="200" swimtime="00:02:55.59" />
                    <SPLIT distance="250" swimtime="00:03:41.11" />
                    <SPLIT distance="300" swimtime="00:04:26.28" />
                    <SPLIT distance="350" swimtime="00:05:10.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-17" firstname="Anna" gender="F" lastname="Zaleska" nation="POL" athleteid="18093">
              <RESULTS>
                <RESULT eventid="1096" status="WDR" swimtime="00:00:00.00" resultid="18094" entrytime="00:03:00.00" />
                <RESULT eventid="1147" status="WDR" swimtime="00:00:00.00" resultid="18095" entrytime="00:12:00.00" />
                <RESULT eventid="1187" status="WDR" swimtime="00:00:00.00" resultid="18096" entrytime="00:00:37.00" />
                <RESULT eventid="1324" status="WDR" swimtime="00:00:00.00" resultid="18097" entrytime="00:02:45.00" />
                <RESULT eventid="1423" status="WDR" swimtime="00:00:00.00" resultid="18098" entrytime="00:00:34.00" />
                <RESULT eventid="1491" status="WDR" swimtime="00:00:00.00" resultid="18099" entrytime="00:02:35.00" />
                <RESULT eventid="1595" status="WDR" swimtime="00:00:00.00" resultid="18100" entrytime="00:01:15.00" />
                <RESULT eventid="1721" status="WDR" swimtime="00:00:00.00" resultid="18101" entrytime="00:05:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-01-29" firstname="Mariusz" gender="M" lastname="Gabiec" nation="POL" athleteid="18211">
              <RESULTS>
                <RESULT eventid="1079" points="349" reactiontime="+88" swimtime="00:00:28.75" resultid="18212" heatid="19294" lane="2" entrytime="00:00:29.25" />
                <RESULT eventid="14189" points="355" reactiontime="+105" swimtime="00:10:25.66" resultid="18213" heatid="19617" lane="2" entrytime="00:10:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                    <SPLIT distance="100" swimtime="00:01:14.31" />
                    <SPLIT distance="150" swimtime="00:01:53.00" />
                    <SPLIT distance="200" swimtime="00:02:31.81" />
                    <SPLIT distance="250" swimtime="00:03:10.58" />
                    <SPLIT distance="300" swimtime="00:04:28.67" />
                    <SPLIT distance="350" swimtime="00:05:07.83" />
                    <SPLIT distance="400" swimtime="00:05:47.43" />
                    <SPLIT distance="450" swimtime="00:06:27.13" />
                    <SPLIT distance="500" swimtime="00:07:06.95" />
                    <SPLIT distance="550" swimtime="00:07:46.74" />
                    <SPLIT distance="600" swimtime="00:08:27.19" />
                    <SPLIT distance="650" swimtime="00:09:07.12" />
                    <SPLIT distance="700" swimtime="00:09:46.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="284" reactiontime="+83" swimtime="00:00:33.79" resultid="18214" heatid="19349" lane="9" entrytime="00:00:34.50" />
                <RESULT eventid="1341" points="273" reactiontime="+93" swimtime="00:02:47.24" resultid="18215" heatid="19415" lane="5" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.80" />
                    <SPLIT distance="100" swimtime="00:01:20.82" />
                    <SPLIT distance="150" swimtime="00:02:04.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="357" reactiontime="+94" swimtime="00:02:20.07" resultid="18216" heatid="19485" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                    <SPLIT distance="100" swimtime="00:01:08.65" />
                    <SPLIT distance="150" swimtime="00:01:44.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="275" reactiontime="+96" swimtime="00:06:01.92" resultid="18217" heatid="19509" lane="8" entrytime="00:06:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.25" />
                    <SPLIT distance="100" swimtime="00:01:24.32" />
                    <SPLIT distance="150" swimtime="00:02:57.11" />
                    <SPLIT distance="250" swimtime="00:03:51.23" />
                    <SPLIT distance="300" swimtime="00:04:44.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="312" reactiontime="+93" swimtime="00:01:10.84" resultid="18218" heatid="19520" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="339" reactiontime="+100" swimtime="00:05:04.33" resultid="18219" heatid="19706" lane="3" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                    <SPLIT distance="100" swimtime="00:01:13.87" />
                    <SPLIT distance="150" swimtime="00:01:52.67" />
                    <SPLIT distance="200" swimtime="00:02:31.30" />
                    <SPLIT distance="250" swimtime="00:03:09.71" />
                    <SPLIT distance="300" swimtime="00:03:48.54" />
                    <SPLIT distance="350" swimtime="00:04:27.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-08-16" firstname="Paweł" gender="M" lastname="Szczuka" nation="POL" athleteid="18164">
              <RESULTS>
                <RESULT eventid="1113" points="443" reactiontime="+87" swimtime="00:02:23.78" resultid="18165" heatid="19317" lane="0" entrytime="00:02:28.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                    <SPLIT distance="100" swimtime="00:01:07.54" />
                    <SPLIT distance="150" swimtime="00:01:49.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="18166" heatid="19351" lane="3" entrytime="00:00:30.80" />
                <RESULT eventid="14243" points="472" reactiontime="+84" swimtime="00:01:04.57" resultid="18167" heatid="19408" lane="3" entrytime="00:01:05.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="454" reactiontime="+91" swimtime="00:05:06.38" resultid="18168" heatid="19512" lane="1" entrytime="00:05:11.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                    <SPLIT distance="100" swimtime="00:01:07.48" />
                    <SPLIT distance="150" swimtime="00:01:46.51" />
                    <SPLIT distance="200" swimtime="00:02:27.45" />
                    <SPLIT distance="250" swimtime="00:03:09.93" />
                    <SPLIT distance="300" swimtime="00:03:54.76" />
                    <SPLIT distance="350" swimtime="00:04:30.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-09-29" firstname="Jakub" gender="M" lastname="Stępień" nation="POL" athleteid="18151">
              <RESULTS>
                <RESULT eventid="1079" points="338" reactiontime="+85" swimtime="00:00:29.08" resultid="18152" heatid="19296" lane="5" entrytime="00:00:28.49" />
                <RESULT eventid="14189" reactiontime="+95" status="OTL" swimtime="00:11:15.35" resultid="18153" heatid="19616" lane="3" entrytime="00:10:57.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                    <SPLIT distance="100" swimtime="00:01:14.36" />
                    <SPLIT distance="150" swimtime="00:01:54.62" />
                    <SPLIT distance="200" swimtime="00:02:35.61" />
                    <SPLIT distance="250" swimtime="00:03:17.67" />
                    <SPLIT distance="300" swimtime="00:04:00.13" />
                    <SPLIT distance="350" swimtime="00:04:42.96" />
                    <SPLIT distance="400" swimtime="00:05:26.26" />
                    <SPLIT distance="450" swimtime="00:06:10.50" />
                    <SPLIT distance="500" swimtime="00:06:53.37" />
                    <SPLIT distance="550" swimtime="00:07:37.05" />
                    <SPLIT distance="600" swimtime="00:08:20.70" />
                    <SPLIT distance="650" swimtime="00:09:05.11" />
                    <SPLIT distance="700" swimtime="00:09:50.02" />
                    <SPLIT distance="750" swimtime="00:10:33.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="18154" heatid="19342" lane="2" />
                <RESULT eventid="1273" points="350" reactiontime="+88" swimtime="00:01:03.76" resultid="18155" heatid="19383" lane="1" entrytime="00:01:02.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="255" reactiontime="+90" swimtime="00:00:34.37" resultid="18156" heatid="19450" lane="2" />
                <RESULT eventid="1508" points="333" reactiontime="+93" swimtime="00:02:23.25" resultid="18157" heatid="19493" lane="6" entrytime="00:02:17.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                    <SPLIT distance="100" swimtime="00:01:08.16" />
                    <SPLIT distance="150" swimtime="00:01:45.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-10-26" firstname="Joanna" gender="F" lastname="Drzewicka" nation="POL" athleteid="18088">
              <RESULTS>
                <RESULT eventid="1062" points="256" reactiontime="+99" swimtime="00:00:36.60" resultid="18089" heatid="19278" lane="3" entrytime="00:00:38.00" />
                <RESULT eventid="1187" points="275" reactiontime="+80" swimtime="00:00:39.47" resultid="18090" heatid="19339" lane="9" entrytime="00:00:41.00" />
                <RESULT eventid="14225" points="183" reactiontime="+97" swimtime="00:01:39.72" resultid="18091" heatid="19391" lane="5" entrytime="00:01:34.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="232" reactiontime="+72" swimtime="00:01:29.45" resultid="18092" heatid="19467" lane="9" entrytime="00:01:31.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-09-15" firstname="Adam" gender="M" lastname="Szmit" nation="POL" athleteid="18110">
              <RESULTS>
                <RESULT eventid="14207" points="252" reactiontime="+112" swimtime="00:22:21.02" resultid="18111" heatid="19622" lane="8" entrytime="00:22:30.00" />
                <RESULT eventid="1273" points="237" reactiontime="+112" swimtime="00:01:12.56" resultid="18112" heatid="19379" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="232" reactiontime="+104" swimtime="00:02:41.56" resultid="18113" heatid="19491" lane="9" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                    <SPLIT distance="150" swimtime="00:02:00.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="244" swimtime="00:05:39.29" resultid="18114" heatid="19704" lane="0" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.07" />
                    <SPLIT distance="200" swimtime="00:02:45.53" />
                    <SPLIT distance="250" swimtime="00:03:28.79" />
                    <SPLIT distance="300" swimtime="00:04:13.10" />
                    <SPLIT distance="350" swimtime="00:04:57.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-03-10" firstname="Katarzyna" gender="F" lastname="Sienkiewicz" nation="POL" athleteid="18143">
              <RESULTS>
                <RESULT eventid="1062" points="214" reactiontime="+97" swimtime="00:00:38.84" resultid="18144" heatid="19275" lane="8" />
                <RESULT eventid="1187" points="126" reactiontime="+82" swimtime="00:00:51.08" resultid="18145" heatid="19336" lane="7" />
                <RESULT eventid="1256" points="174" reactiontime="+91" swimtime="00:01:31.08" resultid="18146" heatid="19366" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="168" reactiontime="+94" swimtime="00:01:52.93" resultid="18147" heatid="19426" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="109" reactiontime="+79" swimtime="00:01:54.88" resultid="18148" heatid="19465" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" status="DNS" swimtime="00:00:00.00" resultid="18149" heatid="19526" lane="8" />
                <RESULT comment="K14 - Praca nóg w płaszczyźnie pionowej w dół (z wyjątkiem jednego ruchu po starcie i nawrocie) (Time: 10:40)" eventid="1664" reactiontime="+93" status="DSQ" swimtime="00:00:49.38" resultid="18150" heatid="19538" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="407" reactiontime="+69" swimtime="00:02:02.11" resultid="18230" heatid="19423" lane="4" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                    <SPLIT distance="100" swimtime="00:01:04.78" />
                    <SPLIT distance="150" swimtime="00:01:33.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18204" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="18164" number="2" reactiontime="+45" />
                    <RELAYPOSITION athleteid="18180" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="18151" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="228" reactiontime="+78" swimtime="00:02:28.15" resultid="18232" heatid="19422" lane="1" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.04" />
                    <SPLIT distance="100" swimtime="00:01:12.48" />
                    <SPLIT distance="150" swimtime="00:01:55.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18173" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="18123" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="18189" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="18110" number="4" reactiontime="+52" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="265" reactiontime="+87" swimtime="00:02:20.87" resultid="18234" heatid="19422" lane="6" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                    <SPLIT distance="100" swimtime="00:01:12.42" />
                    <SPLIT distance="150" swimtime="00:01:49.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18211" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="18137" number="2" reactiontime="+43" />
                    <RELAYPOSITION athleteid="18220" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="18115" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1548" status="DNS" swimtime="00:00:00.00" resultid="18231" heatid="19502" lane="1" entrytime="00:01:49.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18180" number="1" />
                    <RELAYPOSITION athleteid="18151" number="2" />
                    <RELAYPOSITION athleteid="18204" number="3" />
                    <RELAYPOSITION athleteid="18164" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1548" status="DNS" swimtime="00:00:00.00" resultid="18233" heatid="19500" lane="1" entrytime="00:02:09.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18123" number="1" />
                    <RELAYPOSITION athleteid="18110" number="2" />
                    <RELAYPOSITION athleteid="18189" number="3" />
                    <RELAYPOSITION athleteid="18220" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1548" points="285" reactiontime="+87" swimtime="00:02:05.46" resultid="18235" heatid="19500" lane="3" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                    <SPLIT distance="100" swimtime="00:01:00.38" />
                    <SPLIT distance="150" swimtime="00:01:32.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18173" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="18137" number="2" reactiontime="+21" />
                    <RELAYPOSITION athleteid="18115" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="18211" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1358" points="251" reactiontime="+73" swimtime="00:02:43.63" resultid="18228" heatid="19420" lane="7" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.96" />
                    <SPLIT distance="150" swimtime="00:02:04.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18088" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="18102" number="2" />
                    <RELAYPOSITION athleteid="18131" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="18143" number="4" reactiontime="+52" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1525" points="286" reactiontime="+83" swimtime="00:02:22.99" resultid="18229" heatid="19498" lane="8" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                    <SPLIT distance="100" swimtime="00:01:08.98" />
                    <SPLIT distance="150" swimtime="00:01:55.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18131" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="18088" number="2" reactiontime="+19" />
                    <RELAYPOSITION athleteid="18143" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="18102" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="304" reactiontime="+71" swimtime="00:02:11.70" resultid="18225" heatid="19321" lane="0" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.26" />
                    <SPLIT distance="100" swimtime="00:01:03.93" />
                    <SPLIT distance="150" swimtime="00:01:42.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18204" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="18088" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="18143" number="3" reactiontime="+17" />
                    <RELAYPOSITION athleteid="18173" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1698" points="340" reactiontime="+76" swimtime="00:02:19.20" resultid="18227" heatid="19563" lane="6" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.34" />
                    <SPLIT distance="100" swimtime="00:01:16.38" />
                    <SPLIT distance="150" swimtime="00:01:46.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18088" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="18123" number="2" reactiontime="+24" />
                    <RELAYPOSITION athleteid="18180" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="18131" number="4" reactiontime="+70" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1698" status="DNS" swimtime="00:00:00.00" resultid="18224" heatid="19561" lane="4" entrytime="00:02:26.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18204" number="1" />
                    <RELAYPOSITION athleteid="18102" number="2" />
                    <RELAYPOSITION athleteid="18211" number="3" />
                    <RELAYPOSITION athleteid="18143" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1130" points="389" reactiontime="+73" swimtime="00:02:01.30" resultid="18226" heatid="19321" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.49" />
                    <SPLIT distance="100" swimtime="00:00:59.65" />
                    <SPLIT distance="150" swimtime="00:01:34.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18164" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="18131" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="18102" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="18180" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="AQUNI" nation="SVK" region="ZSO" clubid="16098" name="AQUATICS Nitra">
          <ATHLETES>
            <ATHLETE birthdate="1970-02-03" firstname="Peter" gender="M" lastname="Čigáš" nation="SVK" license="SVK15844" athleteid="16982">
              <RESULTS>
                <RESULT eventid="1079" status="WDR" swimtime="00:00:00.00" resultid="16983" entrytime="00:00:27.22" entrycourse="SCM" />
                <RESULT eventid="1205" status="WDR" swimtime="00:00:00.00" resultid="16984" entrytime="00:00:30.18" entrycourse="SCM" />
                <RESULT eventid="1273" status="WDR" swimtime="00:00:00.00" resultid="16985" entrytime="00:00:59.71" entrycourse="SCM" />
                <RESULT eventid="1474" status="WDR" swimtime="00:00:00.00" resultid="16986" entrytime="00:01:04.96" entrycourse="SCM" />
                <RESULT eventid="1647" status="WDR" swimtime="00:00:00.00" resultid="16987" entrytime="00:02:23.22" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-06-08" firstname="Miroslav" gender="M" lastname="Ábel" nation="SVK" license="SVK12721" athleteid="16969" firstname.en="Abel" lastname.en="Miroslav">
              <RESULTS>
                <RESULT eventid="1113" points="489" reactiontime="+73" swimtime="00:02:19.07" resultid="16970" heatid="19318" lane="9" entrytime="00:02:20.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.88" />
                    <SPLIT distance="100" swimtime="00:01:04.99" />
                    <SPLIT distance="150" swimtime="00:01:45.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="408" reactiontime="+84" swimtime="00:02:26.28" resultid="16971" heatid="19418" lane="2" entrytime="00:02:21.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                    <SPLIT distance="100" swimtime="00:01:08.53" />
                    <SPLIT distance="150" swimtime="00:01:46.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="436" reactiontime="+85" swimtime="00:02:10.99" resultid="16972" heatid="19494" lane="5" entrytime="00:02:10.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.13" />
                    <SPLIT distance="100" swimtime="00:01:02.73" />
                    <SPLIT distance="150" swimtime="00:01:37.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="475" reactiontime="+77" swimtime="00:01:01.61" resultid="16973" heatid="19525" lane="7" entrytime="00:00:59.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="404" reactiontime="+82" swimtime="00:04:46.89" resultid="16974" heatid="19707" lane="0" entrytime="00:04:49.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                    <SPLIT distance="100" swimtime="00:01:09.36" />
                    <SPLIT distance="150" swimtime="00:01:46.69" />
                    <SPLIT distance="200" swimtime="00:02:23.63" />
                    <SPLIT distance="250" swimtime="00:03:00.51" />
                    <SPLIT distance="300" swimtime="00:03:36.36" />
                    <SPLIT distance="350" swimtime="00:04:12.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-05-08" firstname="Karol" gender="M" lastname="Lacko" nation="SVK" license="SVK16793" athleteid="16994">
              <RESULTS>
                <RESULT eventid="14207" points="337" reactiontime="+97" swimtime="00:20:18.48" resultid="16995" heatid="19623" lane="9" entrytime="00:20:55.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.50" />
                    <SPLIT distance="100" swimtime="00:01:17.66" />
                    <SPLIT distance="150" swimtime="00:01:58.07" />
                    <SPLIT distance="200" swimtime="00:02:38.67" />
                    <SPLIT distance="250" swimtime="00:03:18.85" />
                    <SPLIT distance="300" swimtime="00:03:59.01" />
                    <SPLIT distance="350" swimtime="00:04:39.20" />
                    <SPLIT distance="400" swimtime="00:05:19.25" />
                    <SPLIT distance="450" swimtime="00:05:59.48" />
                    <SPLIT distance="500" swimtime="00:06:39.94" />
                    <SPLIT distance="550" swimtime="00:07:20.66" />
                    <SPLIT distance="600" swimtime="00:08:01.07" />
                    <SPLIT distance="650" swimtime="00:08:41.46" />
                    <SPLIT distance="700" swimtime="00:09:22.09" />
                    <SPLIT distance="750" swimtime="00:10:02.48" />
                    <SPLIT distance="800" swimtime="00:10:42.79" />
                    <SPLIT distance="850" swimtime="00:11:23.48" />
                    <SPLIT distance="900" swimtime="00:12:03.90" />
                    <SPLIT distance="950" swimtime="00:12:44.66" />
                    <SPLIT distance="1000" swimtime="00:13:25.76" />
                    <SPLIT distance="1050" swimtime="00:14:06.98" />
                    <SPLIT distance="1100" swimtime="00:14:48.34" />
                    <SPLIT distance="1150" swimtime="00:15:29.47" />
                    <SPLIT distance="1200" swimtime="00:16:11.45" />
                    <SPLIT distance="1250" swimtime="00:16:53.19" />
                    <SPLIT distance="1300" swimtime="00:17:34.85" />
                    <SPLIT distance="1350" swimtime="00:18:16.25" />
                    <SPLIT distance="1400" swimtime="00:18:57.76" />
                    <SPLIT distance="1450" swimtime="00:19:38.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="384" reactiontime="+87" swimtime="00:02:16.66" resultid="16996" heatid="19494" lane="1" entrytime="00:02:13.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                    <SPLIT distance="100" swimtime="00:01:06.37" />
                    <SPLIT distance="150" swimtime="00:01:41.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="365" reactiontime="+90" swimtime="00:04:56.80" resultid="16997" heatid="19707" lane="1" entrytime="00:04:45.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                    <SPLIT distance="100" swimtime="00:01:12.54" />
                    <SPLIT distance="200" swimtime="00:02:27.48" />
                    <SPLIT distance="250" swimtime="00:03:05.57" />
                    <SPLIT distance="300" swimtime="00:03:42.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-09-12" firstname="Peter" gender="M" lastname="Korobov" nation="SVK" license="SVK16881" athleteid="16988">
              <RESULTS>
                <RESULT eventid="1079" status="WDR" swimtime="00:00:00.00" resultid="16989" entrytime="00:00:27.52" entrycourse="SCM" />
                <RESULT eventid="1205" status="WDR" swimtime="00:00:00.00" resultid="16990" entrytime="00:00:33.12" entrycourse="SCM" />
                <RESULT eventid="1273" status="WDR" swimtime="00:00:00.00" resultid="16991" entrytime="00:01:00.76" entrycourse="SCM" />
                <RESULT eventid="1440" status="WDR" swimtime="00:00:00.00" resultid="16992" entrytime="00:00:32.28" entrycourse="SCM" />
                <RESULT eventid="1681" status="WDR" swimtime="00:00:00.00" resultid="16993" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-04-01" firstname="Lucia" gender="F" lastname="Ábelová" nation="SVK" license="SVK19294" athleteid="16975">
              <RESULTS>
                <RESULT eventid="1062" points="185" reactiontime="+96" swimtime="00:00:40.74" resultid="16976" heatid="19277" lane="8" entrytime="00:00:43.78" entrycourse="SCM" />
                <RESULT eventid="1187" points="133" swimtime="00:00:50.23" resultid="16977" heatid="19337" lane="7" entrytime="00:00:52.67" entrycourse="SCM" />
                <RESULT eventid="14225" points="134" reactiontime="+107" swimtime="00:01:50.57" resultid="16978" heatid="19390" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.77" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K16 - Niejednoczesne dotknięcie ściany dłońmi przy nawrocie lub na zakończenie wyścigu (Time: 16:18)" eventid="1388" reactiontime="+101" status="DSQ" swimtime="00:01:42.46" resultid="16979" heatid="19428" lane="4" entrytime="00:01:48.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="233" reactiontime="+90" swimtime="00:00:46.51" resultid="16980" heatid="19541" lane="7" entrytime="00:00:46.09" entrycourse="SCM" />
                <RESULT eventid="1491" points="118" reactiontime="+101" swimtime="00:03:45.64" resultid="16981" heatid="19480" lane="2" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.50" />
                    <SPLIT distance="100" swimtime="00:01:48.13" />
                    <SPLIT distance="150" swimtime="00:02:49.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" status="DNS" swimtime="00:00:00.00" resultid="18541" heatid="19499" lane="8">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16982" number="1" />
                    <RELAYPOSITION athleteid="16994" number="2" />
                    <RELAYPOSITION athleteid="16988" number="3" />
                    <RELAYPOSITION athleteid="16969" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" status="DNS" swimtime="00:00:00.00" resultid="18542" heatid="19421" lane="8">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16982" number="1" />
                    <RELAYPOSITION athleteid="16969" number="2" />
                    <RELAYPOSITION athleteid="16988" number="3" />
                    <RELAYPOSITION athleteid="16994" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00611" nation="POL" region="SLA" clubid="16681" name="AZS AWF Katowice">
          <CONTACT city="Katowice" email="m.skora@awf.katowice.pl" name="Michał Skóra" phone="501 370 222" state="ŚLĄSK" street="Mikołowska 72a" zip="40-065" />
          <ATHLETES>
            <ATHLETE birthdate="1986-12-21" firstname="Marcin" gender="M" lastname="Unold" nation="POL" athleteid="16682">
              <RESULTS>
                <RESULT eventid="1079" points="600" reactiontime="+77" swimtime="00:00:24.02" resultid="16683" heatid="19304" lane="2" entrytime="00:00:23.80" />
                <RESULT eventid="1205" points="588" reactiontime="+75" swimtime="00:00:26.52" resultid="16684" heatid="19353" lane="6" entrytime="00:00:27.00" />
                <RESULT eventid="1273" points="663" reactiontime="+77" swimtime="00:00:51.53" resultid="16685" heatid="19388" lane="5" entrytime="00:00:52.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZS WSB" nation="POL" region="SLA" clubid="14982" name="AZS WSB Dąbrowa Górnicza">
          <CONTACT city="Dąbrowa Górnicza" email="msadowski@wsb.edu.pl" internet="azs.wsb.edu.pl" name="Sadowski Maciej" state="ŚLĄSK" street="Cieplaka 1C" zip="41-300" />
          <ATHLETES>
            <ATHLETE birthdate="1996-05-27" firstname="Monika" gender="F" lastname="Kisiel" nation="POL" athleteid="14983">
              <RESULTS>
                <RESULT eventid="1147" points="386" reactiontime="+86" swimtime="00:10:58.16" resultid="14984" heatid="19596" lane="5" entrytime="00:10:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.51" />
                    <SPLIT distance="100" swimtime="00:01:12.39" />
                    <SPLIT distance="150" swimtime="00:01:51.36" />
                    <SPLIT distance="200" swimtime="00:02:31.79" />
                    <SPLIT distance="250" swimtime="00:03:13.37" />
                    <SPLIT distance="300" swimtime="00:03:55.30" />
                    <SPLIT distance="350" swimtime="00:04:37.96" />
                    <SPLIT distance="400" swimtime="00:05:21.02" />
                    <SPLIT distance="450" swimtime="00:06:03.36" />
                    <SPLIT distance="500" swimtime="00:06:46.43" />
                    <SPLIT distance="550" swimtime="00:07:29.47" />
                    <SPLIT distance="600" swimtime="00:08:11.59" />
                    <SPLIT distance="650" swimtime="00:08:53.56" />
                    <SPLIT distance="700" swimtime="00:09:36.05" />
                    <SPLIT distance="750" swimtime="00:10:18.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="480" reactiontime="+73" swimtime="00:01:10.24" resultid="14985" heatid="19469" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZS PWSZ R" nation="POL" region="SLA" clubid="14725" name="AZSPWSZ Raciborz" shortname="Akademicki Związek Sportowy Pa">
          <CONTACT city="Raciborz" email="adip45@poczta.onet.pl" name="Kunicki" state="ŚL" street="Słowackiego 55" zip="47-400" />
          <ATHLETES>
            <ATHLETE birthdate="1957-04-11" firstname="Adolf" gender="M" lastname="Piechula" nation="POL" athleteid="14726">
              <RESULTS>
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="14727" heatid="19310" lane="9" entrytime="00:03:07.34" entrycourse="SCM" />
                <RESULT eventid="1239" points="227" reactiontime="+90" swimtime="00:03:17.23" resultid="14728" heatid="19361" lane="6" entrytime="00:03:23.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.43" />
                    <SPLIT distance="100" swimtime="00:01:34.68" />
                    <SPLIT distance="150" swimtime="00:02:26.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="177" reactiontime="+97" swimtime="00:03:13.04" resultid="14729" heatid="19415" lane="6" entrytime="00:03:15.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.96" />
                    <SPLIT distance="100" swimtime="00:01:31.34" />
                    <SPLIT distance="150" swimtime="00:02:22.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="250" reactiontime="+86" swimtime="00:01:28.24" resultid="14730" heatid="19437" lane="2" entrytime="00:01:29.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="205" reactiontime="+95" swimtime="00:06:39.01" resultid="14731" heatid="19508" lane="4" entrytime="00:06:42.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.92" />
                    <SPLIT distance="100" swimtime="00:01:33.36" />
                    <SPLIT distance="150" swimtime="00:02:24.89" />
                    <SPLIT distance="200" swimtime="00:03:16.20" />
                    <SPLIT distance="250" swimtime="00:04:13.45" />
                    <SPLIT distance="300" swimtime="00:05:08.71" />
                    <SPLIT distance="350" swimtime="00:05:56.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="179" reactiontime="+93" swimtime="00:01:25.23" resultid="14732" heatid="19519" lane="3" entrytime="00:01:25.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="273" reactiontime="+83" swimtime="00:00:38.89" resultid="14733" heatid="19552" lane="9" entrytime="00:00:39.50" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CMUJKR" nation="POL" region="MAL" clubid="15985" name="Collegium Medicum UJ Masters Kraków" shortname="Collegium Medicum UJ Masters K">
          <CONTACT city="Kraków" email="mariuszbaranik@gmail.com" name="Mariusz Baranik" phone="698128222" state="MAL" street="Białopradnicka 32c/3" zip="31-221" />
          <ATHLETES>
            <ATHLETE birthdate="1969-08-22" firstname="Mirosław" gender="M" lastname="Woźniak" nation="POL" athleteid="15986">
              <RESULTS>
                <RESULT eventid="1079" points="351" reactiontime="+82" swimtime="00:00:28.72" resultid="15987" heatid="19297" lane="7" entrytime="00:00:28.00" />
                <RESULT eventid="1113" points="294" reactiontime="+91" swimtime="00:02:44.81" resultid="15988" heatid="19313" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                    <SPLIT distance="100" swimtime="00:01:18.05" />
                    <SPLIT distance="150" swimtime="00:02:06.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="UKR" clubid="17570" name="Crazy Fish">
          <CONTACT city="Poltava" email="maksym.yakovenko@skazhenikarasi.com.ua" fax="+380 50 131 1623" internet="www.skazhenikarasi.com.ua" name="Yakovenko Maksym" phone="+380 97 643 6156" />
          <ATHLETES>
            <ATHLETE birthdate="1957-05-11" firstname="Mykola" gender="M" lastname="Klymko" nation="UKR" athleteid="17571">
              <RESULTS>
                <RESULT eventid="1079" points="338" reactiontime="+88" swimtime="00:00:29.08" resultid="17572" heatid="19294" lane="7" entrytime="00:00:29.32" />
                <RESULT eventid="1205" points="238" reactiontime="+81" swimtime="00:00:35.83" resultid="17573" heatid="19347" lane="2" entrytime="00:00:37.18" />
                <RESULT eventid="1440" points="317" reactiontime="+95" swimtime="00:00:31.94" resultid="17574" heatid="19456" lane="1" entrytime="00:00:32.64" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="UKR" clubid="17575" name="Euro-Lviv MSC">
          <CONTACT city="Lviv" email="madam57@ukr.net, riff.lviv@gmail.com" fax="+38 067 673 4796" internet="www.mastersswim.com.ua" name="Khiresh Lyudmyla" phone="+38 067 371 2151" zip="79000" />
          <ATHLETES>
            <ATHLETE birthdate="1976-02-03" firstname="Romana" gender="F" lastname="Sirenko" nation="UKR" athleteid="17631">
              <RESULTS>
                <RESULT eventid="1096" status="DNS" swimtime="00:00:00.00" resultid="17632" heatid="19307" lane="8" entrytime="00:03:07.50" />
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="17633" heatid="19339" lane="6" entrytime="00:00:38.50" />
                <RESULT eventid="14225" status="DNS" swimtime="00:00:00.00" resultid="17634" heatid="19393" lane="6" entrytime="00:01:24.00" />
                <RESULT eventid="1423" status="DNS" swimtime="00:00:00.00" resultid="17635" heatid="19447" lane="8" entrytime="00:00:37.00" />
                <RESULT eventid="1457" status="DNS" swimtime="00:00:00.00" resultid="17636" heatid="19467" lane="6" entrytime="00:01:25.50" />
                <RESULT eventid="1595" status="DNS" swimtime="00:00:00.00" resultid="17637" heatid="19514" lane="1" entrytime="00:01:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-01-07" firstname="Ruslan" gender="M" lastname="Friauf" nation="UKR" athleteid="17648">
              <RESULTS>
                <RESULT eventid="1113" points="202" reactiontime="+82" swimtime="00:03:06.58" resultid="17649" heatid="19312" lane="7" entrytime="00:03:05.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.90" />
                    <SPLIT distance="100" swimtime="00:01:27.93" />
                    <SPLIT distance="150" swimtime="00:02:22.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="193" swimtime="00:00:38.43" resultid="17650" heatid="19347" lane="8" entrytime="00:00:38.56" />
                <RESULT eventid="14243" points="255" reactiontime="+88" swimtime="00:01:19.29" resultid="17651" heatid="19401" lane="3" entrytime="00:01:22.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="174" reactiontime="+78" swimtime="00:01:27.58" resultid="17652" heatid="19474" lane="9" entrytime="00:01:26.33" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-06-23" firstname="Nadiya" gender="F" lastname="Sannikova" nation="UKR" athleteid="17604">
              <RESULTS>
                <RESULT eventid="1222" points="162" swimtime="00:04:06.70" resultid="17605" heatid="19356" lane="0" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.31" />
                    <SPLIT distance="100" swimtime="00:01:56.45" />
                    <SPLIT distance="150" swimtime="00:03:02.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="195" reactiontime="+101" swimtime="00:00:49.35" resultid="17606" heatid="19540" lane="5" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-02-05" firstname="Lyudmyla" gender="F" lastname="Khiresh" nation="UKR" athleteid="17627">
              <RESULTS>
                <RESULT eventid="1062" points="239" reactiontime="+89" swimtime="00:00:37.40" resultid="17628" heatid="19279" lane="8" entrytime="00:00:36.00" />
                <RESULT eventid="14225" points="252" reactiontime="+101" swimtime="00:01:29.67" resultid="17629" heatid="19392" lane="3" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="237" swimtime="00:01:28.90" resultid="17630" heatid="19467" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-18" firstname="Dmytro" gender="M" lastname="Melnyk" nation="UKR" athleteid="17585">
              <RESULTS>
                <RESULT eventid="1079" points="487" reactiontime="+78" swimtime="00:00:25.74" resultid="17586" heatid="19300" lane="2" entrytime="00:00:26.25" />
                <RESULT eventid="1273" points="491" reactiontime="+70" swimtime="00:00:56.95" resultid="17587" heatid="19385" lane="7" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="450" reactiontime="+76" swimtime="00:01:12.54" resultid="17588" heatid="19441" lane="0" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="490" reactiontime="+71" swimtime="00:00:32.02" resultid="17589" heatid="19558" lane="0" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-11-30" firstname="Tetiana" gender="F" lastname="Kozakova" nation="UKR" athleteid="17638">
              <RESULTS>
                <RESULT eventid="1062" points="105" reactiontime="+108" swimtime="00:00:49.18" resultid="17639" heatid="19276" lane="5" entrytime="00:00:48.00" />
                <RESULT eventid="1187" points="99" reactiontime="+89" swimtime="00:00:55.46" resultid="17640" heatid="19337" lane="8" entrytime="00:00:54.00" />
                <RESULT eventid="14225" points="106" reactiontime="+104" swimtime="00:01:59.64" resultid="17641" heatid="19391" lane="9" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="80" reactiontime="+122" swimtime="00:00:56.44" resultid="17642" heatid="19445" lane="0" entrytime="00:00:58.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-07-31" firstname="Roman" gender="M" lastname="Koretskyy" nation="UKR" athleteid="17601">
              <RESULTS>
                <RESULT eventid="1079" points="126" reactiontime="+114" swimtime="00:00:40.33" resultid="17602" heatid="19286" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="1273" points="106" reactiontime="+90" swimtime="00:01:34.67" resultid="17603" heatid="19377" lane="9" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-10-31" firstname="Dmytro" gender="M" lastname="Ishchenko" nation="UKR" athleteid="17622">
              <RESULTS>
                <RESULT eventid="1079" points="333" reactiontime="+78" swimtime="00:00:29.21" resultid="17623" heatid="19296" lane="8" entrytime="00:00:28.90" />
                <RESULT eventid="1273" points="345" reactiontime="+86" swimtime="00:01:04.06" resultid="17624" heatid="19382" lane="7" entrytime="00:01:04.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="312" reactiontime="+91" swimtime="00:00:32.13" resultid="17625" heatid="19458" lane="4" entrytime="00:00:30.90" />
                <RESULT eventid="1613" points="262" reactiontime="+79" swimtime="00:01:15.08" resultid="17626" heatid="19521" lane="0" entrytime="00:01:14.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-05-24" firstname="Larysa" gender="F" lastname="Tsovkh" nation="UKR" athleteid="17618">
              <RESULTS>
                <RESULT eventid="1062" points="182" reactiontime="+92" swimtime="00:00:40.98" resultid="17619" heatid="19277" lane="6" entrytime="00:00:42.00" />
                <RESULT eventid="1388" points="200" reactiontime="+89" swimtime="00:01:46.59" resultid="17620" heatid="19429" lane="8" entrytime="00:01:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" status="DNS" swimtime="00:00:00.00" resultid="17621" heatid="19541" lane="8" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-06-24" firstname="Inna" gender="F" lastname="Hordii" nation="UKR" athleteid="17595">
              <RESULTS>
                <RESULT eventid="1062" points="371" swimtime="00:00:32.34" resultid="17596" heatid="19282" lane="0" entrytime="00:00:31.50" />
                <RESULT eventid="1187" points="285" reactiontime="+80" swimtime="00:00:39.00" resultid="17597" heatid="19339" lane="1" entrytime="00:00:39.00" />
                <RESULT eventid="14225" points="316" reactiontime="+89" swimtime="00:01:23.15" resultid="17598" heatid="19393" lane="4" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="323" reactiontime="+88" swimtime="00:00:35.50" resultid="17599" heatid="19447" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="1595" points="294" reactiontime="+97" swimtime="00:01:22.05" resultid="17600" heatid="19514" lane="4" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-05-19" firstname="Maryna" gender="F" lastname="Marchuk" nation="UKR" athleteid="17643">
              <RESULTS>
                <RESULT eventid="1062" points="403" swimtime="00:00:31.45" resultid="17644" heatid="19282" lane="9" entrytime="00:00:31.50" />
                <RESULT eventid="14225" status="DNS" swimtime="00:00:00.00" resultid="17645" heatid="19393" lane="1" entrytime="00:01:25.00" />
                <RESULT eventid="1388" points="280" reactiontime="+78" swimtime="00:01:35.25" resultid="17646" heatid="19430" lane="2" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="307" reactiontime="+76" swimtime="00:00:42.43" resultid="17647" heatid="19545" lane="9" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-09-13" firstname="Oleksandr" gender="M" lastname="Syrbu" nation="UKR" athleteid="17607">
              <RESULTS>
                <RESULT eventid="1079" points="478" reactiontime="+74" swimtime="00:00:25.91" resultid="17608" heatid="19302" lane="9" entrytime="00:00:25.92" />
                <RESULT eventid="1273" points="466" reactiontime="+80" swimtime="00:00:57.94" resultid="17609" heatid="19386" lane="3" entrytime="00:00:57.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="387" reactiontime="+84" swimtime="00:02:28.93" resultid="17610" heatid="19418" lane="0" entrytime="00:02:29.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.48" />
                    <SPLIT distance="100" swimtime="00:01:13.30" />
                    <SPLIT distance="150" swimtime="00:01:51.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="523" reactiontime="+73" swimtime="00:00:27.05" resultid="17611" heatid="19463" lane="9" entrytime="00:00:27.12" />
                <RESULT eventid="1613" points="422" reactiontime="+80" swimtime="00:01:04.08" resultid="17612" heatid="19524" lane="0" entrytime="00:01:04.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-11" firstname="Oleksandr" gender="M" lastname="Rekunkov" nation="UKR" athleteid="18519">
              <RESULTS>
                <RESULT eventid="1079" points="151" reactiontime="+106" swimtime="00:00:38.04" resultid="18520" heatid="19287" lane="8" entrytime="00:00:38.00" />
                <RESULT eventid="1205" points="115" reactiontime="+95" swimtime="00:00:45.65" resultid="18521" heatid="19345" lane="3" entrytime="00:00:43.00" />
                <RESULT eventid="1273" points="144" reactiontime="+128" swimtime="00:01:25.63" resultid="18522" heatid="19376" lane="1" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="155" reactiontime="+105" swimtime="00:01:43.38" resultid="18523" heatid="19436" lane="6" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="176" reactiontime="+95" swimtime="00:00:45.04" resultid="18524" heatid="19550" lane="8" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-07-18" firstname="Ihor" gender="M" lastname="Shchotkin" nation="UKR" athleteid="17613">
              <RESULTS>
                <RESULT eventid="1079" points="520" reactiontime="+73" swimtime="00:00:25.19" resultid="17614" heatid="19303" lane="8" entrytime="00:00:25.00" />
                <RESULT eventid="1273" points="539" reactiontime="+73" swimtime="00:00:55.21" resultid="17615" heatid="19387" lane="7" entrytime="00:00:56.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="490" reactiontime="+83" swimtime="00:00:27.64" resultid="17616" heatid="19462" lane="1" entrytime="00:00:27.50" />
                <RESULT eventid="1681" points="546" reactiontime="+69" swimtime="00:00:30.88" resultid="17617" heatid="19559" lane="5" entrytime="00:00:31.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-06-28" firstname="Valentyna" gender="F" lastname="Kvita" nation="UKR" athleteid="17590">
              <RESULTS>
                <RESULT eventid="1096" points="527" reactiontime="+92" swimtime="00:02:30.80" resultid="17591" heatid="19309" lane="3" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                    <SPLIT distance="100" swimtime="00:01:10.41" />
                    <SPLIT distance="150" swimtime="00:01:54.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="604" reactiontime="+89" swimtime="00:01:00.21" resultid="17592" heatid="19372" lane="5" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="580" reactiontime="+93" swimtime="00:02:12.78" resultid="17593" heatid="19484" lane="3" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.39" />
                    <SPLIT distance="100" swimtime="00:01:03.50" />
                    <SPLIT distance="150" swimtime="00:01:37.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="545" reactiontime="+100" swimtime="00:04:47.01" resultid="17594" heatid="19694" lane="2" entrytime="00:04:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                    <SPLIT distance="100" swimtime="00:01:06.69" />
                    <SPLIT distance="150" swimtime="00:01:42.41" />
                    <SPLIT distance="200" swimtime="00:02:18.82" />
                    <SPLIT distance="250" swimtime="00:02:55.80" />
                    <SPLIT distance="300" swimtime="00:03:33.02" />
                    <SPLIT distance="350" swimtime="00:04:10.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-04-22" firstname="Volodymyr" gender="M" lastname="Rybko" nation="UKR" athleteid="17576">
              <RESULTS>
                <RESULT eventid="1113" points="311" reactiontime="+79" swimtime="00:02:41.70" resultid="17577" heatid="19315" lane="2" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                    <SPLIT distance="100" swimtime="00:01:15.28" />
                    <SPLIT distance="150" swimtime="00:02:05.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14207" points="344" reactiontime="+93" swimtime="00:20:09.46" resultid="17578" heatid="19623" lane="2" entrytime="00:19:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.03" />
                    <SPLIT distance="100" swimtime="00:01:11.91" />
                    <SPLIT distance="150" swimtime="00:01:51.24" />
                    <SPLIT distance="200" swimtime="00:02:31.50" />
                    <SPLIT distance="250" swimtime="00:03:11.29" />
                    <SPLIT distance="350" swimtime="00:04:32.02" />
                    <SPLIT distance="400" swimtime="00:05:12.33" />
                    <SPLIT distance="600" swimtime="00:07:52.97" />
                    <SPLIT distance="700" swimtime="00:09:13.32" />
                    <SPLIT distance="750" swimtime="00:09:52.78" />
                    <SPLIT distance="900" swimtime="00:11:58.42" />
                    <SPLIT distance="950" swimtime="00:12:41.94" />
                    <SPLIT distance="1050" swimtime="00:14:04.77" />
                    <SPLIT distance="1150" swimtime="00:15:28.56" />
                    <SPLIT distance="1200" swimtime="00:16:10.04" />
                    <SPLIT distance="1400" swimtime="00:18:54.00" />
                    <SPLIT distance="1450" swimtime="00:19:33.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="419" reactiontime="+81" swimtime="00:01:00.05" resultid="17579" heatid="19385" lane="6" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="362" reactiontime="+80" swimtime="00:01:10.55" resultid="17580" heatid="19406" lane="6" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="360" reactiontime="+75" swimtime="00:00:30.64" resultid="17581" heatid="19461" lane="0" entrytime="00:00:29.00" />
                <RESULT eventid="1578" points="319" reactiontime="+87" swimtime="00:05:44.38" resultid="17582" heatid="19511" lane="8" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                    <SPLIT distance="100" swimtime="00:01:23.34" />
                    <SPLIT distance="150" swimtime="00:02:52.10" />
                    <SPLIT distance="200" swimtime="00:03:43.75" />
                    <SPLIT distance="250" swimtime="00:04:34.03" />
                    <SPLIT distance="300" swimtime="00:05:10.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="17583" heatid="19523" lane="9" entrytime="00:01:09.00" />
                <RESULT eventid="1744" points="372" reactiontime="+80" swimtime="00:04:54.91" resultid="17584" heatid="19707" lane="8" entrytime="00:04:49.00">
                  <SPLITS>
                    <SPLIT distance="250" swimtime="00:03:03.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Euro-Lviv MSC - kat.C" number="2">
              <RESULTS>
                <RESULT eventid="1381" points="473" reactiontime="+64" swimtime="00:01:56.09" resultid="17654" heatid="19424" lane="8" entrytime="00:02:00.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.49" />
                    <SPLIT distance="100" swimtime="00:01:03.38" />
                    <SPLIT distance="150" swimtime="00:01:30.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17576" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="17613" number="2" reactiontime="+21" />
                    <RELAYPOSITION athleteid="17607" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="17585" number="4" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Euro-Lviv MSC - kat.C" number="3">
              <RESULTS>
                <RESULT eventid="1548" points="517" reactiontime="+77" swimtime="00:01:42.86" resultid="17655" heatid="19502" lane="3" entrytime="00:01:44.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.71" />
                    <SPLIT distance="100" swimtime="00:00:50.24" />
                    <SPLIT distance="150" swimtime="00:01:17.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17613" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="17585" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="17576" number="3" reactiontime="+26" />
                    <RELAYPOSITION athleteid="17607" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" name="Euro-Lviv MSC - kat.C" number="4">
              <RESULTS>
                <RESULT eventid="1525" points="395" reactiontime="+84" swimtime="00:02:08.37" resultid="17656" heatid="19498" lane="3" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                    <SPLIT distance="100" swimtime="00:01:08.52" />
                    <SPLIT distance="150" swimtime="00:01:40.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17643" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="17627" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="17595" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="17590" number="4" reactiontime="+52" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Euro-Lviv MSC - kat.C" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="530" reactiontime="+80" swimtime="00:01:49.38" resultid="17653" heatid="19322" lane="5" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.99" />
                    <SPLIT distance="100" swimtime="00:00:50.20" />
                    <SPLIT distance="150" swimtime="00:01:21.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17613" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="17585" number="2" reactiontime="+38" />
                    <RELAYPOSITION athleteid="17595" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="17590" number="4" reactiontime="+52" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Euro-Lviv MSC - kat.D" number="5">
              <RESULTS>
                <RESULT eventid="1698" points="429" reactiontime="+78" swimtime="00:02:08.78" resultid="17657" heatid="19564" lane="1" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.94" />
                    <SPLIT distance="100" swimtime="00:01:10.98" />
                    <SPLIT distance="150" swimtime="00:01:37.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17627" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="17613" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="17607" number="3" reactiontime="+29" />
                    <RELAYPOSITION athleteid="17595" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="DOL" clubid="18479" name="Fitness Academy Wrocław">
          <CONTACT name="Wolny Dariusz" phone="603630870" />
          <ATHLETES>
            <ATHLETE birthdate="1986-08-04" firstname="Joanna" gender="F" lastname="Chojcan" nation="POL" athleteid="18480">
              <RESULTS>
                <RESULT eventid="1096" status="DNS" swimtime="00:00:00.00" resultid="18481" heatid="19307" lane="1" entrytime="00:03:07.00" />
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="18482" heatid="19340" lane="9" entrytime="00:00:37.50" />
                <RESULT eventid="1324" status="DNS" swimtime="00:00:00.00" resultid="18483" heatid="19412" lane="6" entrytime="00:03:15.00" />
                <RESULT eventid="1457" status="DNS" swimtime="00:00:00.00" resultid="18484" heatid="19468" lane="8" entrytime="00:01:23.00" />
                <RESULT eventid="1555" status="DNS" swimtime="00:00:00.00" resultid="18485" heatid="19504" lane="3" entrytime="00:06:35.00" />
                <RESULT eventid="1595" status="DNS" swimtime="00:00:00.00" resultid="18486" heatid="19514" lane="9" entrytime="00:01:30.00" />
                <RESULT eventid="1630" status="DNS" swimtime="00:00:00.00" resultid="18487" heatid="19528" lane="8" entrytime="00:03:05.00" />
                <RESULT eventid="1062" status="DNS" swimtime="00:00:00.00" resultid="18953" heatid="19280" lane="6" entrytime="00:00:33.33" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="15682" name="Gdynia Masters">
          <CONTACT email="k.mysiak@wpit.am.gdynia.pl" name="Mysiak" />
          <ATHLETES>
            <ATHLETE birthdate="1950-01-01" firstname="Czesław" gender="M" lastname="Mikołajczyk" nation="POL" athleteid="15824">
              <RESULTS>
                <RESULT eventid="14189" points="103" reactiontime="+100" swimtime="00:15:45.60" resultid="15825" heatid="19615" lane="0" entrytime="00:16:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.65" />
                    <SPLIT distance="100" swimtime="00:01:46.31" />
                    <SPLIT distance="150" swimtime="00:03:47.18" />
                    <SPLIT distance="200" swimtime="00:05:48.73" />
                    <SPLIT distance="250" swimtime="00:06:50.57" />
                    <SPLIT distance="600" swimtime="00:12:52.66" />
                    <SPLIT distance="650" swimtime="00:13:52.17" />
                    <SPLIT distance="750" swimtime="00:14:49.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="56" reactiontime="+106" swimtime="00:04:42.89" resultid="15826" heatid="19414" lane="5" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.00" />
                    <SPLIT distance="100" swimtime="00:02:16.48" />
                    <SPLIT distance="150" swimtime="00:03:29.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="90" reactiontime="+105" swimtime="00:08:45.23" resultid="15827" heatid="19507" lane="6" entrytime="00:08:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.01" />
                    <SPLIT distance="100" swimtime="00:03:33.15" />
                    <SPLIT distance="150" swimtime="00:04:43.45" />
                    <SPLIT distance="200" swimtime="00:05:51.41" />
                    <SPLIT distance="250" swimtime="00:06:55.37" />
                    <SPLIT distance="350" swimtime="00:07:53.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="15828" heatid="19517" lane="2" entrytime="00:02:05.00" />
                <RESULT eventid="1681" points="138" reactiontime="+99" swimtime="00:00:48.86" resultid="15829" heatid="19549" lane="8" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Andrzej" gender="M" lastname="Jacaszek" nation="POL" athleteid="15820">
              <RESULTS>
                <RESULT eventid="1239" points="209" reactiontime="+106" swimtime="00:03:22.84" resultid="15821" heatid="19361" lane="7" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.81" />
                    <SPLIT distance="150" swimtime="00:02:31.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="233" reactiontime="+89" swimtime="00:01:30.33" resultid="15822" heatid="19437" lane="0" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="223" reactiontime="+109" swimtime="00:00:41.63" resultid="15823" heatid="19551" lane="1" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="Jan Maciej" gender="M" lastname="Boboli" nation="POL" athleteid="15800">
              <RESULTS>
                <RESULT eventid="1079" points="152" reactiontime="+83" swimtime="00:00:37.96" resultid="15801" heatid="19287" lane="7" entrytime="00:00:37.00" />
                <RESULT eventid="1205" points="54" reactiontime="+78" swimtime="00:00:58.50" resultid="15802" heatid="19343" lane="3" entrytime="00:00:57.00" />
                <RESULT eventid="1273" points="96" reactiontime="+90" swimtime="00:01:37.94" resultid="15803" heatid="19375" lane="5" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="139" reactiontime="+88" swimtime="00:00:42.02" resultid="15804" heatid="19452" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1681" points="58" reactiontime="+92" swimtime="00:01:05.19" resultid="15805" heatid="19547" lane="4" entrytime="00:00:58.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-01-01" firstname="Andrzej" gender="M" lastname="Skwarło" nation="POL" athleteid="15806">
              <RESULTS>
                <RESULT eventid="1079" points="120" swimtime="00:00:41.01" resultid="15807" heatid="19287" lane="9" entrytime="00:00:38.00" />
                <RESULT eventid="1113" points="86" reactiontime="+114" swimtime="00:04:08.10" resultid="15808" heatid="19310" lane="3" entrytime="00:04:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.13" />
                    <SPLIT distance="100" swimtime="00:02:08.05" />
                    <SPLIT distance="150" swimtime="00:03:14.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="86" reactiontime="+100" swimtime="00:00:50.26" resultid="15809" heatid="19344" lane="4" entrytime="00:00:49.00" />
                <RESULT eventid="14243" points="89" reactiontime="+106" swimtime="00:01:52.28" resultid="15810" heatid="19399" lane="0" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="107" reactiontime="+114" swimtime="00:01:57.00" resultid="15811" heatid="19435" lane="6" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="62" swimtime="00:00:54.90" resultid="15812" heatid="19452" lane="0" entrytime="00:00:45.00" />
                <RESULT eventid="1613" points="51" reactiontime="+109" swimtime="00:02:09.56" resultid="15813" heatid="19518" lane="8" entrytime="00:01:52.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="148" reactiontime="+116" swimtime="00:00:47.71" resultid="15814" heatid="19549" lane="6" entrytime="00:00:46.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1934-01-01" firstname="Bogdan" gender="M" lastname="Ciundziewicki" nation="POL" athleteid="15815">
              <RESULTS>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="15816" heatid="19343" lane="6" entrytime="00:00:58.50" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="15817" heatid="19435" lane="9" entrytime="00:01:59.00" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="15818" heatid="19471" lane="5" entrytime="00:02:02.00" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="15819" heatid="19548" lane="8" entrytime="00:00:57.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="132" reactiontime="+102" swimtime="00:02:57.46" resultid="15830" heatid="19421" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.06" />
                    <SPLIT distance="100" swimtime="00:01:33.49" />
                    <SPLIT distance="150" swimtime="00:02:15.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15815" number="1" reactiontime="+102" />
                    <RELAYPOSITION athleteid="15820" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="15800" number="3" reactiontime="+29" />
                    <RELAYPOSITION athleteid="15806" number="4" reactiontime="+75" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="S4 - Przedwczesna zmiana sztafetowa (stopy pływaka utraciły kontakt z platformą startową słupka zanim poprzedzający go pływak dotkną ściany) (Time: 19:39), Na trzeciej zmianie" eventid="1548" reactiontime="+99" status="DSQ" swimtime="00:02:35.73" resultid="15831" heatid="19499" lane="6" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.89" />
                    <SPLIT distance="100" swimtime="00:01:19.00" />
                    <SPLIT distance="150" swimtime="00:01:59.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15806" number="1" reactiontime="+99" />
                    <RELAYPOSITION athleteid="15815" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="15800" number="3" reactiontime="+64" />
                    <RELAYPOSITION athleteid="15820" number="4" reactiontime="-29" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="NZWAW" nation="POL" region="WA" clubid="14975" name="K.S.niezrzeszeni.pl">
          <CONTACT name="K.S.niezrzeszeni.pl" />
          <ATHLETES>
            <ATHLETE birthdate="1959-12-27" firstname="Wojciech" gender="M" lastname="Korpetta" nation="POL" athleteid="14976">
              <RESULTS>
                <RESULT eventid="14207" points="193" reactiontime="+120" swimtime="00:24:27.23" resultid="14977" heatid="19621" lane="8" entrytime="00:24:36.59">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.96" />
                    <SPLIT distance="150" swimtime="00:02:17.69" />
                    <SPLIT distance="200" swimtime="00:03:06.85" />
                    <SPLIT distance="250" swimtime="00:03:55.94" />
                    <SPLIT distance="300" swimtime="00:04:45.89" />
                    <SPLIT distance="350" swimtime="00:05:35.21" />
                    <SPLIT distance="400" swimtime="00:06:26.06" />
                    <SPLIT distance="450" swimtime="00:07:15.29" />
                    <SPLIT distance="500" swimtime="00:08:55.26" />
                    <SPLIT distance="550" swimtime="00:10:35.23" />
                    <SPLIT distance="600" swimtime="00:11:25.31" />
                    <SPLIT distance="650" swimtime="00:13:04.79" />
                    <SPLIT distance="700" swimtime="00:15:33.61" />
                    <SPLIT distance="750" swimtime="00:16:24.22" />
                    <SPLIT distance="800" swimtime="00:17:14.17" />
                    <SPLIT distance="850" swimtime="00:18:04.02" />
                    <SPLIT distance="900" swimtime="00:18:54.82" />
                    <SPLIT distance="950" swimtime="00:19:44.65" />
                    <SPLIT distance="1000" swimtime="00:20:34.04" />
                    <SPLIT distance="1050" swimtime="00:21:22.01" />
                    <SPLIT distance="1100" swimtime="00:22:58.19" />
                    <SPLIT distance="1450" swimtime="00:23:44.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" status="DNS" swimtime="00:00:00.00" resultid="14978" heatid="19413" lane="3" />
                <RESULT eventid="1440" points="139" reactiontime="+123" swimtime="00:00:42.00" resultid="14979" heatid="19450" lane="1" />
                <RESULT eventid="1474" points="172" reactiontime="+73" swimtime="00:01:27.88" resultid="14980" heatid="19473" lane="3" entrytime="00:01:27.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="175" reactiontime="+69" swimtime="00:03:08.83" resultid="14981" heatid="19534" lane="6" entrytime="00:03:06.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.17" />
                    <SPLIT distance="100" swimtime="00:01:30.83" />
                    <SPLIT distance="150" swimtime="00:02:19.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="PDK" clubid="15647" name="Klub Plywacki Masters Krosno">
          <CONTACT city="Krosno" email="konrad_szydlo@yahoo.co.uk" internet="masters.krosoft.pl" name="Konrad Szydlo" phone="531304943" state="PDK" street="Sportowa 8" street2="(Zespol Krytych Plywalni w Krosnie)" zip="38-400" />
          <ATHLETES>
            <ATHLETE birthdate="1986-03-13" firstname="Konrad" gender="M" lastname="Szydlo" nation="POL" athleteid="15677">
              <RESULTS>
                <RESULT eventid="1079" points="299" reactiontime="+86" swimtime="00:00:30.28" resultid="15678" heatid="19293" lane="4" entrytime="00:00:29.52" />
                <RESULT eventid="14207" points="318" reactiontime="+93" swimtime="00:20:41.50" resultid="15679" heatid="19622" lane="6" entrytime="00:21:30.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                    <SPLIT distance="100" swimtime="00:01:17.50" />
                    <SPLIT distance="150" swimtime="00:01:58.75" />
                    <SPLIT distance="200" swimtime="00:02:40.85" />
                    <SPLIT distance="250" swimtime="00:03:23.26" />
                    <SPLIT distance="300" swimtime="00:04:06.01" />
                    <SPLIT distance="350" swimtime="00:04:49.02" />
                    <SPLIT distance="400" swimtime="00:05:31.32" />
                    <SPLIT distance="450" swimtime="00:06:14.57" />
                    <SPLIT distance="500" swimtime="00:06:56.93" />
                    <SPLIT distance="550" swimtime="00:07:39.81" />
                    <SPLIT distance="600" swimtime="00:08:20.98" />
                    <SPLIT distance="650" swimtime="00:09:03.27" />
                    <SPLIT distance="700" swimtime="00:09:45.81" />
                    <SPLIT distance="750" swimtime="00:10:28.35" />
                    <SPLIT distance="800" swimtime="00:11:12.04" />
                    <SPLIT distance="850" swimtime="00:11:55.18" />
                    <SPLIT distance="900" swimtime="00:12:38.60" />
                    <SPLIT distance="950" swimtime="00:13:22.17" />
                    <SPLIT distance="1000" swimtime="00:14:05.31" />
                    <SPLIT distance="1050" swimtime="00:14:49.40" />
                    <SPLIT distance="1100" swimtime="00:15:32.16" />
                    <SPLIT distance="1150" swimtime="00:16:15.46" />
                    <SPLIT distance="1200" swimtime="00:16:59.58" />
                    <SPLIT distance="1250" swimtime="00:17:43.54" />
                    <SPLIT distance="1300" swimtime="00:18:28.69" />
                    <SPLIT distance="1350" swimtime="00:19:13.97" />
                    <SPLIT distance="1400" swimtime="00:19:58.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="259" reactiontime="+75" swimtime="00:02:45.69" resultid="15680" heatid="19534" lane="4" entrytime="00:02:56.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.83" />
                    <SPLIT distance="100" swimtime="00:01:21.70" />
                    <SPLIT distance="150" swimtime="00:02:04.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="303" reactiontime="+92" swimtime="00:05:15.83" resultid="15681" heatid="19704" lane="5" entrytime="00:05:20.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.15" />
                    <SPLIT distance="100" swimtime="00:01:12.02" />
                    <SPLIT distance="150" swimtime="00:01:51.54" />
                    <SPLIT distance="200" swimtime="00:02:31.83" />
                    <SPLIT distance="250" swimtime="00:03:12.72" />
                    <SPLIT distance="300" swimtime="00:03:53.84" />
                    <SPLIT distance="350" swimtime="00:04:35.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="100504" nation="POL" region="ZG" clubid="15410" name="Klub Pływacki &quot;Totis Viribus&quot; Świebodzin" shortname="Klub Pływacki &quot;Totis Viribus&quot; ">
          <CONTACT city="Świebodzin" email="totisviribus@totisviribus.pl" internet="www.totisviribus.pl" name="Jaworski Sławomir" phone="531942331" state="LUBUS" street="Okrężna 3" zip="66-200" />
          <ATHLETES>
            <ATHLETE birthdate="1980-10-12" firstname="Ewelina" gender="F" lastname="Solak" nation="POL" athleteid="15411">
              <RESULTS>
                <RESULT eventid="1062" points="154" reactiontime="+155" swimtime="00:00:43.33" resultid="15412" heatid="19275" lane="2" />
                <RESULT eventid="1256" points="138" reactiontime="+131" swimtime="00:01:38.45" resultid="15413" heatid="19366" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="184" reactiontime="+123" swimtime="00:01:49.53" resultid="15414" heatid="19427" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="195" reactiontime="+107" swimtime="00:00:49.36" resultid="15415" heatid="19538" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-03-10" firstname="Anna" gender="F" lastname="Dunaj" nation="POL" athleteid="15421">
              <RESULTS>
                <RESULT eventid="1062" status="DNS" swimtime="00:00:00.00" resultid="15422" heatid="19275" lane="7" />
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="15423" heatid="19367" lane="1" />
                <RESULT eventid="1388" status="DNS" swimtime="00:00:00.00" resultid="15424" heatid="19426" lane="4" />
                <RESULT eventid="1664" status="DNS" swimtime="00:00:00.00" resultid="15425" heatid="19538" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-10-17" firstname="Małgorzata" gender="F" lastname="Maciecka" nation="POL" athleteid="15416">
              <RESULTS>
                <RESULT eventid="1062" status="DNS" swimtime="00:00:00.00" resultid="15417" heatid="19275" lane="6" />
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="15418" heatid="19367" lane="0" />
                <RESULT eventid="1388" status="DNS" swimtime="00:00:00.00" resultid="15419" heatid="19426" lane="6" />
                <RESULT eventid="1664" status="DNS" swimtime="00:00:00.00" resultid="15420" heatid="19538" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-07-24" firstname="Katarzyna" gender="F" lastname="Bubienko" nation="POL" athleteid="15426">
              <RESULTS>
                <RESULT eventid="1062" points="359" reactiontime="+79" swimtime="00:00:32.68" resultid="15427" heatid="19275" lane="5" />
                <RESULT eventid="1324" status="DNS" swimtime="00:00:00.00" resultid="15428" heatid="19411" lane="1" />
                <RESULT eventid="1388" points="263" reactiontime="+85" swimtime="00:01:37.33" resultid="15429" heatid="19426" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="213" reactiontime="+85" swimtime="00:00:40.80" resultid="15430" heatid="19444" lane="3" />
                <RESULT eventid="1664" points="302" reactiontime="+83" swimtime="00:00:42.65" resultid="15431" heatid="19538" lane="4" />
                <RESULT eventid="1222" points="234" reactiontime="+84" swimtime="00:03:38.28" resultid="15433" heatid="19354" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.89" />
                    <SPLIT distance="100" swimtime="00:01:41.02" />
                    <SPLIT distance="150" swimtime="00:02:38.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="15432" heatid="19497" lane="6">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15426" number="1" />
                    <RELAYPOSITION athleteid="15411" number="2" />
                    <RELAYPOSITION athleteid="15421" number="3" />
                    <RELAYPOSITION athleteid="15416" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MAKO" nation="POL" region="WAR" clubid="16894" name="Klub Sportowy MAKO">
          <CONTACT email="ania.plywanie@gmail.com" name="Dąbrowska Anna" phone="601480280" />
          <ATHLETES>
            <ATHLETE birthdate="1980-06-07" firstname="Piotr" gender="M" lastname="Kieżun" nation="POL" athleteid="16938">
              <RESULTS>
                <RESULT eventid="1079" points="266" reactiontime="+100" swimtime="00:00:31.47" resultid="16939" heatid="19290" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1273" points="214" reactiontime="+85" swimtime="00:01:15.07" resultid="16940" heatid="19379" lane="7" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="197" reactiontime="+87" swimtime="00:02:50.57" resultid="16941" heatid="19488" lane="2" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.73" />
                    <SPLIT distance="100" swimtime="00:01:21.74" />
                    <SPLIT distance="150" swimtime="00:02:07.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="227" reactiontime="+96" swimtime="00:00:41.38" resultid="16942" heatid="19551" lane="0" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-30" firstname="Piotr" gender="M" lastname="Safrończyk" nation="POL" athleteid="16922">
              <RESULTS>
                <RESULT eventid="1079" points="605" reactiontime="+71" swimtime="00:00:23.95" resultid="16923" heatid="19304" lane="5" entrytime="00:00:23.20" />
                <RESULT eventid="1205" points="478" reactiontime="+68" swimtime="00:00:28.40" resultid="16924" heatid="19353" lane="3" entrytime="00:00:26.80" />
                <RESULT eventid="14243" status="DNS" swimtime="00:00:00.00" resultid="16925" heatid="19410" lane="3" entrytime="00:00:58.20" />
                <RESULT eventid="1440" points="592" reactiontime="+71" swimtime="00:00:25.96" resultid="16926" heatid="19464" lane="4" entrytime="00:00:24.90" />
                <RESULT eventid="1681" points="671" reactiontime="+67" swimtime="00:00:28.83" resultid="16927" heatid="19560" lane="5" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-04-29" firstname="Artur" gender="M" lastname="Pietrzak" nation="POL" athleteid="16950">
              <RESULTS>
                <RESULT eventid="1440" points="521" reactiontime="+73" swimtime="00:00:27.09" resultid="16951" heatid="19463" lane="7" entrytime="00:00:27.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-05-20" firstname="Anna" gender="F" lastname="Dąbrowska" nation="POL" athleteid="16916">
              <RESULTS>
                <RESULT eventid="1062" points="266" reactiontime="+97" swimtime="00:00:36.11" resultid="16917" heatid="19279" lane="5" entrytime="00:00:34.58" />
                <RESULT eventid="1256" points="254" reactiontime="+106" swimtime="00:01:20.30" resultid="16918" heatid="19370" lane="8" entrytime="00:01:18.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="207" reactiontime="+99" swimtime="00:00:41.18" resultid="16919" heatid="19446" lane="3" entrytime="00:00:39.20" />
                <RESULT eventid="1491" points="225" reactiontime="+89" swimtime="00:03:02.04" resultid="16920" heatid="19482" lane="0" entrytime="00:03:01.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.41" />
                    <SPLIT distance="100" swimtime="00:01:27.24" />
                    <SPLIT distance="150" swimtime="00:02:15.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="176" reactiontime="+126" swimtime="00:01:37.34" resultid="16921" heatid="19513" lane="4" entrytime="00:01:32.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-05-14" firstname="Dominik" gender="M" lastname="Markowski" nation="POL" athleteid="16932">
              <RESULTS>
                <RESULT eventid="1079" points="186" reactiontime="+87" swimtime="00:00:35.47" resultid="16933" heatid="19287" lane="2" entrytime="00:00:37.00" />
                <RESULT eventid="1205" points="159" reactiontime="+80" swimtime="00:00:41.00" resultid="16934" heatid="19342" lane="1" />
                <RESULT eventid="1273" points="170" reactiontime="+81" swimtime="00:01:21.09" resultid="16935" heatid="19376" lane="7" entrytime="00:01:27.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="141" reactiontime="+78" swimtime="00:01:33.78" resultid="16936" heatid="19472" lane="2" entrytime="00:01:41.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="16937" heatid="19701" lane="8" entrytime="00:06:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-09" firstname="Paweł" gender="M" lastname="Rurak" nation="POL" athleteid="16928">
              <RESULTS>
                <RESULT eventid="1079" points="624" reactiontime="+73" swimtime="00:00:23.70" resultid="16929" heatid="19304" lane="4" entrytime="00:00:23.20" />
                <RESULT eventid="1205" points="586" reactiontime="+70" swimtime="00:00:26.54" resultid="16930" heatid="19353" lane="4" entrytime="00:00:25.90" />
                <RESULT eventid="14243" status="DNS" swimtime="00:00:00.00" resultid="16931" heatid="19410" lane="5" entrytime="00:00:57.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-07-11" firstname="Paweł" gender="M" lastname="Adamowicz" nation="POL" athleteid="16943">
              <RESULTS>
                <RESULT eventid="1079" points="128" reactiontime="+78" swimtime="00:00:40.12" resultid="16944" heatid="19286" lane="7" entrytime="00:00:39.39" />
                <RESULT eventid="14243" points="95" reactiontime="+85" swimtime="00:01:50.10" resultid="16945" heatid="19397" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="149" reactiontime="+87" swimtime="00:01:44.86" resultid="16946" heatid="19436" lane="1" entrytime="00:01:41.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="178" reactiontime="+82" swimtime="00:00:44.84" resultid="16947" heatid="19550" lane="1" entrytime="00:00:44.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-06-01" firstname="Robert" gender="M" lastname="Wilk" nation="POL" athleteid="16948" />
            <ATHLETE birthdate="1989-06-25" firstname="Krzysztof" gender="M" lastname="Wilk" nation="POL" athleteid="16949" />
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="626" reactiontime="+66" swimtime="00:01:45.78" resultid="16952" heatid="19424" lane="4" entrytime="00:01:42.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.66" />
                    <SPLIT distance="100" swimtime="00:00:55.53" />
                    <SPLIT distance="150" swimtime="00:01:22.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16928" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="16922" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="16950" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="16948" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="16953" points="671" reactiontime="+70" status="EXH" swimtime="00:03:29.36" resultid="16962" heatid="19425" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.84" />
                    <SPLIT distance="100" swimtime="00:00:51.94" />
                    <SPLIT distance="150" swimtime="00:01:15.89" />
                    <SPLIT distance="200" swimtime="00:01:43.51" />
                    <SPLIT distance="250" swimtime="00:02:08.85" />
                    <SPLIT distance="300" swimtime="00:02:37.53" />
                    <SPLIT distance="350" swimtime="00:03:01.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16928" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="16948" number="2" reactiontime="+28" />
                    <RELAYPOSITION athleteid="16949" number="3" reactiontime="+28" />
                    <RELAYPOSITION athleteid="16922" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="KS WAR" nation="POL" region="WIE" clubid="17144" name="Klub Sportowy Warta Poznań">
          <CONTACT city="Poznań" email="jacek.thiem@gmail.com" name="Thiem Jacek" phone="502499565" state="WIE" street="Osiedle Dębina 19 m 34" zip="61-450" />
          <ATHLETES>
            <ATHLETE birthdate="1957-10-01" firstname="Grażyna" gender="F" lastname="Drela" nation="POL" license="100115700493" athleteid="17152">
              <RESULTS>
                <RESULT eventid="1062" points="277" reactiontime="+93" swimtime="00:00:35.61" resultid="17153" heatid="19279" lane="1" entrytime="00:00:36.00" />
                <RESULT eventid="1222" points="290" reactiontime="+94" swimtime="00:03:23.09" resultid="17154" heatid="19356" lane="5" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.34" />
                    <SPLIT distance="100" swimtime="00:01:37.84" />
                    <SPLIT distance="150" swimtime="00:02:31.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="278" reactiontime="+96" swimtime="00:01:26.77" resultid="17155" heatid="19392" lane="1" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="301" reactiontime="+86" swimtime="00:01:32.99" resultid="17156" heatid="19430" lane="8" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="233" reactiontime="+99" swimtime="00:02:59.95" resultid="17157" heatid="19482" lane="1" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.88" />
                    <SPLIT distance="100" swimtime="00:01:26.30" />
                    <SPLIT distance="150" swimtime="00:02:13.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="294" reactiontime="+87" swimtime="00:00:43.04" resultid="17158" heatid="19542" lane="9" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-19" firstname="Przemysław" gender="M" lastname="Waraczewski" nation="POL" license="100115700344" athleteid="17177">
              <RESULTS>
                <RESULT eventid="1113" points="235" reactiontime="+91" swimtime="00:02:57.62" resultid="17178" heatid="19312" lane="4" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.62" />
                    <SPLIT distance="100" swimtime="00:01:27.24" />
                    <SPLIT distance="150" swimtime="00:02:15.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="267" reactiontime="+89" swimtime="00:03:06.81" resultid="17179" heatid="19363" lane="8" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.80" />
                    <SPLIT distance="100" swimtime="00:01:26.66" />
                    <SPLIT distance="150" swimtime="00:02:15.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="290" reactiontime="+83" swimtime="00:01:23.97" resultid="17180" heatid="19439" lane="9" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="308" reactiontime="+95" swimtime="00:00:37.35" resultid="17181" heatid="19553" lane="0" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-27" firstname="Dariusz" gender="M" lastname="Janyga" nation="POL" license="100115700346" athleteid="17219">
              <RESULTS>
                <RESULT comment="O4 - Start wykonany przed sygnłem (przedwczesny start) (Time: 15:34)" eventid="1079" reactiontime="+72" status="DSQ" swimtime="00:00:28.21" resultid="17220" heatid="19294" lane="9" entrytime="00:00:29.50" />
                <RESULT eventid="14189" points="323" reactiontime="+103" swimtime="00:10:45.66" resultid="17221" heatid="19616" lane="5" entrytime="00:10:45.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                    <SPLIT distance="100" swimtime="00:01:15.32" />
                    <SPLIT distance="150" swimtime="00:01:54.94" />
                    <SPLIT distance="200" swimtime="00:02:35.47" />
                    <SPLIT distance="250" swimtime="00:03:15.76" />
                    <SPLIT distance="300" swimtime="00:03:56.60" />
                    <SPLIT distance="350" swimtime="00:04:37.58" />
                    <SPLIT distance="400" swimtime="00:05:18.23" />
                    <SPLIT distance="450" swimtime="00:05:59.04" />
                    <SPLIT distance="500" swimtime="00:06:40.13" />
                    <SPLIT distance="550" swimtime="00:07:21.42" />
                    <SPLIT distance="600" swimtime="00:08:03.03" />
                    <SPLIT distance="650" swimtime="00:08:44.08" />
                    <SPLIT distance="700" swimtime="00:09:25.50" />
                    <SPLIT distance="750" swimtime="00:10:06.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="308" swimtime="00:00:32.89" resultid="17222" heatid="19349" lane="7" entrytime="00:00:33.50" />
                <RESULT eventid="1474" points="333" reactiontime="+80" swimtime="00:01:10.56" resultid="17223" heatid="19476" lane="1" entrytime="00:01:12.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="340" reactiontime="+93" swimtime="00:02:22.31" resultid="17224" heatid="19492" lane="4" entrytime="00:02:22.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                    <SPLIT distance="100" swimtime="00:01:09.02" />
                    <SPLIT distance="150" swimtime="00:01:45.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="295" swimtime="00:02:38.62" resultid="17225" heatid="19536" lane="7" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.32" />
                    <SPLIT distance="150" swimtime="00:01:58.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="335" reactiontime="+97" swimtime="00:05:05.45" resultid="17226" heatid="19704" lane="3" entrytime="00:05:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.17" />
                    <SPLIT distance="100" swimtime="00:01:12.86" />
                    <SPLIT distance="150" swimtime="00:01:51.33" />
                    <SPLIT distance="200" swimtime="00:02:30.45" />
                    <SPLIT distance="250" swimtime="00:03:09.66" />
                    <SPLIT distance="300" swimtime="00:03:48.38" />
                    <SPLIT distance="350" swimtime="00:04:27.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-05-08" firstname="Anna" gender="F" lastname="Kotecka" nation="POL" license="100115600357" athleteid="17202">
              <RESULTS>
                <RESULT eventid="1165" points="231" swimtime="00:24:58.90" resultid="17203" heatid="19624" lane="7" entrytime="00:27:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.28" />
                    <SPLIT distance="100" swimtime="00:01:30.25" />
                    <SPLIT distance="150" swimtime="00:02:18.61" />
                    <SPLIT distance="200" swimtime="00:03:07.07" />
                    <SPLIT distance="250" swimtime="00:03:55.23" />
                    <SPLIT distance="300" swimtime="00:04:44.31" />
                    <SPLIT distance="350" swimtime="00:05:34.02" />
                    <SPLIT distance="400" swimtime="00:06:23.56" />
                    <SPLIT distance="450" swimtime="00:07:13.64" />
                    <SPLIT distance="500" swimtime="00:08:04.48" />
                    <SPLIT distance="550" swimtime="00:08:54.27" />
                    <SPLIT distance="600" swimtime="00:09:44.73" />
                    <SPLIT distance="650" swimtime="00:10:35.73" />
                    <SPLIT distance="700" swimtime="00:11:26.27" />
                    <SPLIT distance="750" swimtime="00:12:17.17" />
                    <SPLIT distance="800" swimtime="00:13:07.45" />
                    <SPLIT distance="850" swimtime="00:13:57.86" />
                    <SPLIT distance="900" swimtime="00:14:47.70" />
                    <SPLIT distance="950" swimtime="00:15:38.66" />
                    <SPLIT distance="1000" swimtime="00:16:29.19" />
                    <SPLIT distance="1050" swimtime="00:17:19.97" />
                    <SPLIT distance="1100" swimtime="00:18:10.40" />
                    <SPLIT distance="1150" swimtime="00:19:01.95" />
                    <SPLIT distance="1200" swimtime="00:19:53.18" />
                    <SPLIT distance="1250" swimtime="00:20:44.63" />
                    <SPLIT distance="1300" swimtime="00:21:35.98" />
                    <SPLIT distance="1350" swimtime="00:22:26.54" />
                    <SPLIT distance="1400" swimtime="00:23:17.88" />
                    <SPLIT distance="1450" swimtime="00:24:09.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="164" reactiontime="+132" swimtime="00:00:46.83" resultid="17204" heatid="19337" lane="4" entrytime="00:00:48.00" />
                <RESULT eventid="1256" points="217" swimtime="00:01:24.65" resultid="17205" heatid="19369" lane="8" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="166" reactiontime="+85" swimtime="00:01:40.05" resultid="17206" heatid="19466" lane="2" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="219" swimtime="00:03:03.52" resultid="17207" heatid="19482" lane="8" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.99" />
                    <SPLIT distance="100" swimtime="00:01:28.51" />
                    <SPLIT distance="150" swimtime="00:02:15.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="186" reactiontime="+79" swimtime="00:03:28.82" resultid="17208" heatid="19527" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.59" />
                    <SPLIT distance="100" swimtime="00:01:42.22" />
                    <SPLIT distance="150" swimtime="00:02:36.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" reactiontime="+105" status="DNS" swimtime="00:00:00.00" resultid="17209" heatid="19696" lane="1" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.54" />
                    <SPLIT distance="100" swimtime="00:01:41.15" />
                    <SPLIT distance="150" swimtime="00:02:36.96" />
                    <SPLIT distance="200" swimtime="00:03:33.24" />
                    <SPLIT distance="250" swimtime="00:04:29.83" />
                    <SPLIT distance="300" swimtime="00:05:26.66" />
                    <SPLIT distance="350" swimtime="00:06:24.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-09-08" firstname="Szymon" gender="M" lastname="Wieja" nation="POL" athleteid="17227">
              <RESULTS>
                <RESULT eventid="1079" points="377" reactiontime="+76" swimtime="00:00:28.03" resultid="17228" heatid="19298" lane="5" entrytime="00:00:27.50" />
                <RESULT eventid="1273" points="399" reactiontime="+74" swimtime="00:01:01.01" resultid="17229" heatid="19385" lane="5" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="319" swimtime="00:01:11.56" resultid="17230" heatid="19477" lane="8" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="281" reactiontime="+76" swimtime="00:01:13.38" resultid="17231" heatid="19522" lane="7" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-07-02" firstname="Tomasz" gender="M" lastname="Tomaszewski" nation="POL" license="500115700350" athleteid="17210">
              <RESULTS>
                <RESULT eventid="1205" points="396" reactiontime="+76" swimtime="00:00:30.25" resultid="17211" heatid="19351" lane="5" entrytime="00:00:30.50" />
                <RESULT eventid="1474" points="448" reactiontime="+75" swimtime="00:01:03.92" resultid="17212" heatid="19476" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="405" reactiontime="+76" swimtime="00:02:22.76" resultid="17213" heatid="19537" lane="9" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                    <SPLIT distance="100" swimtime="00:01:08.57" />
                    <SPLIT distance="150" swimtime="00:01:46.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-12" firstname="Marcin" gender="M" lastname="Szymkowiak" nation="POL" athleteid="17195">
              <RESULTS>
                <RESULT eventid="1079" points="470" reactiontime="+78" swimtime="00:00:26.05" resultid="17196" heatid="19301" lane="8" entrytime="00:00:26.00" />
                <RESULT eventid="1273" points="440" reactiontime="+89" swimtime="00:00:59.06" resultid="17197" heatid="19386" lane="1" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="418" reactiontime="+77" swimtime="00:01:07.26" resultid="17198" heatid="19407" lane="5" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="461" reactiontime="+85" swimtime="00:01:11.96" resultid="17199" heatid="19441" lane="4" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="446" reactiontime="+82" swimtime="00:00:28.52" resultid="17200" heatid="19462" lane="6" entrytime="00:00:27.50" />
                <RESULT eventid="1681" points="521" reactiontime="+73" swimtime="00:00:31.36" resultid="17201" heatid="19560" lane="9" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-10-01" firstname="Natlia" gender="F" lastname="Wiśniewska" nation="POL" athleteid="17232">
              <RESULTS>
                <RESULT eventid="1096" points="501" reactiontime="+96" swimtime="00:02:33.35" resultid="17233" heatid="19309" lane="2" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                    <SPLIT distance="100" swimtime="00:01:11.90" />
                    <SPLIT distance="150" swimtime="00:01:55.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="516" reactiontime="+86" swimtime="00:02:47.73" resultid="17234" heatid="19358" lane="4" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.92" />
                    <SPLIT distance="100" swimtime="00:01:21.10" />
                    <SPLIT distance="150" swimtime="00:02:04.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="511" reactiontime="+84" swimtime="00:01:10.84" resultid="17235" heatid="19396" lane="5" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="527" reactiontime="+87" swimtime="00:01:17.19" resultid="17236" heatid="19432" lane="4" entrytime="00:01:16.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="489" reactiontime="+89" swimtime="00:05:29.15" resultid="17237" heatid="19505" lane="3" entrytime="00:05:32.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.14" />
                    <SPLIT distance="100" swimtime="00:01:13.82" />
                    <SPLIT distance="150" swimtime="00:01:56.53" />
                    <SPLIT distance="200" swimtime="00:02:38.77" />
                    <SPLIT distance="250" swimtime="00:03:23.19" />
                    <SPLIT distance="300" swimtime="00:04:09.12" />
                    <SPLIT distance="350" swimtime="00:04:50.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="503" reactiontime="+86" swimtime="00:00:36.00" resultid="17238" heatid="19545" lane="7" entrytime="00:00:36.83" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-26" firstname="Stanisław" gender="M" lastname="Kaczmarek" nation="POL" license="100115700354" athleteid="17168">
              <RESULTS>
                <RESULT eventid="1113" points="511" reactiontime="+72" swimtime="00:02:17.05" resultid="17169" heatid="19318" lane="7" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.50" />
                    <SPLIT distance="100" swimtime="00:01:05.90" />
                    <SPLIT distance="150" swimtime="00:01:45.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14189" points="513" reactiontime="+73" swimtime="00:09:13.63" resultid="17170" heatid="19618" lane="4" entrytime="00:08:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.15" />
                    <SPLIT distance="100" swimtime="00:01:05.43" />
                    <SPLIT distance="150" swimtime="00:01:40.25" />
                    <SPLIT distance="200" swimtime="00:02:14.98" />
                    <SPLIT distance="250" swimtime="00:02:49.58" />
                    <SPLIT distance="300" swimtime="00:03:24.23" />
                    <SPLIT distance="350" swimtime="00:03:59.05" />
                    <SPLIT distance="400" swimtime="00:04:33.99" />
                    <SPLIT distance="450" swimtime="00:05:08.76" />
                    <SPLIT distance="500" swimtime="00:05:43.29" />
                    <SPLIT distance="550" swimtime="00:06:18.29" />
                    <SPLIT distance="600" swimtime="00:06:53.53" />
                    <SPLIT distance="650" swimtime="00:07:29.02" />
                    <SPLIT distance="700" swimtime="00:08:04.16" />
                    <SPLIT distance="750" swimtime="00:08:39.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="484" reactiontime="+74" swimtime="00:02:33.39" resultid="17171" heatid="19365" lane="6" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                    <SPLIT distance="100" swimtime="00:01:14.45" />
                    <SPLIT distance="150" swimtime="00:01:54.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="498" reactiontime="+74" swimtime="00:02:16.88" resultid="17172" heatid="19418" lane="3" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.40" />
                    <SPLIT distance="100" swimtime="00:01:05.14" />
                    <SPLIT distance="150" swimtime="00:01:40.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="534" reactiontime="+71" swimtime="00:02:02.47" resultid="17173" heatid="19496" lane="6" entrytime="00:01:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.97" />
                    <SPLIT distance="100" swimtime="00:01:00.05" />
                    <SPLIT distance="150" swimtime="00:01:31.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="511" reactiontime="+74" swimtime="00:04:54.54" resultid="17174" heatid="19512" lane="6" entrytime="00:04:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.09" />
                    <SPLIT distance="100" swimtime="00:01:05.69" />
                    <SPLIT distance="150" swimtime="00:01:45.41" />
                    <SPLIT distance="200" swimtime="00:02:24.32" />
                    <SPLIT distance="250" swimtime="00:03:05.81" />
                    <SPLIT distance="300" swimtime="00:03:48.43" />
                    <SPLIT distance="350" swimtime="00:04:22.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="481" reactiontime="+85" swimtime="00:00:32.22" resultid="17175" heatid="19559" lane="1" entrytime="00:00:31.80" />
                <RESULT eventid="1744" points="536" reactiontime="+72" swimtime="00:04:21.14" resultid="17176" heatid="19708" lane="5" entrytime="00:04:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.93" />
                    <SPLIT distance="100" swimtime="00:01:02.41" />
                    <SPLIT distance="150" swimtime="00:01:35.23" />
                    <SPLIT distance="200" swimtime="00:02:08.39" />
                    <SPLIT distance="250" swimtime="00:02:41.68" />
                    <SPLIT distance="300" swimtime="00:03:15.10" />
                    <SPLIT distance="350" swimtime="00:03:48.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-02-03" firstname="Paweł" gender="M" lastname="Olszewski" nation="POL" license="100115700350" athleteid="17214">
              <RESULTS>
                <RESULT eventid="1273" points="406" reactiontime="+78" swimtime="00:01:00.66" resultid="17215" heatid="19384" lane="9" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="367" reactiontime="+75" swimtime="00:00:30.44" resultid="17216" heatid="19457" lane="6" entrytime="00:00:31.50" />
                <RESULT eventid="1508" points="398" reactiontime="+79" swimtime="00:02:15.06" resultid="17217" heatid="19493" lane="7" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                    <SPLIT distance="100" swimtime="00:01:07.29" />
                    <SPLIT distance="150" swimtime="00:01:42.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="374" reactiontime="+84" swimtime="00:04:54.56" resultid="17218" heatid="19706" lane="2" entrytime="00:04:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:09.96" />
                    <SPLIT distance="150" swimtime="00:01:47.64" />
                    <SPLIT distance="200" swimtime="00:02:26.10" />
                    <SPLIT distance="250" swimtime="00:03:04.20" />
                    <SPLIT distance="300" swimtime="00:03:42.25" />
                    <SPLIT distance="350" swimtime="00:04:19.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-02-17" firstname="Jacek" gender="M" lastname="Thiem" nation="POL" license="100115700345" athleteid="17145">
              <RESULTS>
                <RESULT eventid="14207" points="175" reactiontime="+122" swimtime="00:25:13.62" resultid="17146" heatid="19620" lane="5" entrytime="00:26:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.17" />
                    <SPLIT distance="100" swimtime="00:01:30.49" />
                    <SPLIT distance="150" swimtime="00:02:19.44" />
                    <SPLIT distance="200" swimtime="00:03:08.20" />
                    <SPLIT distance="250" swimtime="00:03:57.92" />
                    <SPLIT distance="300" swimtime="00:04:48.74" />
                    <SPLIT distance="350" swimtime="00:05:39.65" />
                    <SPLIT distance="400" swimtime="00:06:30.61" />
                    <SPLIT distance="450" swimtime="00:07:22.60" />
                    <SPLIT distance="500" swimtime="00:08:14.08" />
                    <SPLIT distance="550" swimtime="00:09:05.60" />
                    <SPLIT distance="600" swimtime="00:09:57.22" />
                    <SPLIT distance="650" swimtime="00:10:47.86" />
                    <SPLIT distance="700" swimtime="00:11:39.33" />
                    <SPLIT distance="750" swimtime="00:12:30.53" />
                    <SPLIT distance="800" swimtime="00:13:21.36" />
                    <SPLIT distance="850" swimtime="00:14:12.90" />
                    <SPLIT distance="900" swimtime="00:15:03.32" />
                    <SPLIT distance="950" swimtime="00:15:54.62" />
                    <SPLIT distance="1000" swimtime="00:16:46.76" />
                    <SPLIT distance="1050" swimtime="00:17:38.10" />
                    <SPLIT distance="1100" swimtime="00:18:29.93" />
                    <SPLIT distance="1150" swimtime="00:19:21.79" />
                    <SPLIT distance="1200" swimtime="00:20:13.79" />
                    <SPLIT distance="1250" swimtime="00:21:05.13" />
                    <SPLIT distance="1300" swimtime="00:21:56.78" />
                    <SPLIT distance="1350" swimtime="00:22:48.04" />
                    <SPLIT distance="1400" swimtime="00:23:37.44" />
                    <SPLIT distance="1450" swimtime="00:24:27.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="187" reactiontime="+113" swimtime="00:03:09.80" resultid="17147" heatid="19415" lane="4" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.95" />
                    <SPLIT distance="100" swimtime="00:01:32.29" />
                    <SPLIT distance="150" swimtime="00:02:21.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="208" reactiontime="+91" swimtime="00:00:36.78" resultid="17148" heatid="19453" lane="2" entrytime="00:00:37.00" />
                <RESULT eventid="1508" points="200" reactiontime="+105" swimtime="00:02:49.74" resultid="17149" heatid="19490" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.18" />
                    <SPLIT distance="150" swimtime="00:02:06.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="180" reactiontime="+104" swimtime="00:01:25.00" resultid="17150" heatid="19519" lane="6" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="17151" heatid="19703" lane="7" entrytime="00:05:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-10-01" firstname="Rusłana" gender="F" lastname="Dembecka" nation="POL" license="100115600353" athleteid="17188">
              <RESULTS>
                <RESULT eventid="1147" status="OTL" swimtime="00:19:06.40" resultid="17189" heatid="19594" lane="5" entrytime="00:17:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.06" />
                    <SPLIT distance="100" swimtime="00:02:10.87" />
                    <SPLIT distance="150" swimtime="00:03:23.47" />
                    <SPLIT distance="200" swimtime="00:04:35.98" />
                    <SPLIT distance="250" swimtime="00:05:50.04" />
                    <SPLIT distance="300" swimtime="00:07:03.81" />
                    <SPLIT distance="350" swimtime="00:08:17.49" />
                    <SPLIT distance="400" swimtime="00:09:31.06" />
                    <SPLIT distance="450" swimtime="00:10:44.58" />
                    <SPLIT distance="500" swimtime="00:11:57.22" />
                    <SPLIT distance="550" swimtime="00:13:09.24" />
                    <SPLIT distance="600" swimtime="00:14:21.50" />
                    <SPLIT distance="650" swimtime="00:15:33.98" />
                    <SPLIT distance="700" swimtime="00:16:46.47" />
                    <SPLIT distance="750" swimtime="00:17:58.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="93" reactiontime="+91" swimtime="00:00:56.64" resultid="17190" heatid="19336" lane="5" entrytime="00:01:00.00" />
                <RESULT eventid="1256" points="82" reactiontime="+124" swimtime="00:01:56.72" resultid="17191" heatid="19367" lane="3" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="64" reactiontime="+90" swimtime="00:02:17.30" resultid="17192" heatid="19465" lane="4" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="67" reactiontime="+105" swimtime="00:04:52.27" resultid="17193" heatid="19526" lane="2" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.12" />
                    <SPLIT distance="100" swimtime="00:02:26.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="75" reactiontime="+137" swimtime="00:09:13.96" resultid="17194" heatid="19695" lane="8" entrytime="00:09:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-08-31" firstname="Bartłomiej" gender="M" lastname="Zadorożny" nation="POL" license="500115700461" athleteid="17182">
              <RESULTS>
                <RESULT eventid="1079" points="436" reactiontime="+78" swimtime="00:00:26.70" resultid="17183" heatid="19298" lane="7" entrytime="00:00:27.53" />
                <RESULT eventid="1239" points="409" reactiontime="+84" swimtime="00:02:42.14" resultid="17184" heatid="19364" lane="1" entrytime="00:02:48.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                    <SPLIT distance="100" swimtime="00:01:16.04" />
                    <SPLIT distance="150" swimtime="00:01:58.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="407" reactiontime="+81" swimtime="00:01:00.64" resultid="17185" heatid="19384" lane="3" entrytime="00:01:00.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="474" reactiontime="+81" swimtime="00:01:11.29" resultid="17186" heatid="19440" lane="4" entrytime="00:01:15.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="462" reactiontime="+84" swimtime="00:00:32.66" resultid="17187" heatid="19556" lane="5" entrytime="00:00:34.37" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1381" points="474" reactiontime="+67" swimtime="00:01:56.01" resultid="17242" heatid="19424" lane="9" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.64" />
                    <SPLIT distance="100" swimtime="00:01:02.64" />
                    <SPLIT distance="150" swimtime="00:01:30.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17210" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="17182" number="2" reactiontime="+70" />
                    <RELAYPOSITION athleteid="17168" number="3" reactiontime="+18" />
                    <RELAYPOSITION athleteid="17195" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="1381" points="292" swimtime="00:02:16.37" resultid="17243" heatid="19422" lane="7" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                    <SPLIT distance="100" swimtime="00:01:11.90" />
                    <SPLIT distance="150" swimtime="00:01:48.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17219" number="1" />
                    <RELAYPOSITION athleteid="17177" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="17145" number="3" reactiontime="+79" />
                    <RELAYPOSITION athleteid="17214" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="7">
              <RESULTS>
                <RESULT eventid="1548" points="469" reactiontime="+86" swimtime="00:01:46.24" resultid="17245" heatid="19502" lane="0" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.64" />
                    <SPLIT distance="100" swimtime="00:00:54.27" />
                    <SPLIT distance="150" swimtime="00:01:20.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17210" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="17227" number="2" reactiontime="+24" />
                    <RELAYPOSITION athleteid="17168" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="17195" number="4" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="8">
              <RESULTS>
                <RESULT eventid="1548" points="318" reactiontime="+98" swimtime="00:02:00.95" resultid="17246" heatid="19500" lane="4" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.67" />
                    <SPLIT distance="100" swimtime="00:01:01.37" />
                    <SPLIT distance="150" swimtime="00:01:33.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17219" number="1" reactiontime="+98" />
                    <RELAYPOSITION athleteid="17177" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="17145" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="17214" number="4" reactiontime="+15" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="3">
              <RESULTS>
                <RESULT eventid="1358" status="DNS" swimtime="00:00:00.00" resultid="17241" heatid="19420" lane="9" entrytime="00:03:10.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17202" number="1" />
                    <RELAYPOSITION athleteid="17188" number="2" />
                    <RELAYPOSITION athleteid="17152" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="6">
              <RESULTS>
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="17244" heatid="19498" lane="0" entrytime="00:02:55.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17202" number="1" />
                    <RELAYPOSITION athleteid="17188" number="2" />
                    <RELAYPOSITION athleteid="17152" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="331" swimtime="00:02:07.96" resultid="17240" heatid="19321" lane="8" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                    <SPLIT distance="100" swimtime="00:01:14.34" />
                    <SPLIT distance="150" swimtime="00:01:41.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17202" number="1" />
                    <RELAYPOSITION athleteid="17152" number="2" reactiontime="+65" />
                    <RELAYPOSITION athleteid="17168" number="3" reactiontime="+192" />
                    <RELAYPOSITION athleteid="17182" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1130" status="DNS" swimtime="00:00:00.00" resultid="17239" heatid="19320" lane="8" entrytime="00:02:39.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17188" number="1" />
                    <RELAYPOSITION athleteid="17214" number="3" />
                    <RELAYPOSITION athleteid="17219" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="9">
              <RESULTS>
                <RESULT eventid="1698" points="296" reactiontime="+104" swimtime="00:02:25.64" resultid="17247" heatid="19563" lane="7" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.67" />
                    <SPLIT distance="100" swimtime="00:01:29.46" />
                    <SPLIT distance="150" swimtime="00:01:59.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17202" number="1" reactiontime="+104" />
                    <RELAYPOSITION athleteid="17152" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="17168" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="17195" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="10">
              <RESULTS>
                <RESULT eventid="1698" status="DNS" swimtime="00:00:00.00" resultid="17248" heatid="19562" lane="0" entrytime="00:02:44.50">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17188" number="2" />
                    <RELAYPOSITION athleteid="17214" number="3" />
                    <RELAYPOSITION athleteid="17219" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="LBS" clubid="14431" name="KP Stilon Gorzów Wlkp.">
          <CONTACT city="Gorzów Wlkp." email="kpstilon@hotmail.com" internet="http://www.kpstilon.gorzow.eu" name="K. Świderski" phone="512 428 265" state="LUB" street="UL. Słowiańska 1/ 42" zip="66-400" />
          <ATHLETES>
            <ATHLETE birthdate="1955-07-15" firstname="Marian" gender="M" lastname="Lasowy" nation="POL" athleteid="14432">
              <RESULTS>
                <RESULT eventid="14207" points="123" reactiontime="+121" swimtime="00:28:20.78" resultid="14433" heatid="19620" lane="1" entrytime="00:29:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.94" />
                    <SPLIT distance="100" swimtime="00:01:42.73" />
                    <SPLIT distance="150" swimtime="00:02:37.46" />
                    <SPLIT distance="200" swimtime="00:03:32.35" />
                    <SPLIT distance="250" swimtime="00:04:27.86" />
                    <SPLIT distance="300" swimtime="00:05:24.24" />
                    <SPLIT distance="350" swimtime="00:06:20.24" />
                    <SPLIT distance="400" swimtime="00:07:17.40" />
                    <SPLIT distance="450" swimtime="00:08:14.28" />
                    <SPLIT distance="500" swimtime="00:09:11.58" />
                    <SPLIT distance="550" swimtime="00:10:08.46" />
                    <SPLIT distance="600" swimtime="00:11:05.81" />
                    <SPLIT distance="650" swimtime="00:12:04.14" />
                    <SPLIT distance="700" swimtime="00:13:01.16" />
                    <SPLIT distance="750" swimtime="00:13:59.07" />
                    <SPLIT distance="800" swimtime="00:14:56.82" />
                    <SPLIT distance="850" swimtime="00:15:54.43" />
                    <SPLIT distance="900" swimtime="00:16:51.80" />
                    <SPLIT distance="950" swimtime="00:17:48.91" />
                    <SPLIT distance="1000" swimtime="00:18:47.59" />
                    <SPLIT distance="1050" swimtime="00:19:45.37" />
                    <SPLIT distance="1100" swimtime="00:20:42.87" />
                    <SPLIT distance="1150" swimtime="00:21:40.52" />
                    <SPLIT distance="1200" swimtime="00:22:37.90" />
                    <SPLIT distance="1250" swimtime="00:23:36.47" />
                    <SPLIT distance="1300" swimtime="00:24:34.97" />
                    <SPLIT distance="1350" swimtime="00:25:32.29" />
                    <SPLIT distance="1400" swimtime="00:26:29.95" />
                    <SPLIT distance="1450" swimtime="00:27:27.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="117" reactiontime="+116" swimtime="00:07:12.84" resultid="14434" heatid="19700" lane="1" entrytime="00:07:26.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.83" />
                    <SPLIT distance="100" swimtime="00:01:40.10" />
                    <SPLIT distance="150" swimtime="00:02:36.20" />
                    <SPLIT distance="200" swimtime="00:03:32.26" />
                    <SPLIT distance="250" swimtime="00:04:28.69" />
                    <SPLIT distance="300" swimtime="00:05:25.28" />
                    <SPLIT distance="350" swimtime="00:06:21.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="14643" name="KS Delfin Gdynia">
          <ATHLETES>
            <ATHLETE birthdate="1971-11-04" firstname="Jakub" gender="M" lastname="Mańczak" nation="POL" athleteid="15037">
              <RESULTS>
                <RESULT eventid="1273" points="369" reactiontime="+81" swimtime="00:01:02.62" resultid="15038" heatid="19384" lane="2" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="260" reactiontime="+79" swimtime="00:02:49.96" resultid="15039" heatid="19417" lane="7" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                    <SPLIT distance="100" swimtime="00:01:20.71" />
                    <SPLIT distance="150" swimtime="00:02:05.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="392" reactiontime="+71" swimtime="00:00:29.77" resultid="15040" heatid="19460" lane="7" entrytime="00:00:29.50" />
                <RESULT eventid="1508" points="329" reactiontime="+78" swimtime="00:02:23.85" resultid="15041" heatid="19493" lane="8" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.53" />
                    <SPLIT distance="100" swimtime="00:01:08.28" />
                    <SPLIT distance="150" swimtime="00:01:46.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="317" reactiontime="+85" swimtime="00:01:10.50" resultid="15042" heatid="19522" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-08-09" firstname="Joanna" gender="F" lastname="Skutkiewicz" nation="POL" athleteid="14644">
              <RESULTS>
                <RESULT eventid="1096" status="WDR" swimtime="00:00:00.00" resultid="14645" entrytime="00:02:53.00" />
                <RESULT eventid="1147" status="WDR" swimtime="00:00:00.00" resultid="14646" entrytime="00:10:55.00" />
                <RESULT eventid="1256" status="WDR" swimtime="00:00:00.00" resultid="14647" entrytime="00:01:10.00" />
                <RESULT eventid="14225" status="WDR" swimtime="00:00:00.00" resultid="14648" entrytime="00:01:20.00" />
                <RESULT eventid="1491" status="WDR" swimtime="00:00:00.00" resultid="14649" entrytime="00:02:55.00" />
                <RESULT eventid="1555" status="WDR" swimtime="00:00:00.00" resultid="14650" entrytime="00:06:05.00" />
                <RESULT eventid="1595" status="WDR" swimtime="00:00:00.00" resultid="14651" entrytime="00:01:33.00" />
                <RESULT eventid="1721" status="WDR" swimtime="00:00:00.00" resultid="14652" entrytime="00:05:20.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="EXOBO" nation="POL" region="WIE" clubid="14740" name="KS Extreme Team Oborniki">
          <CONTACT city="OBORNIKI" email="janwol@poczta.onet.pl" name="WOLNIEWICZ" phone="791064667" state="WIE" street="CZARNKOWSKA 84" zip="64-600" />
          <ATHLETES>
            <ATHLETE birthdate="1948-12-22" firstname="Janusz" gender="M" lastname="Wolniewicz" nation="POL" athleteid="14741">
              <RESULTS>
                <RESULT eventid="1079" points="171" reactiontime="+89" swimtime="00:00:36.45" resultid="14742" heatid="19288" lane="1" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="14207" points="113" reactiontime="+97" swimtime="00:29:10.69" resultid="14743" heatid="19620" lane="7" entrytime="00:29:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.19" />
                    <SPLIT distance="100" swimtime="00:01:40.12" />
                    <SPLIT distance="150" swimtime="00:02:35.75" />
                    <SPLIT distance="200" swimtime="00:03:32.69" />
                    <SPLIT distance="250" swimtime="00:04:29.86" />
                    <SPLIT distance="300" swimtime="00:05:27.08" />
                    <SPLIT distance="350" swimtime="00:06:24.83" />
                    <SPLIT distance="400" swimtime="00:07:22.29" />
                    <SPLIT distance="450" swimtime="00:08:20.73" />
                    <SPLIT distance="500" swimtime="00:09:19.29" />
                    <SPLIT distance="550" swimtime="00:10:17.21" />
                    <SPLIT distance="600" swimtime="00:11:15.12" />
                    <SPLIT distance="650" swimtime="00:12:13.04" />
                    <SPLIT distance="700" swimtime="00:13:11.61" />
                    <SPLIT distance="750" swimtime="00:14:11.91" />
                    <SPLIT distance="800" swimtime="00:15:13.86" />
                    <SPLIT distance="850" swimtime="00:16:11.34" />
                    <SPLIT distance="900" swimtime="00:17:11.39" />
                    <SPLIT distance="950" swimtime="00:18:11.85" />
                    <SPLIT distance="1000" swimtime="00:19:13.28" />
                    <SPLIT distance="1050" swimtime="00:20:14.03" />
                    <SPLIT distance="1100" swimtime="00:21:13.78" />
                    <SPLIT distance="1150" swimtime="00:22:13.81" />
                    <SPLIT distance="1200" swimtime="00:23:14.16" />
                    <SPLIT distance="1250" swimtime="00:24:14.61" />
                    <SPLIT distance="1300" swimtime="00:25:15.99" />
                    <SPLIT distance="1350" swimtime="00:26:15.78" />
                    <SPLIT distance="1400" swimtime="00:27:15.42" />
                    <SPLIT distance="1450" swimtime="00:28:14.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="134" reactiontime="+94" swimtime="00:01:27.81" resultid="14744" heatid="19377" lane="0" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="111" reactiontime="+84" swimtime="00:03:26.27" resultid="14745" heatid="19488" lane="8" entrytime="00:03:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:02:32.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="97" reactiontime="+87" swimtime="00:07:41.63" resultid="14746" heatid="19701" lane="9" entrytime="00:07:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.50" />
                    <SPLIT distance="100" swimtime="00:01:47.18" />
                    <SPLIT distance="150" swimtime="00:02:46.23" />
                    <SPLIT distance="200" swimtime="00:03:46.13" />
                    <SPLIT distance="250" swimtime="00:04:46.74" />
                    <SPLIT distance="300" swimtime="00:05:46.85" />
                    <SPLIT distance="350" swimtime="00:06:47.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KORONAKR" nation="POL" region="KR" clubid="15460" name="KS Korona Kraków">
          <CONTACT city="Kraków" name="Mariola Kuliś" phone="500677133" state="MAŁ" />
          <ATHLETES>
            <ATHLETE birthdate="1966-12-07" firstname="Jarosław" gender="M" lastname="Zadrożny" nation="POL" athleteid="16410">
              <RESULTS>
                <RESULT eventid="1079" points="200" reactiontime="+91" swimtime="00:00:34.62" resultid="16411" heatid="19289" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="14207" points="206" reactiontime="+103" swimtime="00:23:54.36" resultid="16412" heatid="19621" lane="6" entrytime="00:24:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.09" />
                    <SPLIT distance="100" swimtime="00:01:23.16" />
                    <SPLIT distance="150" swimtime="00:02:08.31" />
                    <SPLIT distance="200" swimtime="00:02:54.76" />
                    <SPLIT distance="250" swimtime="00:03:41.75" />
                    <SPLIT distance="300" swimtime="00:04:29.76" />
                    <SPLIT distance="350" swimtime="00:05:17.44" />
                    <SPLIT distance="400" swimtime="00:06:05.09" />
                    <SPLIT distance="450" swimtime="00:06:53.04" />
                    <SPLIT distance="500" swimtime="00:07:41.87" />
                    <SPLIT distance="550" swimtime="00:08:30.20" />
                    <SPLIT distance="600" swimtime="00:09:19.08" />
                    <SPLIT distance="650" swimtime="00:10:07.72" />
                    <SPLIT distance="700" swimtime="00:10:57.03" />
                    <SPLIT distance="750" swimtime="00:11:46.04" />
                    <SPLIT distance="800" swimtime="00:12:35.05" />
                    <SPLIT distance="850" swimtime="00:13:24.29" />
                    <SPLIT distance="900" swimtime="00:14:13.32" />
                    <SPLIT distance="950" swimtime="00:15:02.37" />
                    <SPLIT distance="1000" swimtime="00:15:51.40" />
                    <SPLIT distance="1050" swimtime="00:16:39.91" />
                    <SPLIT distance="1100" swimtime="00:17:28.38" />
                    <SPLIT distance="1150" swimtime="00:18:16.64" />
                    <SPLIT distance="1200" swimtime="00:19:05.62" />
                    <SPLIT distance="1250" swimtime="00:19:54.44" />
                    <SPLIT distance="1300" swimtime="00:20:42.78" />
                    <SPLIT distance="1350" swimtime="00:21:31.88" />
                    <SPLIT distance="1400" swimtime="00:22:20.71" />
                    <SPLIT distance="1450" swimtime="00:23:09.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-03-21" firstname="Janusz" gender="M" lastname="Gołębiowski" nation="POL" athleteid="16383">
              <RESULTS>
                <RESULT eventid="1079" points="28" reactiontime="+112" swimtime="00:01:05.95" resultid="16384" heatid="19284" lane="8" />
                <RESULT eventid="1205" points="11" swimtime="00:01:39.61" resultid="16385" heatid="19342" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-05-16" firstname="Tadeusz" gender="M" lastname="Krawczyk" nation="POL" athleteid="16452">
              <RESULTS>
                <RESULT eventid="1079" points="69" reactiontime="+128" swimtime="00:00:49.20" resultid="16453" heatid="19284" lane="4" entrytime="00:00:46.00" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="16454" heatid="19342" lane="4" entrytime="00:01:10.00" />
                <RESULT eventid="14243" status="DNS" swimtime="00:00:00.00" resultid="16455" heatid="19397" lane="5" entrytime="00:02:30.00" />
                <RESULT eventid="1440" points="17" reactiontime="+124" swimtime="00:01:24.15" resultid="16456" heatid="19450" lane="4" entrytime="00:01:30.00" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="16457" heatid="19486" lane="6" entrytime="00:04:10.00" />
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="16458" heatid="19531" lane="6" entrytime="00:05:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-07-26" firstname="Anna" gender="F" lastname="Koźmin" nation="POL" athleteid="16404">
              <RESULTS>
                <RESULT eventid="1096" points="77" reactiontime="+119" swimtime="00:04:46.19" resultid="16405" heatid="19305" lane="6" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.37" />
                    <SPLIT distance="100" swimtime="00:02:21.69" />
                    <SPLIT distance="150" swimtime="00:03:35.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="89" reactiontime="+124" swimtime="00:02:06.80" resultid="16406" heatid="19390" lane="3" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="104" reactiontime="+126" swimtime="00:02:12.40" resultid="16407" heatid="19428" lane="1" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="82" reactiontime="+121" swimtime="00:00:55.99" resultid="16408" heatid="19445" lane="7" entrytime="00:00:53.00" />
                <RESULT eventid="1664" points="130" reactiontime="+109" swimtime="00:00:56.49" resultid="16409" heatid="19540" lane="9" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-02" firstname="Wojciech" gender="M" lastname="Kaczmarczyk" nation="POL" athleteid="16395">
              <RESULTS>
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="16396" heatid="19359" lane="3" />
                <RESULT eventid="1273" points="63" reactiontime="+106" swimtime="00:01:52.55" resultid="16397" heatid="19374" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-07-29" firstname="Jolanta" gender="F" lastname="Uczarczyk" nation="POL" athleteid="16377">
              <RESULTS>
                <RESULT eventid="1062" points="239" reactiontime="+102" swimtime="00:00:37.43" resultid="16378" heatid="19278" lane="4" entrytime="00:00:37.90" />
                <RESULT eventid="1096" points="170" reactiontime="+77" swimtime="00:03:39.64" resultid="16379" heatid="19305" lane="4" entrytime="00:03:51.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.31" />
                    <SPLIT distance="100" swimtime="00:01:44.31" />
                    <SPLIT distance="150" swimtime="00:02:47.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="188" reactiontime="+118" swimtime="00:01:28.86" resultid="16380" heatid="19369" lane="1" entrytime="00:01:26.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="135" reactiontime="+117" swimtime="00:03:53.11" resultid="16381" heatid="19411" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.77" />
                    <SPLIT distance="100" swimtime="00:01:48.70" />
                    <SPLIT distance="150" swimtime="00:02:50.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="174" reactiontime="+107" swimtime="00:00:43.63" resultid="16382" heatid="19445" lane="4" entrytime="00:00:44.29" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-07-24" firstname="Bogusław" gender="M" lastname="Kwiatkowski" nation="POL" athleteid="16420">
              <RESULTS>
                <RESULT eventid="1079" points="52" reactiontime="+106" swimtime="00:00:54.23" resultid="16421" heatid="19284" lane="7" />
                <RESULT eventid="1205" points="33" reactiontime="+87" swimtime="00:01:09.13" resultid="16422" heatid="19342" lane="8" />
                <RESULT eventid="1239" points="55" reactiontime="+105" swimtime="00:05:15.81" resultid="16423" heatid="19359" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.39" />
                    <SPLIT distance="100" swimtime="00:02:32.42" />
                    <SPLIT distance="150" swimtime="00:03:56.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="53" reactiontime="+104" swimtime="00:02:27.58" resultid="16424" heatid="19433" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="45" reactiontime="+110" swimtime="00:04:37.67" resultid="16425" heatid="19486" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.48" />
                    <SPLIT distance="100" swimtime="00:02:09.77" />
                    <SPLIT distance="150" swimtime="00:03:24.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="34" reactiontime="+96" swimtime="00:05:25.95" resultid="16426" heatid="19530" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.81" />
                    <SPLIT distance="100" swimtime="00:02:34.82" />
                    <SPLIT distance="150" swimtime="00:04:01.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="58" reactiontime="+115" swimtime="00:01:05.08" resultid="16427" heatid="19546" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-21" firstname="Adam" gender="M" lastname="Pycia" nation="POL" athleteid="16473">
              <RESULTS>
                <RESULT eventid="1239" points="222" reactiontime="+98" swimtime="00:03:18.67" resultid="16474" heatid="19360" lane="4" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.58" />
                    <SPLIT distance="100" swimtime="00:01:30.14" />
                    <SPLIT distance="150" swimtime="00:02:23.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="281" reactiontime="+93" swimtime="00:01:08.54" resultid="16475" heatid="19380" lane="8" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="258" reactiontime="+89" swimtime="00:01:27.28" resultid="16476" heatid="19437" lane="5" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="187" reactiontime="+96" swimtime="00:00:38.11" resultid="16477" heatid="19454" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1681" points="273" reactiontime="+98" swimtime="00:00:38.88" resultid="16478" heatid="19554" lane="3" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-06-03" firstname="Antoni" gender="M" lastname="Kubis" nation="POL" athleteid="16413">
              <RESULTS>
                <RESULT comment="G8 - Ukończenie wyścigu nie w położeniu na plecach (Time: 11:49), Z-2" eventid="14243" status="DSQ" swimtime="00:01:49.29" resultid="16414" heatid="19398" lane="7" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="91" reactiontime="+131" swimtime="00:00:55.95" resultid="16415" heatid="19548" lane="7" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-07-17" firstname="Wojciech" gender="M" lastname="Liszkowski" nation="POL" athleteid="16437">
              <RESULTS>
                <RESULT eventid="1205" points="347" reactiontime="+71" swimtime="00:00:31.60" resultid="16438" heatid="19349" lane="2" entrytime="00:00:33.50" />
                <RESULT eventid="1440" points="431" reactiontime="+80" swimtime="00:00:28.86" resultid="16439" heatid="19457" lane="3" entrytime="00:00:31.50" />
                <RESULT eventid="1681" points="381" reactiontime="+93" swimtime="00:00:34.80" resultid="16440" heatid="19553" lane="3" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-10-22" firstname="Maria" gender="F" lastname="Mleczko" nation="POL" athleteid="16338">
              <RESULTS>
                <RESULT eventid="1062" points="47" reactiontime="+120" swimtime="00:01:04.38" resultid="16339" heatid="19275" lane="4" entrytime="00:01:02.00" />
                <RESULT eventid="1096" points="33" reactiontime="+127" swimtime="00:06:18.86" resultid="16340" heatid="19305" lane="7" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:32.94" />
                    <SPLIT distance="100" swimtime="00:03:30.59" />
                    <SPLIT distance="150" swimtime="00:05:02.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="47" reactiontime="+120" swimtime="00:02:20.40" resultid="16341" heatid="19367" lane="2" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="35" reactiontime="+114" swimtime="00:02:52.37" resultid="16342" heatid="19390" lane="9" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:34.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="55" reactiontime="+116" swimtime="00:02:43.69" resultid="16343" heatid="19427" lane="3" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.21" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="(Time: 17:02), Nieprawidłowa praca nóg" eventid="1423" reactiontime="+106" status="DSQ" swimtime="00:01:30.73" resultid="16344" heatid="19445" lane="9" entrytime="00:01:12.00" />
                <RESULT eventid="1595" points="19" reactiontime="+114" swimtime="00:03:22.90" resultid="16345" heatid="19513" lane="8" entrytime="00:03:00.00" />
                <RESULT eventid="1664" points="55" reactiontime="+129" swimtime="00:01:15.07" resultid="16346" heatid="19539" lane="1" entrytime="00:01:08.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-27" firstname="Wacław" gender="M" lastname="Brożek" nation="POL" athleteid="16428">
              <RESULTS>
                <RESULT eventid="1079" points="192" reactiontime="+114" swimtime="00:00:35.09" resultid="16429" heatid="19288" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1113" points="131" reactiontime="+115" swimtime="00:03:35.74" resultid="16430" heatid="19311" lane="1" entrytime="00:03:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.31" />
                    <SPLIT distance="100" swimtime="00:01:50.85" />
                    <SPLIT distance="150" swimtime="00:02:52.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="71" swimtime="00:00:53.57" resultid="16431" heatid="19344" lane="1" entrytime="00:00:53.00" />
                <RESULT eventid="1239" points="131" reactiontime="+115" swimtime="00:03:56.96" resultid="16432" heatid="19359" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.72" />
                    <SPLIT distance="100" swimtime="00:01:59.29" />
                    <SPLIT distance="150" swimtime="00:02:59.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="16433" heatid="19471" lane="4" entrytime="00:02:00.00" />
                <RESULT eventid="1578" points="114" reactiontime="+108" swimtime="00:08:05.55" resultid="16434" heatid="19506" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.73" />
                    <SPLIT distance="100" swimtime="00:02:05.88" />
                    <SPLIT distance="150" swimtime="00:03:12.02" />
                    <SPLIT distance="200" swimtime="00:04:18.68" />
                    <SPLIT distance="250" swimtime="00:05:27.93" />
                    <SPLIT distance="300" swimtime="00:06:35.40" />
                    <SPLIT distance="350" swimtime="00:07:22.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="16435" heatid="19517" lane="5" entrytime="00:01:57.00" />
                <RESULT eventid="1647" points="82" reactiontime="+48" swimtime="00:04:02.66" resultid="16436" heatid="19532" lane="2" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.34" />
                    <SPLIT distance="100" swimtime="00:01:59.69" />
                    <SPLIT distance="150" swimtime="00:03:02.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-07-27" firstname="Mariola" gender="F" lastname="Kuliś" nation="POL" athleteid="16308">
              <RESULTS>
                <RESULT eventid="1062" points="479" reactiontime="+75" swimtime="00:00:29.69" resultid="16309" heatid="19282" lane="4" entrytime="00:00:29.80" />
                <RESULT eventid="1187" points="398" reactiontime="+61" swimtime="00:00:34.88" resultid="16310" heatid="19340" lane="3" entrytime="00:00:35.30" />
                <RESULT eventid="14225" points="417" reactiontime="+71" swimtime="00:01:15.83" resultid="16311" heatid="19395" lane="9" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="424" reactiontime="+73" swimtime="00:00:32.44" resultid="16312" heatid="19448" lane="3" entrytime="00:00:32.70" />
                <RESULT eventid="1457" points="341" reactiontime="+65" swimtime="00:01:18.70" resultid="16313" heatid="19468" lane="6" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="477" reactiontime="+82" swimtime="00:00:36.63" resultid="16314" heatid="19545" lane="2" entrytime="00:00:36.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-09-18" firstname="Izabela" gender="F" lastname="Frączek" nation="POL" athleteid="16459">
              <RESULTS>
                <RESULT eventid="1062" points="507" swimtime="00:00:29.14" resultid="16460" heatid="19283" lane="0" entrytime="00:00:29.00" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1256" points="488" reactiontime="+85" swimtime="00:01:04.66" resultid="16461" heatid="19371" lane="4" entrytime="00:01:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="438" reactiontime="+81" swimtime="00:00:32.10" resultid="16462" heatid="19448" lane="5" entrytime="00:00:32.60" />
                <RESULT eventid="1595" points="375" reactiontime="+80" swimtime="00:01:15.67" resultid="16463" heatid="19515" lane="2" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-07-04" firstname="Stanisław" gender="M" lastname="Waga" nation="POL" athleteid="16441">
              <RESULTS>
                <RESULT eventid="1079" points="76" reactiontime="+111" swimtime="00:00:47.67" resultid="16442" heatid="19285" lane="7" entrytime="00:00:44.00" />
                <RESULT eventid="14207" points="75" reactiontime="+125" swimtime="00:33:27.10" resultid="16443" heatid="19620" lane="8" entrytime="00:42:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.58" />
                    <SPLIT distance="100" swimtime="00:02:04.10" />
                    <SPLIT distance="150" swimtime="00:03:13.80" />
                    <SPLIT distance="200" swimtime="00:04:22.11" />
                    <SPLIT distance="250" swimtime="00:05:28.72" />
                    <SPLIT distance="300" swimtime="00:06:38.94" />
                    <SPLIT distance="350" swimtime="00:07:46.94" />
                    <SPLIT distance="400" swimtime="00:08:53.91" />
                    <SPLIT distance="450" swimtime="00:10:02.29" />
                    <SPLIT distance="500" swimtime="00:11:11.51" />
                    <SPLIT distance="550" swimtime="00:12:17.33" />
                    <SPLIT distance="600" swimtime="00:13:24.76" />
                    <SPLIT distance="650" swimtime="00:14:32.21" />
                    <SPLIT distance="700" swimtime="00:15:38.55" />
                    <SPLIT distance="750" swimtime="00:16:47.48" />
                    <SPLIT distance="800" swimtime="00:17:55.78" />
                    <SPLIT distance="850" swimtime="00:19:03.87" />
                    <SPLIT distance="900" swimtime="00:20:11.38" />
                    <SPLIT distance="950" swimtime="00:21:17.76" />
                    <SPLIT distance="1000" swimtime="00:22:26.69" />
                    <SPLIT distance="1050" swimtime="00:23:33.33" />
                    <SPLIT distance="1100" swimtime="00:24:39.66" />
                    <SPLIT distance="1150" swimtime="00:25:46.62" />
                    <SPLIT distance="1200" swimtime="00:26:52.66" />
                    <SPLIT distance="1250" swimtime="00:27:59.05" />
                    <SPLIT distance="1300" swimtime="00:29:05.49" />
                    <SPLIT distance="1350" swimtime="00:30:12.55" />
                    <SPLIT distance="1400" swimtime="00:31:18.46" />
                    <SPLIT distance="1450" swimtime="00:32:25.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="68" reactiontime="+109" swimtime="00:01:49.57" resultid="16444" heatid="19375" lane="0" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="64" reactiontime="+119" swimtime="00:04:08.00" resultid="16445" heatid="19487" lane="9" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.95" />
                    <SPLIT distance="100" swimtime="00:01:55.86" />
                    <SPLIT distance="150" swimtime="00:03:02.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="59" reactiontime="+116" swimtime="00:01:04.54" resultid="16446" heatid="19547" lane="6" entrytime="00:01:02.00" />
                <RESULT eventid="1744" points="64" reactiontime="+121" swimtime="00:08:49.18" resultid="16447" heatid="19699" lane="5" entrytime="00:08:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.05" />
                    <SPLIT distance="100" swimtime="00:02:04.63" />
                    <SPLIT distance="150" swimtime="00:03:13.83" />
                    <SPLIT distance="200" swimtime="00:04:23.39" />
                    <SPLIT distance="250" swimtime="00:05:31.74" />
                    <SPLIT distance="300" swimtime="00:06:40.25" />
                    <SPLIT distance="350" swimtime="00:07:46.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-21" firstname="Klaudia" gender="F" lastname="Wysocka" nation="POL" athleteid="16398">
              <RESULTS>
                <RESULT eventid="1096" points="295" reactiontime="+86" swimtime="00:03:02.89" resultid="16399" heatid="19307" lane="7" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.51" />
                    <SPLIT distance="100" swimtime="00:01:26.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="313" reactiontime="+84" swimtime="00:01:23.38" resultid="16400" heatid="19393" lane="7" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="267" reactiontime="+101" swimtime="00:01:36.75" resultid="16401" heatid="19430" lane="0" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="273" reactiontime="+106" swimtime="00:06:39.62" resultid="16402" heatid="19504" lane="2" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.25" />
                    <SPLIT distance="100" swimtime="00:01:26.71" />
                    <SPLIT distance="150" swimtime="00:02:19.92" />
                    <SPLIT distance="250" swimtime="00:04:09.46" />
                    <SPLIT distance="300" swimtime="00:05:07.96" />
                    <SPLIT distance="350" swimtime="00:05:54.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="278" reactiontime="+85" swimtime="00:01:23.58" resultid="16403" heatid="19515" lane="9" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-10-20" firstname="Janusz" gender="M" lastname="Toporski" nation="POL" athleteid="16320">
              <RESULTS>
                <RESULT eventid="1079" points="117" reactiontime="+100" swimtime="00:00:41.42" resultid="16321" heatid="19284" lane="3" entrytime="00:00:50.00" />
                <RESULT eventid="1113" points="120" reactiontime="+103" swimtime="00:03:41.68" resultid="16322" heatid="19310" lane="4" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.16" />
                    <SPLIT distance="100" swimtime="00:01:55.07" />
                    <SPLIT distance="150" swimtime="00:02:51.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="160" reactiontime="+105" swimtime="00:03:41.42" resultid="16323" heatid="19360" lane="2" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.24" />
                    <SPLIT distance="100" swimtime="00:01:49.61" />
                    <SPLIT distance="150" swimtime="00:02:46.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="112" reactiontime="+89" swimtime="00:01:44.32" resultid="16324" heatid="19398" lane="8" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="148" reactiontime="+87" swimtime="00:01:45.04" resultid="16325" heatid="19434" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="100" reactiontime="+95" swimtime="00:00:46.95" resultid="16326" heatid="19451" lane="0" entrytime="00:01:00.00" />
                <RESULT eventid="1681" points="134" reactiontime="+85" swimtime="00:00:49.32" resultid="16327" heatid="19547" lane="3" entrytime="00:01:00.00" />
                <RESULT eventid="1744" points="115" reactiontime="+95" swimtime="00:07:16.23" resultid="16328" heatid="19700" lane="9" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.69" />
                    <SPLIT distance="100" swimtime="00:01:44.59" />
                    <SPLIT distance="150" swimtime="00:02:40.78" />
                    <SPLIT distance="200" swimtime="00:03:36.54" />
                    <SPLIT distance="250" swimtime="00:04:33.04" />
                    <SPLIT distance="300" swimtime="00:05:29.59" />
                    <SPLIT distance="350" swimtime="00:06:25.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-09-15" firstname="Mirosława" gender="F" lastname="Legutko" nation="POL" athleteid="16386">
              <RESULTS>
                <RESULT eventid="1062" points="243" swimtime="00:00:37.21" resultid="16387" heatid="19279" lane="0" entrytime="00:00:37.00" />
                <RESULT eventid="1147" points="148" reactiontime="+109" swimtime="00:15:05.27" resultid="16388" heatid="19595" lane="9" entrytime="00:15:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.97" />
                    <SPLIT distance="100" swimtime="00:01:43.70" />
                    <SPLIT distance="150" swimtime="00:02:41.76" />
                    <SPLIT distance="200" swimtime="00:03:40.03" />
                    <SPLIT distance="250" swimtime="00:04:36.84" />
                    <SPLIT distance="300" swimtime="00:05:34.69" />
                    <SPLIT distance="350" swimtime="00:06:32.57" />
                    <SPLIT distance="400" swimtime="00:07:30.31" />
                    <SPLIT distance="450" swimtime="00:08:27.46" />
                    <SPLIT distance="500" swimtime="00:09:26.16" />
                    <SPLIT distance="550" swimtime="00:10:23.17" />
                    <SPLIT distance="600" swimtime="00:11:20.96" />
                    <SPLIT distance="650" swimtime="00:13:14.15" />
                    <SPLIT distance="700" swimtime="00:14:11.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="171" reactiontime="+110" swimtime="00:01:31.57" resultid="16389" heatid="19367" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:31.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="116" reactiontime="+113" swimtime="00:04:04.62" resultid="16390" heatid="19412" lane="9" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.51" />
                    <SPLIT distance="100" swimtime="00:01:56.58" />
                    <SPLIT distance="150" swimtime="00:03:00.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="165" reactiontime="+109" swimtime="00:00:44.39" resultid="16391" heatid="19445" lane="5" entrytime="00:00:45.00" />
                <RESULT eventid="1555" points="144" reactiontime="+112" swimtime="00:08:14.53" resultid="16392" heatid="19503" lane="5" entrytime="00:08:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.63" />
                    <SPLIT distance="100" swimtime="00:02:01.13" />
                    <SPLIT distance="150" swimtime="00:03:04.18" />
                    <SPLIT distance="200" swimtime="00:04:09.08" />
                    <SPLIT distance="250" swimtime="00:05:17.83" />
                    <SPLIT distance="300" swimtime="00:06:25.80" />
                    <SPLIT distance="350" swimtime="00:07:21.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="116" reactiontime="+112" swimtime="00:01:51.90" resultid="16393" heatid="19513" lane="6" entrytime="00:01:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="159" reactiontime="+112" swimtime="00:07:12.35" resultid="16394" heatid="19695" lane="5" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.29" />
                    <SPLIT distance="100" swimtime="00:01:42.05" />
                    <SPLIT distance="150" swimtime="00:02:38.05" />
                    <SPLIT distance="200" swimtime="00:03:33.85" />
                    <SPLIT distance="250" swimtime="00:04:29.79" />
                    <SPLIT distance="300" swimtime="00:05:26.67" />
                    <SPLIT distance="350" swimtime="00:06:22.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-30" firstname="Piotr" gender="M" lastname="Łysiak" nation="POL" athleteid="16315">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="16316" heatid="19294" lane="6" entrytime="00:00:29.06" />
                <RESULT eventid="1239" points="339" reactiontime="+85" swimtime="00:02:52.73" resultid="16317" heatid="19364" lane="9" entrytime="00:02:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.77" />
                    <SPLIT distance="100" swimtime="00:01:21.60" />
                    <SPLIT distance="150" swimtime="00:02:05.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="343" reactiontime="+96" swimtime="00:01:19.42" resultid="16318" heatid="19440" lane="2" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="16319" heatid="19555" lane="8" entrytime="00:00:36.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-05-29" firstname="Małgorzata" gender="F" lastname="Orlewicz-Musiał" nation="POL" athleteid="16347">
              <RESULTS>
                <RESULT eventid="1062" points="109" reactiontime="+107" swimtime="00:00:48.55" resultid="16348" heatid="19276" lane="4" entrytime="00:00:45.90" />
                <RESULT eventid="1147" reactiontime="+111" status="OTL" swimtime="00:00:00.00" resultid="16349" heatid="19595" lane="1" entrytime="00:15:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.90" />
                    <SPLIT distance="100" swimtime="00:01:55.51" />
                    <SPLIT distance="150" swimtime="00:02:59.94" />
                    <SPLIT distance="200" swimtime="00:04:04.13" />
                    <SPLIT distance="250" swimtime="00:05:09.81" />
                    <SPLIT distance="300" swimtime="00:06:16.98" />
                    <SPLIT distance="350" swimtime="00:07:22.99" />
                    <SPLIT distance="400" swimtime="00:08:28.84" />
                    <SPLIT distance="450" swimtime="00:09:35.52" />
                    <SPLIT distance="500" swimtime="00:10:41.92" />
                    <SPLIT distance="550" swimtime="00:11:50.84" />
                    <SPLIT distance="600" swimtime="00:12:56.32" />
                    <SPLIT distance="650" swimtime="00:14:01.09" />
                    <SPLIT distance="700" swimtime="00:15:06.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="63" swimtime="00:01:04.46" resultid="16350" heatid="19336" lane="6" entrytime="00:01:01.52" />
                <RESULT eventid="1324" status="DNS" swimtime="00:00:00.00" resultid="16351" heatid="19411" lane="6" entrytime="00:04:49.79" />
                <RESULT eventid="1457" points="51" swimtime="00:02:28.25" resultid="16352" heatid="19465" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="102" reactiontime="+106" swimtime="00:03:57.08" resultid="16353" heatid="19480" lane="1" entrytime="00:03:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.46" />
                    <SPLIT distance="100" swimtime="00:01:52.13" />
                    <SPLIT distance="150" swimtime="00:02:56.75" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="M12 - Niejednoczesne dotknięcie ściany dłońmi przy nawrocie lub na zakończenie wyścigu (Time: 9:07)" eventid="1595" reactiontime="+113" status="DSQ" swimtime="00:02:25.12" resultid="16354" heatid="19513" lane="1" entrytime="00:02:13.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="95" reactiontime="+113" swimtime="00:08:33.66" resultid="16355" heatid="19695" lane="6" entrytime="00:08:16.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.74" />
                    <SPLIT distance="100" swimtime="00:01:57.08" />
                    <SPLIT distance="150" swimtime="00:03:02.37" />
                    <SPLIT distance="200" swimtime="00:04:07.69" />
                    <SPLIT distance="250" swimtime="00:05:15.78" />
                    <SPLIT distance="300" swimtime="00:06:22.46" />
                    <SPLIT distance="350" swimtime="00:07:28.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-04-20" firstname="Agnieszka" gender="F" lastname="Macierzewska" nation="POL" athleteid="16464">
              <RESULTS>
                <RESULT eventid="1062" points="309" swimtime="00:00:34.35" resultid="16465" heatid="19280" lane="9" entrytime="00:00:34.00" />
                <RESULT eventid="1147" points="270" reactiontime="+111" swimtime="00:12:21.49" resultid="16466" heatid="19595" lane="5" entrytime="00:12:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.25" />
                    <SPLIT distance="100" swimtime="00:01:23.11" />
                    <SPLIT distance="150" swimtime="00:02:09.52" />
                    <SPLIT distance="200" swimtime="00:02:56.32" />
                    <SPLIT distance="250" swimtime="00:03:43.66" />
                    <SPLIT distance="300" swimtime="00:04:31.19" />
                    <SPLIT distance="350" swimtime="00:05:18.65" />
                    <SPLIT distance="400" swimtime="00:06:05.99" />
                    <SPLIT distance="450" swimtime="00:06:53.30" />
                    <SPLIT distance="500" swimtime="00:07:40.57" />
                    <SPLIT distance="550" swimtime="00:08:28.03" />
                    <SPLIT distance="600" swimtime="00:09:15.95" />
                    <SPLIT distance="650" swimtime="00:10:03.00" />
                    <SPLIT distance="700" swimtime="00:10:50.71" />
                    <SPLIT distance="750" swimtime="00:11:37.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="299" reactiontime="+95" swimtime="00:01:16.06" resultid="16467" heatid="19370" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="210" reactiontime="+104" swimtime="00:03:20.95" resultid="16468" heatid="19412" lane="8" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.41" />
                    <SPLIT distance="100" swimtime="00:01:33.70" />
                    <SPLIT distance="150" swimtime="00:02:27.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="258" reactiontime="+96" swimtime="00:00:38.28" resultid="16469" heatid="19446" lane="5" entrytime="00:00:39.00" />
                <RESULT eventid="1555" points="232" reactiontime="+104" swimtime="00:07:02.24" resultid="16470" heatid="19504" lane="1" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.17" />
                    <SPLIT distance="150" swimtime="00:02:33.32" />
                    <SPLIT distance="200" swimtime="00:03:27.51" />
                    <SPLIT distance="250" swimtime="00:04:28.26" />
                    <SPLIT distance="300" swimtime="00:05:29.22" />
                    <SPLIT distance="350" swimtime="00:06:17.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="224" swimtime="00:01:29.82" resultid="16471" heatid="19514" lane="0" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="268" reactiontime="+102" swimtime="00:06:03.55" resultid="16472" heatid="19697" lane="3" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.03" />
                    <SPLIT distance="100" swimtime="00:01:25.11" />
                    <SPLIT distance="150" swimtime="00:02:11.32" />
                    <SPLIT distance="200" swimtime="00:02:57.73" />
                    <SPLIT distance="250" swimtime="00:03:45.09" />
                    <SPLIT distance="300" swimtime="00:04:32.56" />
                    <SPLIT distance="350" swimtime="00:05:19.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-02-18" firstname="Bartosz" gender="M" lastname="Próchniewicz" nation="POL" athleteid="16356">
              <RESULTS>
                <RESULT eventid="1205" points="92" reactiontime="+89" swimtime="00:00:49.21" resultid="16357" heatid="19344" lane="6" entrytime="00:00:50.00" />
                <RESULT eventid="14243" points="96" reactiontime="+88" swimtime="00:01:49.72" resultid="16358" heatid="19398" lane="3" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="80" swimtime="00:01:53.23" resultid="16359" heatid="19472" lane="8" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="16360" heatid="19547" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-11-10" firstname="Waldemar" gender="M" lastname="Piszczek" nation="POL" athleteid="16361">
              <RESULTS>
                <RESULT eventid="1079" points="296" reactiontime="+84" swimtime="00:00:30.39" resultid="16362" heatid="19292" lane="9" entrytime="00:00:31.00" />
                <RESULT eventid="1205" points="254" reactiontime="+74" swimtime="00:00:35.08" resultid="16363" heatid="19348" lane="9" entrytime="00:00:36.00" />
                <RESULT eventid="14243" points="295" reactiontime="+94" swimtime="00:01:15.54" resultid="16364" heatid="19403" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="334" reactiontime="+89" swimtime="00:00:31.42" resultid="16365" heatid="19457" lane="7" entrytime="00:00:32.00" />
                <RESULT eventid="1474" points="227" reactiontime="+77" swimtime="00:01:20.08" resultid="16366" heatid="19475" lane="9" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="266" reactiontime="+103" swimtime="00:01:14.68" resultid="16367" heatid="19520" lane="6" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="312" reactiontime="+104" swimtime="00:00:37.21" resultid="16368" heatid="19553" lane="1" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-08-26" firstname="Andrzej" gender="M" lastname="Mleczko" nation="POL" athleteid="16329">
              <RESULTS>
                <RESULT eventid="1113" points="119" reactiontime="+129" swimtime="00:03:42.40" resultid="16330" heatid="19311" lane="2" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.24" />
                    <SPLIT distance="100" swimtime="00:01:47.32" />
                    <SPLIT distance="150" swimtime="00:02:54.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14207" points="136" reactiontime="+145" swimtime="00:27:25.35" resultid="16331" heatid="19620" lane="2" entrytime="00:26:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.77" />
                    <SPLIT distance="100" swimtime="00:01:43.30" />
                    <SPLIT distance="150" swimtime="00:02:37.64" />
                    <SPLIT distance="200" swimtime="00:03:32.10" />
                    <SPLIT distance="250" swimtime="00:04:28.20" />
                    <SPLIT distance="300" swimtime="00:05:24.14" />
                    <SPLIT distance="350" swimtime="00:06:20.50" />
                    <SPLIT distance="400" swimtime="00:07:16.49" />
                    <SPLIT distance="450" swimtime="00:08:11.52" />
                    <SPLIT distance="500" swimtime="00:09:05.71" />
                    <SPLIT distance="550" swimtime="00:10:01.31" />
                    <SPLIT distance="600" swimtime="00:10:56.15" />
                    <SPLIT distance="650" swimtime="00:11:51.80" />
                    <SPLIT distance="700" swimtime="00:12:47.29" />
                    <SPLIT distance="750" swimtime="00:13:42.11" />
                    <SPLIT distance="800" swimtime="00:14:37.42" />
                    <SPLIT distance="850" swimtime="00:15:32.95" />
                    <SPLIT distance="900" swimtime="00:16:28.83" />
                    <SPLIT distance="950" swimtime="00:17:24.10" />
                    <SPLIT distance="1000" swimtime="00:18:19.74" />
                    <SPLIT distance="1050" swimtime="00:19:15.40" />
                    <SPLIT distance="1100" swimtime="00:20:10.72" />
                    <SPLIT distance="1150" swimtime="00:21:06.57" />
                    <SPLIT distance="1200" swimtime="00:22:01.43" />
                    <SPLIT distance="1250" swimtime="00:22:55.79" />
                    <SPLIT distance="1300" swimtime="00:23:50.99" />
                    <SPLIT distance="1350" swimtime="00:24:46.49" />
                    <SPLIT distance="1400" swimtime="00:25:43.13" />
                    <SPLIT distance="1450" swimtime="00:26:38.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="200" reactiontime="+131" swimtime="00:01:16.77" resultid="16332" heatid="19378" lane="1" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="131" reactiontime="+122" swimtime="00:01:38.86" resultid="16333" heatid="19399" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="165" reactiontime="+128" swimtime="00:03:00.84" resultid="16334" heatid="19488" lane="3" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.77" />
                    <SPLIT distance="100" swimtime="00:01:27.50" />
                    <SPLIT distance="150" swimtime="00:02:13.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="91" reactiontime="+135" swimtime="00:08:42.82" resultid="16335" heatid="19507" lane="5" entrytime="00:08:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.49" />
                    <SPLIT distance="100" swimtime="00:02:03.34" />
                    <SPLIT distance="150" swimtime="00:03:16.90" />
                    <SPLIT distance="200" swimtime="00:04:30.14" />
                    <SPLIT distance="250" swimtime="00:05:43.17" />
                    <SPLIT distance="300" swimtime="00:06:55.52" />
                    <SPLIT distance="350" swimtime="00:07:56.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="78" reactiontime="+142" swimtime="00:01:52.22" resultid="16336" heatid="19518" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="141" reactiontime="+141" swimtime="00:06:47.26" resultid="16337" heatid="19701" lane="2" entrytime="00:06:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.81" />
                    <SPLIT distance="100" swimtime="00:01:38.66" />
                    <SPLIT distance="150" swimtime="00:02:30.36" />
                    <SPLIT distance="200" swimtime="00:03:22.62" />
                    <SPLIT distance="250" swimtime="00:04:13.84" />
                    <SPLIT distance="300" swimtime="00:05:05.78" />
                    <SPLIT distance="350" swimtime="00:05:56.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-02-08" firstname="Tomasz" gender="M" lastname="Czerniecki" nation="POL" athleteid="16416">
              <RESULTS>
                <RESULT eventid="1079" points="470" reactiontime="+72" swimtime="00:00:26.05" resultid="16417" heatid="19301" lane="6" entrytime="00:00:26.00" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="16418" heatid="19373" lane="3" />
                <RESULT eventid="14243" points="411" reactiontime="+81" swimtime="00:01:07.62" resultid="16419" heatid="19408" lane="1" entrytime="00:01:07.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-12-23" firstname="Anna" gender="F" lastname="Janeczko" nation="POL" athleteid="16369">
              <RESULTS>
                <RESULT eventid="1062" points="314" reactiontime="+97" swimtime="00:00:34.18" resultid="16370" heatid="19280" lane="3" entrytime="00:00:33.20" />
                <RESULT eventid="1187" points="242" reactiontime="+84" swimtime="00:00:41.15" resultid="16371" heatid="19338" lane="6" entrytime="00:00:42.00" />
                <RESULT eventid="1256" points="282" reactiontime="+104" swimtime="00:01:17.58" resultid="16372" heatid="19369" lane="4" entrytime="00:01:19.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="251" reactiontime="+98" swimtime="00:00:38.61" resultid="16373" heatid="19447" lane="2" entrytime="00:00:36.50" />
                <RESULT eventid="1555" points="214" reactiontime="+101" swimtime="00:07:13.77" resultid="16374" heatid="19504" lane="9" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.40" />
                    <SPLIT distance="100" swimtime="00:01:47.54" />
                    <SPLIT distance="150" swimtime="00:02:41.91" />
                    <SPLIT distance="200" swimtime="00:03:35.34" />
                    <SPLIT distance="250" swimtime="00:04:38.20" />
                    <SPLIT distance="300" swimtime="00:05:39.60" />
                    <SPLIT distance="350" swimtime="00:06:28.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="145" reactiontime="+105" swimtime="00:01:43.76" resultid="16375" heatid="19513" lane="3" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="196" reactiontime="+89" swimtime="00:03:25.12" resultid="16376" heatid="19527" lane="6" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.14" />
                    <SPLIT distance="100" swimtime="00:01:41.73" />
                    <SPLIT distance="150" swimtime="00:02:36.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-03-26" firstname="Józef" gender="M" lastname="Śmigielski" nation="POL" athleteid="16448">
              <RESULTS>
                <RESULT eventid="1205" points="49" reactiontime="+100" swimtime="00:01:00.66" resultid="16449" heatid="19343" lane="8" entrytime="00:01:00.00" />
                <RESULT eventid="1474" points="55" reactiontime="+98" swimtime="00:02:08.58" resultid="16450" heatid="19471" lane="1" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="52" reactiontime="+106" swimtime="00:04:42.14" resultid="16451" heatid="19532" lane="8" entrytime="00:04:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.17" />
                    <SPLIT distance="100" swimtime="00:02:16.65" />
                    <SPLIT distance="150" swimtime="00:03:31.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Korona Kraków C" number="6">
              <RESULTS>
                <RESULT eventid="1381" points="376" reactiontime="+67" swimtime="00:02:05.38" resultid="16484" heatid="19423" lane="5" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.91" />
                    <SPLIT distance="100" swimtime="00:01:08.11" />
                    <SPLIT distance="150" swimtime="00:01:39.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16437" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="16315" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="16361" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="16416" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" name="Korona Kraków E" number="7">
              <RESULTS>
                <RESULT eventid="1381" points="85" reactiontime="+89" swimtime="00:03:25.48" resultid="16485" heatid="19421" lane="2" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.18" />
                    <SPLIT distance="100" swimtime="00:01:58.20" />
                    <SPLIT distance="150" swimtime="00:02:40.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16420" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="16320" number="2" reactiontime="+6" />
                    <RELAYPOSITION athleteid="16473" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="16452" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" name="Korona Kraków F" number="8">
              <RESULTS>
                <RESULT eventid="1381" points="77" reactiontime="+107" swimtime="00:03:31.89" resultid="16486" heatid="19421" lane="1" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.53" />
                    <SPLIT distance="100" swimtime="00:02:57.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16448" number="1" reactiontime="+107" />
                    <RELAYPOSITION athleteid="16441" number="2" reactiontime="+94" />
                    <RELAYPOSITION athleteid="16413" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="16329" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" name="Korona Kraków E" number="11">
              <RESULTS>
                <RESULT eventid="1548" points="236" reactiontime="+92" swimtime="00:02:13.66" resultid="16489" heatid="19500" lane="7" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.19" />
                    <SPLIT distance="100" swimtime="00:01:11.33" />
                    <SPLIT distance="150" swimtime="00:01:45.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16361" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="16413" number="2" reactiontime="+81" />
                    <RELAYPOSITION athleteid="16329" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="16437" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" name="Korona Kraków F" number="12">
              <RESULTS>
                <RESULT eventid="1548" points="86" reactiontime="+138" swimtime="00:03:07.04" resultid="16490" heatid="19499" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.98" />
                    <SPLIT distance="150" swimtime="00:02:29.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16448" number="1" reactiontime="+138" />
                    <RELAYPOSITION athleteid="16441" number="2" reactiontime="+14" />
                    <RELAYPOSITION athleteid="16452" number="3" />
                    <RELAYPOSITION athleteid="16320" number="4" reactiontime="+20" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="Korona Kraków D" number="4">
              <RESULTS>
                <RESULT eventid="1358" points="376" reactiontime="+82" swimtime="00:02:23.06" resultid="16482" heatid="19420" lane="6" entrytime="00:02:22.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.21" />
                    <SPLIT distance="100" swimtime="00:01:18.91" />
                    <SPLIT distance="150" swimtime="00:01:54.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16464" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="16308" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="16398" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="16459" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="F" name="Korona Kraków E" number="5">
              <RESULTS>
                <RESULT eventid="1358" points="125" reactiontime="+97" swimtime="00:03:26.20" resultid="16483" heatid="19420" lane="0" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.38" />
                    <SPLIT distance="100" swimtime="00:01:56.29" />
                    <SPLIT distance="150" swimtime="00:02:34.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16386" number="1" reactiontime="+97" />
                    <RELAYPOSITION athleteid="16338" number="2" reactiontime="+68" />
                    <RELAYPOSITION athleteid="16369" number="3" reactiontime="+91" />
                    <RELAYPOSITION athleteid="16404" number="4" reactiontime="+89" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="Korona Kraków D" number="9">
              <RESULTS>
                <RESULT eventid="1525" points="408" reactiontime="+78" swimtime="00:02:06.99" resultid="16487" heatid="19498" lane="5" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                    <SPLIT distance="100" swimtime="00:01:04.94" />
                    <SPLIT distance="150" swimtime="00:01:38.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16308" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="16464" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="16369" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="16459" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="F" name="Korona Kraków E" number="10">
              <RESULTS>
                <RESULT eventid="1525" points="107" reactiontime="+122" swimtime="00:03:18.30" resultid="16488" heatid="19497" lane="4" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.38" />
                    <SPLIT distance="100" swimtime="00:02:02.82" />
                    <SPLIT distance="150" swimtime="00:02:42.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16404" number="1" reactiontime="+122" />
                    <RELAYPOSITION athleteid="16338" number="2" reactiontime="+90" />
                    <RELAYPOSITION athleteid="16386" number="3" reactiontime="+74" />
                    <RELAYPOSITION athleteid="16398" number="4" reactiontime="+62" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Korona Kraków D" number="1">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1130" points="418" reactiontime="+83" swimtime="00:01:58.44" resultid="16479" heatid="19322" lane="0" entrytime="00:01:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.91" />
                    <SPLIT distance="100" swimtime="00:01:04.20" />
                    <SPLIT distance="150" swimtime="00:01:32.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16308" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="16329" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="16459" number="3" reactiontime="+18" />
                    <RELAYPOSITION athleteid="16416" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" name="Korona Kraków E" number="2">
              <RESULTS>
                <RESULT eventid="1130" points="223" reactiontime="+92" swimtime="00:02:25.93" resultid="16480" heatid="19320" lane="6" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.47" />
                    <SPLIT distance="100" swimtime="00:01:08.43" />
                    <SPLIT distance="150" swimtime="00:01:51.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16361" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="16386" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="16413" number="3" reactiontime="+95" />
                    <RELAYPOSITION athleteid="16464" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" name="Korona Kraków F" number="3">
              <RESULTS>
                <RESULT eventid="1130" points="69" reactiontime="+112" swimtime="00:03:35.43" resultid="16481" heatid="19319" lane="5" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.91" />
                    <SPLIT distance="100" swimtime="00:01:56.41" />
                    <SPLIT distance="150" swimtime="00:02:43.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16338" number="1" reactiontime="+112" />
                    <RELAYPOSITION athleteid="16452" number="2" reactiontime="+84" />
                    <RELAYPOSITION athleteid="16441" number="3" reactiontime="+24" />
                    <RELAYPOSITION athleteid="16404" number="4" reactiontime="+104" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="Korona Kraków C" number="13">
              <RESULTS>
                <RESULT eventid="1698" points="433" reactiontime="+70" swimtime="00:02:08.38" resultid="16491" heatid="19564" lane="2" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                    <SPLIT distance="100" swimtime="00:01:11.37" />
                    <SPLIT distance="150" swimtime="00:01:40.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16308" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="16315" number="2" reactiontime="+27" />
                    <RELAYPOSITION athleteid="16437" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="16459" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" name="Korona Kraków E" number="14">
              <RESULTS>
                <RESULT eventid="1698" points="248" reactiontime="+80" swimtime="00:02:34.65" resultid="16492" heatid="19562" lane="7" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.29" />
                    <SPLIT distance="100" swimtime="00:01:20.76" />
                    <SPLIT distance="150" swimtime="00:02:00.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16386" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="16361" number="2" reactiontime="+33" />
                    <RELAYPOSITION athleteid="16464" number="3" reactiontime="+60" />
                    <RELAYPOSITION athleteid="16329" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" name="Korona Kraków F" number="15">
              <RESULTS>
                <RESULT eventid="1698" points="70" reactiontime="+109" swimtime="00:03:55.26" resultid="16493" heatid="19562" lane="3" entrytime="00:03:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.26" />
                    <SPLIT distance="100" swimtime="00:02:11.73" />
                    <SPLIT distance="150" swimtime="00:03:08.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16413" number="1" reactiontime="+109" />
                    <RELAYPOSITION athleteid="16338" number="2" />
                    <RELAYPOSITION athleteid="16404" number="3" reactiontime="+102" />
                    <RELAYPOSITION athleteid="16441" number="4" reactiontime="+18" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02001" nation="POL" region="DOL" clubid="18064" name="KS Rekin Świebodzice">
          <CONTACT city="Świebodzice" email="winiar182@wp.pl" internet="www.klubrekin.pl" name="WINIARCZYK Krzysztof" phone="606626274" state="DOL" street="Mieszka Starego 4" zip="58-160" />
          <ATHLETES>
            <ATHLETE birthdate="1984-12-12" firstname="Karolina" gender="F" lastname="Jahnz" nation="POL" athleteid="18359">
              <RESULTS>
                <RESULT eventid="1096" points="374" reactiontime="+74" swimtime="00:02:49.02" resultid="18360" heatid="19305" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                    <SPLIT distance="100" swimtime="00:01:20.59" />
                    <SPLIT distance="150" swimtime="00:02:09.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="395" reactiontime="+82" swimtime="00:10:52.92" resultid="18361" heatid="19595" lane="4" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                    <SPLIT distance="100" swimtime="00:01:14.71" />
                    <SPLIT distance="150" swimtime="00:01:55.74" />
                    <SPLIT distance="200" swimtime="00:02:36.52" />
                    <SPLIT distance="250" swimtime="00:03:18.17" />
                    <SPLIT distance="300" swimtime="00:03:59.95" />
                    <SPLIT distance="350" swimtime="00:04:41.60" />
                    <SPLIT distance="400" swimtime="00:05:23.59" />
                    <SPLIT distance="450" swimtime="00:06:06.17" />
                    <SPLIT distance="500" swimtime="00:06:48.44" />
                    <SPLIT distance="550" swimtime="00:07:29.85" />
                    <SPLIT distance="600" swimtime="00:08:11.22" />
                    <SPLIT distance="650" swimtime="00:08:52.88" />
                    <SPLIT distance="700" swimtime="00:09:33.95" />
                    <SPLIT distance="750" swimtime="00:10:14.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="390" reactiontime="+83" swimtime="00:03:04.12" resultid="18362" heatid="19357" lane="2" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.99" />
                    <SPLIT distance="100" swimtime="00:01:29.24" />
                    <SPLIT distance="150" swimtime="00:02:16.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="285" reactiontime="+81" swimtime="00:03:01.60" resultid="18363" heatid="19412" lane="3" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                    <SPLIT distance="100" swimtime="00:01:24.33" />
                    <SPLIT distance="150" swimtime="00:02:13.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="395" reactiontime="+85" swimtime="00:02:30.86" resultid="18364" heatid="19479" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                    <SPLIT distance="100" swimtime="00:01:11.90" />
                    <SPLIT distance="150" swimtime="00:01:52.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="375" reactiontime="+84" swimtime="00:05:59.48" resultid="18365" heatid="19505" lane="0" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.30" />
                    <SPLIT distance="100" swimtime="00:01:26.30" />
                    <SPLIT distance="150" swimtime="00:02:13.35" />
                    <SPLIT distance="200" swimtime="00:02:59.30" />
                    <SPLIT distance="250" swimtime="00:03:49.06" />
                    <SPLIT distance="300" swimtime="00:04:39.68" />
                    <SPLIT distance="350" swimtime="00:05:20.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="310" reactiontime="+82" swimtime="00:02:56.03" resultid="18366" heatid="19526" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.57" />
                    <SPLIT distance="100" swimtime="00:01:24.60" />
                    <SPLIT distance="150" swimtime="00:02:10.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="392" reactiontime="+67" swimtime="00:05:20.42" resultid="18367" heatid="19698" lane="0" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                    <SPLIT distance="100" swimtime="00:01:16.15" />
                    <SPLIT distance="150" swimtime="00:01:56.97" />
                    <SPLIT distance="200" swimtime="00:02:37.91" />
                    <SPLIT distance="250" swimtime="00:03:19.92" />
                    <SPLIT distance="300" swimtime="00:04:00.83" />
                    <SPLIT distance="350" swimtime="00:04:41.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-06-21" firstname="Alfred" gender="M" lastname="Żemier" nation="POL" athleteid="18385">
              <RESULTS>
                <RESULT eventid="1079" points="484" reactiontime="+66" swimtime="00:00:25.80" resultid="18386" heatid="19303" lane="9" entrytime="00:00:25.00" />
                <RESULT eventid="1113" points="330" reactiontime="+71" swimtime="00:02:38.64" resultid="18387" heatid="19317" lane="8" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.49" />
                    <SPLIT distance="100" swimtime="00:01:12.33" />
                    <SPLIT distance="150" swimtime="00:01:58.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="406" reactiontime="+72" swimtime="00:00:29.99" resultid="18388" heatid="19351" lane="0" entrytime="00:00:31.00" />
                <RESULT eventid="1273" points="471" reactiontime="+79" swimtime="00:00:57.72" resultid="18389" heatid="19387" lane="1" entrytime="00:00:56.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="494" reactiontime="+78" swimtime="00:00:27.56" resultid="18390" heatid="19462" lane="5" entrytime="00:00:27.20" />
                <RESULT eventid="1474" points="391" reactiontime="+69" swimtime="00:01:06.89" resultid="18391" heatid="19478" lane="0" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="18392" heatid="19496" lane="9" entrytime="00:02:05.00" />
                <RESULT eventid="1613" points="449" reactiontime="+68" swimtime="00:01:02.78" resultid="18393" heatid="19524" lane="7" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="467" reactiontime="+72" swimtime="00:00:32.53" resultid="18394" heatid="19556" lane="6" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-02-18" firstname="Marek" gender="M" lastname="Stuczyński" nation="POL" athleteid="18368">
              <RESULTS>
                <RESULT eventid="1079" points="530" reactiontime="+81" swimtime="00:00:25.03" resultid="18369" heatid="19303" lane="1" entrytime="00:00:25.00" entrycourse="SCM" />
                <RESULT eventid="1273" points="522" reactiontime="+81" swimtime="00:00:55.80" resultid="18370" heatid="19387" lane="5" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="514" reactiontime="+76" swimtime="00:01:09.38" resultid="18371" heatid="19443" lane="7" entrytime="00:01:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="548" reactiontime="+82" swimtime="00:00:30.85" resultid="18372" heatid="19558" lane="1" entrytime="00:00:32.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-20" firstname="Veronica" gender="F" lastname="Campbell-Żemier" nation="POL" athleteid="18395">
              <RESULTS>
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="18396" heatid="19372" lane="0" entrytime="00:01:04.50" />
                <RESULT eventid="1388" points="436" reactiontime="+79" swimtime="00:01:22.20" resultid="18397" heatid="19432" lane="9" entrytime="00:01:25.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="476" reactiontime="+84" swimtime="00:00:36.67" resultid="18398" heatid="19544" lane="0" entrytime="00:00:39.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-06-22" firstname="Aleksandra" gender="F" lastname="Hebel" nation="POL" athleteid="18351">
              <RESULTS>
                <RESULT eventid="1062" points="352" swimtime="00:00:32.90" resultid="18352" heatid="19281" lane="9" entrytime="00:00:32.90" entrycourse="SCM" />
                <RESULT eventid="1222" points="217" reactiontime="+101" swimtime="00:03:43.82" resultid="18353" heatid="19355" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.74" />
                    <SPLIT distance="100" swimtime="00:01:44.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="312" reactiontime="+111" swimtime="00:01:15.00" resultid="18354" heatid="19371" lane="0" entrytime="00:01:14.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="230" reactiontime="+116" swimtime="00:01:41.77" resultid="18355" heatid="19427" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="297" reactiontime="+110" swimtime="00:02:45.88" resultid="18356" heatid="19483" lane="0" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                    <SPLIT distance="100" swimtime="00:01:18.58" />
                    <SPLIT distance="150" swimtime="00:02:02.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="226" reactiontime="+91" swimtime="00:03:15.64" resultid="18357" heatid="19527" lane="4" entrytime="00:03:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.67" />
                    <SPLIT distance="100" swimtime="00:01:35.88" />
                    <SPLIT distance="150" swimtime="00:02:26.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="244" reactiontime="+106" swimtime="00:00:45.79" resultid="18358" heatid="19541" lane="1" entrytime="00:00:46.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-04-16" firstname="Filip" gender="M" lastname="Żemier" nation="POL" athleteid="18380">
              <RESULTS>
                <RESULT eventid="1079" points="455" reactiontime="+71" swimtime="00:00:26.34" resultid="18381" heatid="19300" lane="3" entrytime="00:00:26.00" />
                <RESULT eventid="1273" points="413" reactiontime="+72" swimtime="00:01:00.34" resultid="18382" heatid="19385" lane="3" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="382" reactiontime="+71" swimtime="00:00:30.02" resultid="18383" heatid="19460" lane="1" entrytime="00:00:29.50" />
                <RESULT eventid="1681" points="331" swimtime="00:00:36.50" resultid="18384" heatid="19556" lane="0" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-11-09" firstname="Karol" gender="M" lastname="Żemier" nation="POL" athleteid="18373">
              <RESULTS>
                <RESULT eventid="1205" points="487" swimtime="00:00:28.24" resultid="18374" heatid="19352" lane="2" entrytime="00:00:29.00" />
                <RESULT eventid="14243" points="542" reactiontime="+74" swimtime="00:01:01.69" resultid="18375" heatid="19409" lane="6" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="521" reactiontime="+76" swimtime="00:00:27.08" resultid="18376" heatid="19461" lane="7" entrytime="00:00:28.50" />
                <RESULT eventid="1474" points="509" reactiontime="+69" swimtime="00:01:01.23" resultid="18377" heatid="19478" lane="2" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="499" reactiontime="+74" swimtime="00:01:00.58" resultid="18378" heatid="19524" lane="6" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="454" reactiontime="+75" swimtime="00:00:32.85" resultid="18379" heatid="19556" lane="7" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="Rekin Świebodzodzice 303" number="1">
              <RESULTS>
                <RESULT eventid="1548" points="572" reactiontime="+76" swimtime="00:01:39.49" resultid="18401" heatid="19502" lane="6" entrytime="00:01:45.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.09" />
                    <SPLIT distance="100" swimtime="00:00:49.55" />
                    <SPLIT distance="150" swimtime="00:01:14.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18368" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="18385" number="2" reactiontime="+29" />
                    <RELAYPOSITION athleteid="18380" number="3" reactiontime="+17" />
                    <RELAYPOSITION athleteid="18373" number="4" reactiontime="+6" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" points="537" reactiontime="+66" swimtime="00:01:51.31" resultid="18402" heatid="19424" lane="2" entrytime="00:01:55.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.13" />
                    <SPLIT distance="100" swimtime="00:00:58.28" />
                    <SPLIT distance="150" swimtime="00:01:25.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18373" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="18368" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="18385" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="18380" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="Rekin Świebodzodzice 303" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="455" reactiontime="+70" swimtime="00:01:55.14" resultid="18399" heatid="19322" lane="7" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.30" />
                    <SPLIT distance="100" swimtime="00:00:58.15" />
                    <SPLIT distance="150" swimtime="00:01:23.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18373" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="18351" number="2" reactiontime="+77" />
                    <RELAYPOSITION athleteid="18368" number="3" reactiontime="+23" />
                    <RELAYPOSITION athleteid="18395" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="469" reactiontime="+64" swimtime="00:02:05.06" resultid="18400" heatid="19564" lane="3" entrytime="00:02:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.00" />
                    <SPLIT distance="100" swimtime="00:01:04.31" />
                    <SPLIT distance="150" swimtime="00:01:32.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18373" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="18395" number="2" reactiontime="+27" />
                    <RELAYPOSITION athleteid="18368" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="18351" number="4" reactiontime="+70" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="03315" nation="POL" region="PO" clubid="16703" name="KU AZS UAM Poznań">
          <CONTACT city="Poznań" email="kukowalazs@gmail.com" name="Kowalik" phone="603965223" state="WLKP" street="Zagajnikowa 9" zip="61-602" />
          <ATHLETES>
            <ATHLETE birthdate="1994-03-19" firstname="Damian" gender="M" lastname="Kowalik" nation="POL" license="103315200009" athleteid="16704">
              <RESULTS>
                <RESULT eventid="1079" points="526" reactiontime="+70" swimtime="00:00:25.09" resultid="16705" heatid="19303" lane="3" entrytime="00:00:24.50" />
                <RESULT eventid="1205" points="425" reactiontime="+55" swimtime="00:00:29.54" resultid="16706" heatid="19353" lane="9" entrytime="00:00:28.43" />
                <RESULT eventid="14243" points="525" reactiontime="+66" swimtime="00:01:02.35" resultid="16707" heatid="19410" lane="8" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="563" reactiontime="+73" swimtime="00:00:26.39" resultid="16708" heatid="19464" lane="2" entrytime="00:00:25.80" />
                <RESULT eventid="1613" points="508" reactiontime="+73" swimtime="00:01:00.22" resultid="16709" heatid="19525" lane="2" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-07-20" firstname="Krzysztof" gender="M" lastname="Strzelczyk" nation="POL" athleteid="16761">
              <RESULTS>
                <RESULT eventid="1079" points="195" reactiontime="+85" swimtime="00:00:34.88" resultid="16762" heatid="19290" lane="0" entrytime="00:00:33.00" />
                <RESULT eventid="1273" points="161" reactiontime="+82" swimtime="00:01:22.58" resultid="16763" heatid="19377" lane="8" entrytime="00:01:23.00" />
                <RESULT eventid="14243" points="131" reactiontime="+102" swimtime="00:01:38.87" resultid="16764" heatid="19399" lane="2" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="124" reactiontime="+89" swimtime="00:00:43.62" resultid="16765" heatid="19452" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="1508" points="144" reactiontime="+101" swimtime="00:03:09.47" resultid="16766" heatid="19488" lane="7" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.26" />
                    <SPLIT distance="100" swimtime="00:01:30.29" />
                    <SPLIT distance="150" swimtime="00:02:20.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="143" reactiontime="+90" swimtime="00:06:45.15" resultid="16767" heatid="19701" lane="0" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.30" />
                    <SPLIT distance="100" swimtime="00:01:34.28" />
                    <SPLIT distance="150" swimtime="00:03:18.24" />
                    <SPLIT distance="200" swimtime="00:04:09.68" />
                    <SPLIT distance="250" swimtime="00:05:02.09" />
                    <SPLIT distance="300" swimtime="00:05:54.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Jakub" gender="M" lastname="Sterczyński" nation="POL" license="103315200002" athleteid="16739">
              <RESULTS>
                <RESULT eventid="1079" points="464" reactiontime="+73" swimtime="00:00:26.16" resultid="16740" heatid="19301" lane="3" entrytime="00:00:26.00" />
                <RESULT eventid="1113" points="468" reactiontime="+74" swimtime="00:02:21.12" resultid="16741" heatid="19317" lane="4" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.16" />
                    <SPLIT distance="100" swimtime="00:01:06.26" />
                    <SPLIT distance="150" swimtime="00:01:46.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="384" reactiontime="+67" swimtime="00:00:30.55" resultid="16742" heatid="19352" lane="9" entrytime="00:00:30.00" />
                <RESULT eventid="14243" points="541" reactiontime="+75" swimtime="00:01:01.71" resultid="16743" heatid="19409" lane="1" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="462" reactiontime="+77" swimtime="00:00:28.19" resultid="16744" heatid="19461" lane="2" entrytime="00:00:28.50" />
                <RESULT eventid="1474" points="447" reactiontime="+81" swimtime="00:01:03.95" resultid="16745" heatid="19478" lane="1" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="446" reactiontime="+77" swimtime="00:01:02.89" resultid="16746" heatid="19524" lane="5" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-03-14" firstname="Jarosław" gender="M" lastname="Bystry" nation="POL" athleteid="16768">
              <RESULTS>
                <RESULT eventid="1079" points="378" reactiontime="+78" swimtime="00:00:28.00" resultid="16769" heatid="19297" lane="8" entrytime="00:00:28.00" />
                <RESULT eventid="1273" points="385" reactiontime="+77" swimtime="00:01:01.73" resultid="16770" heatid="19383" lane="8" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="340" reactiontime="+80" swimtime="00:00:31.23" resultid="16771" heatid="19455" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1508" points="333" reactiontime="+85" swimtime="00:02:23.30" resultid="16772" heatid="19491" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                    <SPLIT distance="100" swimtime="00:01:09.23" />
                    <SPLIT distance="150" swimtime="00:01:46.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-05" firstname="Piotr" gender="M" lastname="Kowalik" nation="POL" license="103315200006" athleteid="16710">
              <RESULTS>
                <RESULT eventid="1079" points="549" reactiontime="+65" swimtime="00:00:24.73" resultid="16711" heatid="19304" lane="9" entrytime="00:00:24.30" />
                <RESULT eventid="1205" points="535" swimtime="00:00:27.36" resultid="16712" heatid="19353" lane="7" entrytime="00:00:27.20" />
                <RESULT eventid="14243" points="549" reactiontime="+66" swimtime="00:01:01.41" resultid="16713" heatid="19410" lane="6" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="627" reactiontime="+68" swimtime="00:00:25.46" resultid="16714" heatid="19464" lane="3" entrytime="00:00:25.20" />
                <RESULT eventid="1613" points="593" reactiontime="+69" swimtime="00:00:57.21" resultid="16715" heatid="19525" lane="5" entrytime="00:00:57.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-02-17" firstname="Jerzy" gender="M" lastname="Gniazdowski" nation="POL" license="103315700026" athleteid="16716">
              <RESULTS>
                <RESULT eventid="1079" points="406" reactiontime="+63" swimtime="00:00:27.36" resultid="16717" heatid="19302" lane="3" entrytime="00:00:25.17" />
                <RESULT eventid="1205" points="274" reactiontime="+71" swimtime="00:00:34.20" resultid="16718" heatid="19350" lane="9" entrytime="00:00:33.00" />
                <RESULT eventid="1273" points="425" reactiontime="+63" swimtime="00:00:59.74" resultid="16719" heatid="19387" lane="4" entrytime="00:00:55.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="388" reactiontime="+72" swimtime="00:00:29.88" resultid="16720" heatid="19461" lane="1" entrytime="00:00:28.94" />
                <RESULT eventid="1508" points="376" reactiontime="+65" swimtime="00:02:17.64" resultid="16721" heatid="19495" lane="4" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                    <SPLIT distance="100" swimtime="00:01:05.30" />
                    <SPLIT distance="150" swimtime="00:01:40.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="16722" heatid="19523" lane="8" entrytime="00:01:08.08" />
                <RESULT eventid="1681" points="342" reactiontime="+66" swimtime="00:00:36.09" resultid="16723" heatid="19553" lane="4" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-11-18" firstname="Marek" gender="M" lastname="Michałkowski" nation="POL" athleteid="16724">
              <RESULTS>
                <RESULT eventid="1079" points="570" reactiontime="+72" swimtime="00:00:24.43" resultid="16725" heatid="19303" lane="5" entrytime="00:00:24.50" />
                <RESULT eventid="14243" points="538" reactiontime="+77" swimtime="00:01:01.82" resultid="16726" heatid="19410" lane="2" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="569" reactiontime="+72" swimtime="00:01:07.09" resultid="16727" heatid="19443" lane="2" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="576" reactiontime="+75" swimtime="00:00:30.33" resultid="16728" heatid="19560" lane="1" entrytime="00:00:30.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-04-18" firstname="Karolina" gender="F" lastname="Sterczyńska" nation="POL" license="103315100003" athleteid="16747">
              <RESULTS>
                <RESULT eventid="1062" points="598" reactiontime="+83" swimtime="00:00:27.58" resultid="16748" heatid="19283" lane="5" entrytime="00:00:27.50" />
                <RESULT eventid="1256" points="597" reactiontime="+80" swimtime="00:01:00.46" resultid="16749" heatid="19372" lane="6" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="529" reactiontime="+92" swimtime="00:01:10.03" resultid="16750" heatid="19396" lane="1" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="499" reactiontime="+85" swimtime="00:01:18.62" resultid="16751" heatid="19432" lane="2" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="500" reactiontime="+81" swimtime="00:00:30.70" resultid="16752" heatid="19449" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1664" points="507" reactiontime="+80" swimtime="00:00:35.91" resultid="16753" heatid="19545" lane="5" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-12-27" firstname="Bartosz" gender="M" lastname="Jankowiak" nation="POL" athleteid="16729">
              <RESULTS>
                <RESULT eventid="1079" points="300" reactiontime="+80" swimtime="00:00:30.24" resultid="16730" heatid="19296" lane="0" entrytime="00:00:29.00" />
                <RESULT eventid="1273" points="296" reactiontime="+82" swimtime="00:01:07.43" resultid="16731" heatid="19381" lane="8" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="249" reactiontime="+89" swimtime="00:01:19.85" resultid="16732" heatid="19401" lane="1" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="258" reactiontime="+83" swimtime="00:02:35.90" resultid="16733" heatid="19490" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="100" swimtime="00:01:14.98" />
                    <SPLIT distance="150" swimtime="00:01:56.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="274" swimtime="00:05:26.63" resultid="16734" heatid="19704" lane="6" entrytime="00:05:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                    <SPLIT distance="100" swimtime="00:01:14.90" />
                    <SPLIT distance="150" swimtime="00:01:56.57" />
                    <SPLIT distance="200" swimtime="00:02:38.85" />
                    <SPLIT distance="250" swimtime="00:03:21.52" />
                    <SPLIT distance="300" swimtime="00:04:04.01" />
                    <SPLIT distance="350" swimtime="00:04:46.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14189" reactiontime="+93" status="OTL" swimtime="00:11:27.50" resultid="18969" heatid="19616" lane="2" entrytime="00:11:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                    <SPLIT distance="100" swimtime="00:01:17.12" />
                    <SPLIT distance="150" swimtime="00:02:00.15" />
                    <SPLIT distance="200" swimtime="00:04:10.50" />
                    <SPLIT distance="350" swimtime="00:04:54.14" />
                    <SPLIT distance="400" swimtime="00:05:38.03" />
                    <SPLIT distance="450" swimtime="00:06:21.99" />
                    <SPLIT distance="550" swimtime="00:08:33.62" />
                    <SPLIT distance="600" swimtime="00:09:17.99" />
                    <SPLIT distance="650" swimtime="00:10:01.83" />
                    <SPLIT distance="700" swimtime="00:10:45.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-07-15" firstname="Marcin" gender="M" lastname="Tomczak" nation="POL" athleteid="16735">
              <RESULTS>
                <RESULT eventid="1273" points="302" reactiontime="+75" swimtime="00:01:06.92" resultid="16736" heatid="19382" lane="5" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="318" reactiontime="+82" swimtime="00:02:25.45" resultid="16737" heatid="19492" lane="2" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.96" />
                    <SPLIT distance="100" swimtime="00:01:10.68" />
                    <SPLIT distance="150" swimtime="00:01:48.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="306" swimtime="00:05:14.64" resultid="16738" heatid="19706" lane="0" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                    <SPLIT distance="100" swimtime="00:01:12.29" />
                    <SPLIT distance="150" swimtime="00:01:50.84" />
                    <SPLIT distance="200" swimtime="00:02:30.59" />
                    <SPLIT distance="250" swimtime="00:03:11.37" />
                    <SPLIT distance="300" swimtime="00:03:52.94" />
                    <SPLIT distance="350" swimtime="00:04:34.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-27" firstname="Maciej" gender="M" lastname="Waliński" nation="POL" athleteid="16754">
              <RESULTS>
                <RESULT eventid="1079" points="320" reactiontime="+79" swimtime="00:00:29.61" resultid="16755" heatid="19293" lane="1" entrytime="00:00:30.00" />
                <RESULT eventid="1273" points="303" reactiontime="+71" swimtime="00:01:06.88" resultid="16756" heatid="19379" lane="9" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="216" reactiontime="+73" swimtime="00:01:23.78" resultid="16757" heatid="19400" lane="7" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="215" reactiontime="+77" swimtime="00:00:36.38" resultid="16758" heatid="19454" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1508" points="258" reactiontime="+81" swimtime="00:02:36.07" resultid="16759" heatid="19489" lane="8" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                    <SPLIT distance="100" swimtime="00:01:14.92" />
                    <SPLIT distance="150" swimtime="00:01:55.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="233" reactiontime="+78" swimtime="00:05:44.68" resultid="16760" heatid="19701" lane="5" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.39" />
                    <SPLIT distance="100" swimtime="00:01:16.42" />
                    <SPLIT distance="150" swimtime="00:01:58.39" />
                    <SPLIT distance="200" swimtime="00:02:42.22" />
                    <SPLIT distance="250" swimtime="00:03:27.61" />
                    <SPLIT distance="300" swimtime="00:04:14.06" />
                    <SPLIT distance="350" swimtime="00:05:00.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" points="511" reactiontime="+75" swimtime="00:01:43.26" resultid="16773" heatid="19502" lane="2" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.47" />
                    <SPLIT distance="100" swimtime="00:00:53.44" />
                    <SPLIT distance="150" swimtime="00:01:18.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16724" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="16754" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="16739" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="16710" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" points="496" reactiontime="+71" swimtime="00:01:54.31" resultid="16774" heatid="19424" lane="6" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.59" />
                    <SPLIT distance="100" swimtime="00:01:00.60" />
                    <SPLIT distance="150" swimtime="00:01:25.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16739" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="16724" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="16710" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="16754" number="4" reactiontime="+62" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT comment="O4 - Start wykonany przed sygnłem (przedwczesny start) (Time: 19:48)" eventid="1548" reactiontime="+66" status="DSQ" swimtime="00:02:03.05" resultid="16775" heatid="19501" lane="8" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.92" />
                    <SPLIT distance="100" swimtime="00:01:05.49" />
                    <SPLIT distance="150" swimtime="00:01:35.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16735" number="1" reactiontime="+66" status="DSQ" />
                    <RELAYPOSITION athleteid="16761" number="2" reactiontime="0" status="DSQ" />
                    <RELAYPOSITION athleteid="16729" number="3" reactiontime="+70" status="DSQ" />
                    <RELAYPOSITION athleteid="16768" number="4" reactiontime="+42" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" points="245" reactiontime="+86" swimtime="00:02:24.57" resultid="16776" heatid="19422" lane="3" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                    <SPLIT distance="100" swimtime="00:01:18.21" />
                    <SPLIT distance="150" swimtime="00:01:49.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16735" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="16729" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="16768" number="3" reactiontime="+77" />
                    <RELAYPOSITION athleteid="16761" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="AZS UW" nation="POL" region="MAZ" clubid="15715" name="KU AZS Uniwersytet Warszawski">
          <CONTACT city="Warszawa" email="marek.baranowski91@gmail.com" name="Baranowski Marek" phone="602445201" state="MAZ" street="Krakowskie Przedmieście 26/28" zip="00-927" />
          <ATHLETES>
            <ATHLETE birthdate="1996-08-27" firstname="Edyta" gender="F" lastname="Ilcewicz" nation="POL" license="108114600029" athleteid="15728">
              <RESULTS>
                <RESULT eventid="1096" points="426" reactiontime="+78" swimtime="00:02:41.93" resultid="15729" heatid="19309" lane="5" entrytime="00:02:29.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.41" />
                    <SPLIT distance="100" swimtime="00:01:16.21" />
                    <SPLIT distance="150" swimtime="00:02:03.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="525" reactiontime="+78" swimtime="00:01:03.09" resultid="15730" heatid="19372" lane="2" entrytime="00:01:00.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="499" reactiontime="+77" swimtime="00:01:11.42" resultid="15731" heatid="19396" lane="3" entrytime="00:01:09.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="478" reactiontime="+77" swimtime="00:01:19.71" resultid="15732" heatid="19432" lane="3" entrytime="00:01:18.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="473" reactiontime="+75" swimtime="00:00:36.74" resultid="15733" heatid="19545" lane="3" entrytime="00:00:35.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-15" firstname="Marek" gender="M" lastname="Baranowski" nation="POL" license="108114700035" athleteid="15723">
              <RESULTS>
                <RESULT eventid="1079" points="479" reactiontime="+81" swimtime="00:00:25.88" resultid="15724" heatid="19302" lane="1" entrytime="00:00:25.87" entrycourse="SCM" />
                <RESULT eventid="1273" points="521" reactiontime="+73" swimtime="00:00:55.82" resultid="15725" heatid="19386" lane="5" entrytime="00:00:57.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="506" reactiontime="+74" swimtime="00:02:04.69" resultid="15726" heatid="19495" lane="3" entrytime="00:02:05.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.62" />
                    <SPLIT distance="100" swimtime="00:01:00.57" />
                    <SPLIT distance="150" swimtime="00:01:32.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="457" reactiontime="+73" swimtime="00:04:35.43" resultid="15727" heatid="19708" lane="9" entrytime="00:04:36.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.74" />
                    <SPLIT distance="100" swimtime="00:01:02.93" />
                    <SPLIT distance="150" swimtime="00:01:36.79" />
                    <SPLIT distance="200" swimtime="00:02:11.67" />
                    <SPLIT distance="250" swimtime="00:02:47.03" />
                    <SPLIT distance="300" swimtime="00:03:22.90" />
                    <SPLIT distance="350" swimtime="00:03:59.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06614" nation="POL" region="MAZ" clubid="14986" name="Legia Warszawa">
          <CONTACT email="janek@plywanielegia.pl" name="Peńsko" phone="600826305" />
          <ATHLETES>
            <ATHLETE birthdate="1981-10-24" firstname="Marcin" gender="M" lastname="Wilczęga" nation="POL" athleteid="14989">
              <RESULTS>
                <RESULT eventid="1079" points="430" reactiontime="+76" swimtime="00:00:26.84" resultid="14990" heatid="19302" lane="7" entrytime="00:00:25.82" />
                <RESULT eventid="14243" points="398" reactiontime="+70" swimtime="00:01:08.38" resultid="14991" heatid="19408" lane="9" entrytime="00:01:07.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-05-11" firstname="Maciej" gender="M" lastname="Rybicki" nation="POL" athleteid="15004">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="15005" heatid="19293" lane="3" entrytime="00:00:29.65" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="15006" heatid="19347" lane="9" entrytime="00:00:39.89" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-08-13" firstname="Roman" gender="M" lastname="Kozłowski" nation="POL" athleteid="15007">
              <RESULTS>
                <RESULT eventid="1079" points="323" swimtime="00:00:29.51" resultid="15008" heatid="19295" lane="0" entrytime="00:00:29.00" />
                <RESULT eventid="1205" points="252" reactiontime="+83" swimtime="00:00:35.16" resultid="15009" heatid="19351" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="14243" points="320" reactiontime="+81" swimtime="00:01:13.48" resultid="15010" heatid="19402" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="324" reactiontime="+73" swimtime="00:00:31.71" resultid="15011" heatid="19458" lane="6" entrytime="00:00:31.00" />
                <RESULT eventid="1681" points="355" reactiontime="+73" swimtime="00:00:35.66" resultid="15012" heatid="19551" lane="2" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-07-12" firstname="Filip" gender="M" lastname="Rowiński" nation="POL" athleteid="14987">
              <RESULTS>
                <RESULT eventid="14207" points="444" reactiontime="+69" swimtime="00:18:31.53" resultid="14988" heatid="19623" lane="3" entrytime="00:19:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                    <SPLIT distance="100" swimtime="00:01:06.13" />
                    <SPLIT distance="150" swimtime="00:01:42.03" />
                    <SPLIT distance="200" swimtime="00:02:18.63" />
                    <SPLIT distance="250" swimtime="00:02:54.95" />
                    <SPLIT distance="300" swimtime="00:03:32.10" />
                    <SPLIT distance="350" swimtime="00:04:09.77" />
                    <SPLIT distance="400" swimtime="00:04:47.11" />
                    <SPLIT distance="450" swimtime="00:05:24.43" />
                    <SPLIT distance="500" swimtime="00:06:02.47" />
                    <SPLIT distance="550" swimtime="00:06:40.13" />
                    <SPLIT distance="600" swimtime="00:07:17.99" />
                    <SPLIT distance="650" swimtime="00:07:55.67" />
                    <SPLIT distance="700" swimtime="00:08:33.57" />
                    <SPLIT distance="750" swimtime="00:09:11.13" />
                    <SPLIT distance="800" swimtime="00:09:48.76" />
                    <SPLIT distance="850" swimtime="00:10:26.41" />
                    <SPLIT distance="900" swimtime="00:11:03.89" />
                    <SPLIT distance="950" swimtime="00:11:41.63" />
                    <SPLIT distance="1000" swimtime="00:12:19.62" />
                    <SPLIT distance="1050" swimtime="00:12:57.67" />
                    <SPLIT distance="1100" swimtime="00:13:35.80" />
                    <SPLIT distance="1150" swimtime="00:14:13.89" />
                    <SPLIT distance="1200" swimtime="00:14:52.07" />
                    <SPLIT distance="1250" swimtime="00:15:30.10" />
                    <SPLIT distance="1300" swimtime="00:16:07.83" />
                    <SPLIT distance="1350" swimtime="00:16:46.26" />
                    <SPLIT distance="1400" swimtime="00:17:23.58" />
                    <SPLIT distance="1450" swimtime="00:17:59.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-05-05" firstname="Bogdan" gender="M" lastname="Dubiński" nation="POL" athleteid="18960">
              <RESULTS>
                <RESULT eventid="1079" points="217" reactiontime="+76" swimtime="00:00:33.69" resultid="18961" heatid="19291" lane="0" entrytime="00:00:32.00" />
                <RESULT eventid="14207" points="157" reactiontime="+98" swimtime="00:26:11.98" resultid="18962" heatid="19620" lane="3" entrytime="00:26:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.45" />
                    <SPLIT distance="100" swimtime="00:01:30.16" />
                    <SPLIT distance="150" swimtime="00:02:18.99" />
                    <SPLIT distance="200" swimtime="00:03:07.66" />
                    <SPLIT distance="250" swimtime="00:03:57.90" />
                    <SPLIT distance="300" swimtime="00:04:49.31" />
                    <SPLIT distance="350" swimtime="00:05:41.82" />
                    <SPLIT distance="400" swimtime="00:06:34.77" />
                    <SPLIT distance="450" swimtime="00:07:28.21" />
                    <SPLIT distance="500" swimtime="00:08:21.92" />
                    <SPLIT distance="550" swimtime="00:09:14.65" />
                    <SPLIT distance="600" swimtime="00:10:09.05" />
                    <SPLIT distance="650" swimtime="00:11:02.55" />
                    <SPLIT distance="700" swimtime="00:11:55.86" />
                    <SPLIT distance="750" swimtime="00:12:50.15" />
                    <SPLIT distance="800" swimtime="00:13:43.47" />
                    <SPLIT distance="850" swimtime="00:14:37.63" />
                    <SPLIT distance="900" swimtime="00:15:32.37" />
                    <SPLIT distance="950" swimtime="00:16:26.58" />
                    <SPLIT distance="1000" swimtime="00:17:20.53" />
                    <SPLIT distance="1050" swimtime="00:18:14.64" />
                    <SPLIT distance="1100" swimtime="00:19:08.67" />
                    <SPLIT distance="1150" swimtime="00:20:02.87" />
                    <SPLIT distance="1200" swimtime="00:20:56.57" />
                    <SPLIT distance="1250" swimtime="00:21:50.23" />
                    <SPLIT distance="1300" swimtime="00:22:43.20" />
                    <SPLIT distance="1350" swimtime="00:23:36.98" />
                    <SPLIT distance="1400" swimtime="00:24:30.39" />
                    <SPLIT distance="1450" swimtime="00:25:22.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="146" reactiontime="+76" swimtime="00:00:42.17" resultid="18963" heatid="19346" lane="7" entrytime="00:00:41.00" />
                <RESULT eventid="1341" points="68" reactiontime="+104" swimtime="00:04:24.80" resultid="18964" heatid="19414" lane="3" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.18" />
                    <SPLIT distance="100" swimtime="00:01:51.65" />
                    <SPLIT distance="150" swimtime="00:02:59.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="143" swimtime="00:01:33.37" resultid="18965" heatid="19473" lane="8" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="131" reactiontime="+96" swimtime="00:07:42.55" resultid="18966" heatid="19508" lane="8" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:59.69" />
                    <SPLIT distance="100" swimtime="00:03:53.66" />
                    <SPLIT distance="150" swimtime="00:05:01.53" />
                    <SPLIT distance="300" swimtime="00:06:06.23" />
                    <SPLIT distance="350" swimtime="00:06:56.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="123" reactiontime="+87" swimtime="00:03:32.26" resultid="18967" heatid="19533" lane="1" entrytime="00:03:35.00" />
                <RESULT eventid="1744" points="154" swimtime="00:06:35.42" resultid="18968" heatid="19702" lane="0" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.04" />
                    <SPLIT distance="100" swimtime="00:01:30.55" />
                    <SPLIT distance="150" swimtime="00:02:20.55" />
                    <SPLIT distance="200" swimtime="00:03:11.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-06-15" firstname="Aleksandra" gender="F" lastname="Marianek" nation="POL" athleteid="14992">
              <RESULTS>
                <RESULT eventid="1222" points="317" reactiontime="+91" swimtime="00:03:17.21" resultid="14993" heatid="19357" lane="0" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.13" />
                    <SPLIT distance="100" swimtime="00:01:35.51" />
                    <SPLIT distance="150" swimtime="00:02:27.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="299" reactiontime="+80" swimtime="00:01:33.25" resultid="14994" heatid="19431" lane="9" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="311" reactiontime="+82" swimtime="00:00:42.26" resultid="14995" heatid="19543" lane="2" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-05-07" firstname="Agnieszka" gender="F" lastname="Kaczmarek" nation="POL" athleteid="14996">
              <RESULTS>
                <RESULT eventid="1062" points="509" reactiontime="+79" swimtime="00:00:29.09" resultid="14997" heatid="19283" lane="8" entrytime="00:00:28.50" />
                <RESULT eventid="1096" points="478" reactiontime="+84" swimtime="00:02:35.79" resultid="14998" heatid="19309" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                    <SPLIT distance="100" swimtime="00:01:13.84" />
                    <SPLIT distance="150" swimtime="00:01:58.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="490" reactiontime="+68" swimtime="00:00:32.54" resultid="14999" heatid="19341" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="14225" points="473" reactiontime="+82" swimtime="00:01:12.69" resultid="15000" heatid="19396" lane="7" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="448" reactiontime="+73" swimtime="00:01:11.87" resultid="15001" heatid="19469" lane="3" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="405" reactiontime="+76" swimtime="00:02:41.09" resultid="15002" heatid="19529" lane="4" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.63" />
                    <SPLIT distance="100" swimtime="00:01:17.06" />
                    <SPLIT distance="150" swimtime="00:01:58.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="428" reactiontime="+89" swimtime="00:00:38.00" resultid="15003" heatid="19544" lane="2" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="15850" name="Masters Białystok">
          <CONTACT internet="mbzgloszenia@gmail.com" name="MASTERS BIAŁYSTOK" />
          <ATHLETES>
            <ATHLETE birthdate="1965-01-01" firstname="Andrzej" gender="M" lastname="Twarowski" nation="POL" athleteid="15856">
              <RESULTS>
                <RESULT eventid="1113" points="189" reactiontime="+105" swimtime="00:03:10.85" resultid="15857" heatid="19312" lane="0" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.91" />
                    <SPLIT distance="100" swimtime="00:01:24.27" />
                    <SPLIT distance="150" swimtime="00:02:20.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="205" reactiontime="+103" swimtime="00:03:24.06" resultid="15858" heatid="19361" lane="3" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.14" />
                    <SPLIT distance="100" swimtime="00:01:37.64" />
                    <SPLIT distance="150" swimtime="00:02:32.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="124" reactiontime="+106" swimtime="00:03:37.28" resultid="15859" heatid="19415" lane="1" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.67" />
                    <SPLIT distance="100" swimtime="00:01:44.08" />
                    <SPLIT distance="150" swimtime="00:02:42.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="212" reactiontime="+101" swimtime="00:01:33.23" resultid="15860" heatid="19437" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="178" reactiontime="+102" swimtime="00:06:58.56" resultid="15861" heatid="19508" lane="5" entrytime="00:06:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.46" />
                    <SPLIT distance="100" swimtime="00:01:42.64" />
                    <SPLIT distance="150" swimtime="00:02:35.62" />
                    <SPLIT distance="200" swimtime="00:03:28.92" />
                    <SPLIT distance="250" swimtime="00:04:26.73" />
                    <SPLIT distance="300" swimtime="00:05:24.19" />
                    <SPLIT distance="350" swimtime="00:06:14.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="191" reactiontime="+77" swimtime="00:03:03.33" resultid="15862" heatid="19534" lane="5" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.59" />
                    <SPLIT distance="100" swimtime="00:01:28.02" />
                    <SPLIT distance="150" swimtime="00:02:15.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="213" reactiontime="+103" swimtime="00:00:42.26" resultid="15863" heatid="19552" lane="3" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-01" firstname="Dominika" gender="F" lastname="Michalik" nation="POL" athleteid="15851">
              <RESULTS>
                <RESULT eventid="1147" points="443" reactiontime="+82" swimtime="00:10:28.58" resultid="15852" heatid="19596" lane="3" entrytime="00:10:17.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                    <SPLIT distance="100" swimtime="00:01:13.49" />
                    <SPLIT distance="150" swimtime="00:01:52.48" />
                    <SPLIT distance="200" swimtime="00:02:32.03" />
                    <SPLIT distance="250" swimtime="00:03:11.73" />
                    <SPLIT distance="300" swimtime="00:03:50.99" />
                    <SPLIT distance="350" swimtime="00:04:30.28" />
                    <SPLIT distance="400" swimtime="00:05:09.23" />
                    <SPLIT distance="450" swimtime="00:05:49.18" />
                    <SPLIT distance="500" swimtime="00:06:29.00" />
                    <SPLIT distance="550" swimtime="00:07:09.38" />
                    <SPLIT distance="600" swimtime="00:07:49.38" />
                    <SPLIT distance="650" swimtime="00:08:30.05" />
                    <SPLIT distance="700" swimtime="00:09:09.76" />
                    <SPLIT distance="750" swimtime="00:09:49.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="458" swimtime="00:01:06.04" resultid="15853" heatid="19372" lane="9" entrytime="00:01:05.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="488" reactiontime="+82" swimtime="00:02:20.70" resultid="15854" heatid="19484" lane="6" entrytime="00:02:19.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                    <SPLIT distance="100" swimtime="00:01:08.25" />
                    <SPLIT distance="150" swimtime="00:01:44.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="482" reactiontime="+82" swimtime="00:04:59.10" resultid="15855" heatid="19698" lane="3" entrytime="00:04:56.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                    <SPLIT distance="100" swimtime="00:01:09.70" />
                    <SPLIT distance="150" swimtime="00:01:47.16" />
                    <SPLIT distance="200" swimtime="00:02:25.29" />
                    <SPLIT distance="250" swimtime="00:03:04.03" />
                    <SPLIT distance="300" swimtime="00:03:43.03" />
                    <SPLIT distance="350" swimtime="00:04:21.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="RZ" clubid="16686" name="Masters Ikar Mielec">
          <CONTACT city="CHORZELÓW" email="sebastianboicetta@gmail.com" name="SEBASTIAN BOICETTA" phone="501072284" street="MALINIE 629" zip="39-331" />
          <ATHLETES>
            <ATHLETE birthdate="1988-06-09" firstname="Daniel" gender="M" lastname="Paduch" nation="POL" license="503208700002" athleteid="16692">
              <RESULTS>
                <RESULT eventid="14207" points="494" reactiontime="+85" swimtime="00:17:52.55" resultid="16693" heatid="19623" lane="4" entrytime="00:18:10.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.89" />
                    <SPLIT distance="100" swimtime="00:01:05.39" />
                    <SPLIT distance="150" swimtime="00:01:40.48" />
                    <SPLIT distance="200" swimtime="00:02:15.12" />
                    <SPLIT distance="250" swimtime="00:02:50.09" />
                    <SPLIT distance="300" swimtime="00:03:25.44" />
                    <SPLIT distance="350" swimtime="00:04:01.10" />
                    <SPLIT distance="400" swimtime="00:04:37.08" />
                    <SPLIT distance="450" swimtime="00:05:12.83" />
                    <SPLIT distance="500" swimtime="00:05:48.92" />
                    <SPLIT distance="550" swimtime="00:06:25.50" />
                    <SPLIT distance="600" swimtime="00:07:01.75" />
                    <SPLIT distance="650" swimtime="00:07:37.68" />
                    <SPLIT distance="700" swimtime="00:08:13.85" />
                    <SPLIT distance="750" swimtime="00:08:50.19" />
                    <SPLIT distance="800" swimtime="00:09:26.68" />
                    <SPLIT distance="850" swimtime="00:10:03.15" />
                    <SPLIT distance="900" swimtime="00:10:39.31" />
                    <SPLIT distance="950" swimtime="00:11:15.55" />
                    <SPLIT distance="1000" swimtime="00:11:52.34" />
                    <SPLIT distance="1050" swimtime="00:12:28.09" />
                    <SPLIT distance="1100" swimtime="00:13:04.11" />
                    <SPLIT distance="1150" swimtime="00:13:40.52" />
                    <SPLIT distance="1200" swimtime="00:14:16.63" />
                    <SPLIT distance="1250" swimtime="00:14:52.76" />
                    <SPLIT distance="1300" swimtime="00:15:29.57" />
                    <SPLIT distance="1350" swimtime="00:16:05.15" />
                    <SPLIT distance="1400" swimtime="00:16:41.77" />
                    <SPLIT distance="1450" swimtime="00:17:17.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="528" reactiontime="+79" swimtime="00:02:14.24" resultid="16694" heatid="19418" lane="6" entrytime="00:02:16.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.01" />
                    <SPLIT distance="100" swimtime="00:01:04.61" />
                    <SPLIT distance="150" swimtime="00:01:39.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="467" reactiontime="+76" swimtime="00:02:08.07" resultid="16695" heatid="19495" lane="8" entrytime="00:02:08.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.71" />
                    <SPLIT distance="100" swimtime="00:01:02.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="431" reactiontime="+83" swimtime="00:05:11.53" resultid="16696" heatid="19511" lane="6" entrytime="00:05:30.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                    <SPLIT distance="100" swimtime="00:01:07.21" />
                    <SPLIT distance="150" swimtime="00:01:52.08" />
                    <SPLIT distance="200" swimtime="00:02:35.18" />
                    <SPLIT distance="250" swimtime="00:03:19.11" />
                    <SPLIT distance="300" swimtime="00:04:03.44" />
                    <SPLIT distance="350" swimtime="00:04:38.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="16697" heatid="19524" lane="9" entrytime="00:01:04.75" />
                <RESULT eventid="1744" points="465" reactiontime="+83" swimtime="00:04:33.92" resultid="16698" heatid="19708" lane="0" entrytime="00:04:35.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                    <SPLIT distance="100" swimtime="00:01:05.16" />
                    <SPLIT distance="150" swimtime="00:01:40.35" />
                    <SPLIT distance="200" swimtime="00:02:15.23" />
                    <SPLIT distance="250" swimtime="00:02:49.87" />
                    <SPLIT distance="300" swimtime="00:03:25.45" />
                    <SPLIT distance="350" swimtime="00:04:00.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-04-01" firstname="Sebastian" gender="M" lastname="Boicetta" nation="POL" athleteid="16687">
              <RESULTS>
                <RESULT eventid="1079" points="285" reactiontime="+83" swimtime="00:00:30.76" resultid="16688" heatid="19291" lane="2" entrytime="00:00:31.48" entrycourse="SCM" />
                <RESULT eventid="1205" points="211" reactiontime="+73" swimtime="00:00:37.31" resultid="16689" heatid="19347" lane="4" entrytime="00:00:36.86" />
                <RESULT eventid="14243" points="236" reactiontime="+86" swimtime="00:01:21.29" resultid="16690" heatid="19401" lane="4" entrytime="00:01:20.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="199" reactiontime="+74" swimtime="00:01:23.70" resultid="16691" heatid="19474" lane="3" entrytime="00:01:21.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="MAL" clubid="14956" name="Masters Oświęcim">
          <CONTACT city="Oświęcim" email="js.formasy@interia.pl" name="Masters Oświęcim" phone="793691105" state="MAL" zip="32-600" />
          <ATHLETES>
            <ATHLETE birthdate="1973-01-27" firstname="Robert" gender="M" lastname="Krulikowski" nation="POL" athleteid="14971">
              <RESULTS>
                <RESULT eventid="14243" points="332" reactiontime="+85" swimtime="00:01:12.59" resultid="14972" heatid="19406" lane="7" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="277" reactiontime="+80" swimtime="00:01:15.01" resultid="14973" heatid="19476" lane="3" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="14974" heatid="19523" lane="1" entrytime="00:01:08.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-11-05" firstname="Sławomir" gender="M" lastname="Formas" nation="POL" athleteid="14964">
              <RESULTS>
                <RESULT eventid="1113" points="446" reactiontime="+85" swimtime="00:02:23.43" resultid="14965" heatid="19317" lane="6" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                    <SPLIT distance="100" swimtime="00:01:08.41" />
                    <SPLIT distance="150" swimtime="00:01:48.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="503" reactiontime="+91" swimtime="00:02:31.40" resultid="14966" heatid="19365" lane="1" entrytime="00:02:36.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                    <SPLIT distance="100" swimtime="00:01:12.77" />
                    <SPLIT distance="150" swimtime="00:01:52.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="489" reactiontime="+85" swimtime="00:01:03.83" resultid="14967" heatid="19407" lane="3" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="526" reactiontime="+78" swimtime="00:01:08.86" resultid="14968" heatid="19442" lane="8" entrytime="00:01:10.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="431" reactiontime="+76" swimtime="00:00:28.84" resultid="14969" heatid="19460" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="1681" points="538" reactiontime="+76" swimtime="00:00:31.04" resultid="14970" heatid="19559" lane="2" entrytime="00:00:31.62" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="17006" name="Masters Team Biała Podlaska">
          <CONTACT email="wilhelmg@poczta.onet.pl" name="Gromisz" />
          <ATHLETES>
            <ATHLETE birthdate="1980-03-03" firstname="Tomasz" gender="M" lastname="Melańczuk" nation="POL" athleteid="17018">
              <RESULTS>
                <RESULT eventid="1113" points="431" reactiontime="+91" swimtime="00:02:25.11" resultid="17019" heatid="19316" lane="8" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.16" />
                    <SPLIT distance="100" swimtime="00:01:06.45" />
                    <SPLIT distance="150" swimtime="00:01:49.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="431" reactiontime="+74" swimtime="00:00:29.41" resultid="17020" heatid="19351" lane="6" entrytime="00:00:30.87" />
                <RESULT eventid="14243" points="477" reactiontime="+97" swimtime="00:01:04.35" resultid="17021" heatid="19407" lane="0" entrytime="00:01:08.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="490" reactiontime="+93" swimtime="00:00:27.65" resultid="17022" heatid="19459" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1474" points="435" reactiontime="+76" swimtime="00:01:04.53" resultid="17023" heatid="19477" lane="1" entrytime="00:01:08.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="413" reactiontime="+78" swimtime="00:02:21.84" resultid="17024" heatid="19536" lane="4" entrytime="00:02:33.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                    <SPLIT distance="100" swimtime="00:01:09.36" />
                    <SPLIT distance="150" swimtime="00:01:45.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-11-25" firstname="Iga" gender="F" lastname="Olszanowska" nation="POL" athleteid="17013">
              <RESULTS>
                <RESULT eventid="1187" points="485" reactiontime="+78" swimtime="00:00:32.65" resultid="17014" heatid="19341" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="14225" points="442" reactiontime="+88" swimtime="00:01:14.39" resultid="17015" heatid="19395" lane="7" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="441" reactiontime="+84" swimtime="00:00:32.02" resultid="17016" heatid="19449" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="1457" points="401" reactiontime="+72" swimtime="00:01:14.58" resultid="17017" heatid="19469" lane="7" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-03" firstname="Wilhelm" gender="M" lastname="Gromisz" nation="POL" athleteid="17007">
              <RESULTS>
                <RESULT eventid="1205" points="463" reactiontime="+80" swimtime="00:00:28.71" resultid="17008" heatid="19353" lane="0" entrytime="00:00:28.00" />
                <RESULT eventid="1273" points="453" reactiontime="+91" swimtime="00:00:58.50" resultid="17009" heatid="19387" lane="9" entrytime="00:00:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="496" reactiontime="+94" swimtime="00:00:27.53" resultid="17010" heatid="19463" lane="6" entrytime="00:00:26.80" />
                <RESULT eventid="1474" points="489" reactiontime="+77" swimtime="00:01:02.09" resultid="17011" heatid="19478" lane="3" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="423" reactiontime="+78" swimtime="00:02:20.61" resultid="17012" heatid="19537" lane="5" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                    <SPLIT distance="100" swimtime="00:01:06.14" />
                    <SPLIT distance="150" swimtime="00:01:43.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WIKRA" nation="POL" region="MAL" clubid="14781" name="Masters Wisła Kraków">
          <CONTACT email="wislaplywanie@gmail.com" internet="http://www.wislaplywanie.pl/sekcja-masters/" name="Tomasz Doniec" phone="693703490" />
          <ATHLETES>
            <ATHLETE birthdate="1969-06-25" firstname="Jerzy" gender="M" lastname="Korba" nation="POL" athleteid="14859">
              <RESULTS>
                <RESULT eventid="1079" points="427" reactiontime="+84" swimtime="00:00:26.89" resultid="14860" heatid="19298" lane="4" entrytime="00:00:27.50" entrycourse="SCM" />
                <RESULT eventid="14189" points="372" reactiontime="+101" swimtime="00:10:16.54" resultid="14861" heatid="19616" lane="4" entrytime="00:10:36.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.99" />
                    <SPLIT distance="100" swimtime="00:01:11.46" />
                    <SPLIT distance="150" swimtime="00:01:49.57" />
                    <SPLIT distance="200" swimtime="00:02:28.48" />
                    <SPLIT distance="250" swimtime="00:03:07.13" />
                    <SPLIT distance="300" swimtime="00:03:46.89" />
                    <SPLIT distance="350" swimtime="00:04:25.82" />
                    <SPLIT distance="400" swimtime="00:05:05.67" />
                    <SPLIT distance="450" swimtime="00:05:45.34" />
                    <SPLIT distance="500" swimtime="00:06:24.74" />
                    <SPLIT distance="550" swimtime="00:07:04.10" />
                    <SPLIT distance="600" swimtime="00:07:43.57" />
                    <SPLIT distance="650" swimtime="00:08:22.57" />
                    <SPLIT distance="700" swimtime="00:09:01.96" />
                    <SPLIT distance="750" swimtime="00:09:40.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="347" reactiontime="+87" swimtime="00:02:51.33" resultid="14862" heatid="19359" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                    <SPLIT distance="100" swimtime="00:01:21.10" />
                    <SPLIT distance="150" swimtime="00:02:06.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="14863" heatid="19385" lane="1" entrytime="00:00:59.90" entrycourse="SCM" />
                <RESULT eventid="1406" points="403" reactiontime="+87" swimtime="00:01:15.23" resultid="14864" heatid="19440" lane="3" entrytime="00:01:17.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="403" reactiontime="+84" swimtime="00:02:14.46" resultid="14865" heatid="19494" lane="9" entrytime="00:02:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                    <SPLIT distance="100" swimtime="00:01:05.68" />
                    <SPLIT distance="150" swimtime="00:01:40.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="425" reactiontime="+81" swimtime="00:00:33.56" resultid="14866" heatid="19556" lane="4" entrytime="00:00:34.19" entrycourse="SCM" />
                <RESULT eventid="1744" points="373" reactiontime="+89" swimtime="00:04:54.61" resultid="14867" heatid="19705" lane="8" entrytime="00:05:14.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:01:49.18" />
                    <SPLIT distance="200" swimtime="00:02:27.10" />
                    <SPLIT distance="250" swimtime="00:03:42.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1930-05-04" firstname="Stanisław" gender="M" lastname="Krokoszyński" nation="POL" athleteid="14822">
              <RESULTS>
                <RESULT eventid="1079" points="86" reactiontime="+127" swimtime="00:00:45.87" resultid="14823" heatid="19285" lane="4" entrytime="00:00:41.00" entrycourse="SCM" />
                <RESULT eventid="1113" points="54" reactiontime="+157" swimtime="00:04:48.36" resultid="14824" heatid="19310" lane="2" entrytime="00:04:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.36" />
                    <SPLIT distance="100" swimtime="00:02:33.30" />
                    <SPLIT distance="150" swimtime="00:03:50.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="52" reactiontime="+93" swimtime="00:00:59.42" resultid="14825" heatid="19343" lane="1" entrytime="00:01:00.00" entrycourse="SCM" />
                <RESULT eventid="1273" points="73" reactiontime="+122" swimtime="00:01:47.09" resultid="14826" heatid="19375" lane="2" entrytime="00:01:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="71" reactiontime="+123" swimtime="00:02:13.75" resultid="14827" heatid="19433" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="71" reactiontime="+117" swimtime="00:01:00.80" resultid="14828" heatid="19548" lane="9" entrytime="00:00:58.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-09-30" firstname="Szymon" gender="M" lastname="Łenyk" nation="POL" athleteid="14882">
              <RESULTS>
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="14883" heatid="19359" lane="7" />
                <RESULT eventid="14243" status="DNS" swimtime="00:00:00.00" resultid="14884" heatid="19398" lane="6" entrytime="00:01:50.00" entrycourse="SCM" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="14885" heatid="19435" lane="2" entrytime="00:01:50.00" entrycourse="SCM" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="14886" heatid="19488" lane="1" entrytime="00:03:05.00" entrycourse="SCM" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="14887" heatid="19549" lane="1" entrytime="00:00:48.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-02-26" firstname="Iwona" gender="F" lastname="Bednarczyk" nation="POL" athleteid="14842">
              <RESULTS>
                <RESULT eventid="1062" points="88" reactiontime="+108" swimtime="00:00:52.11" resultid="14843" heatid="19276" lane="3" entrytime="00:00:48.00" entrycourse="SCM" />
                <RESULT eventid="1147" reactiontime="+120" status="OTL" swimtime="00:19:14.58" resultid="14844" heatid="19594" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.08" />
                    <SPLIT distance="100" swimtime="00:02:06.68" />
                    <SPLIT distance="150" swimtime="00:03:18.94" />
                    <SPLIT distance="200" swimtime="00:04:33.34" />
                    <SPLIT distance="250" swimtime="00:05:48.85" />
                    <SPLIT distance="300" swimtime="00:07:03.85" />
                    <SPLIT distance="350" swimtime="00:08:19.37" />
                    <SPLIT distance="400" swimtime="00:09:32.84" />
                    <SPLIT distance="450" swimtime="00:10:45.71" />
                    <SPLIT distance="500" swimtime="00:11:58.10" />
                    <SPLIT distance="550" swimtime="00:13:10.50" />
                    <SPLIT distance="600" swimtime="00:14:22.40" />
                    <SPLIT distance="650" swimtime="00:15:35.10" />
                    <SPLIT distance="700" swimtime="00:16:48.87" />
                    <SPLIT distance="750" swimtime="00:18:02.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="62" reactiontime="+94" swimtime="00:01:04.52" resultid="14845" heatid="19336" lane="9" />
                <RESULT eventid="1256" points="70" swimtime="00:02:03.19" resultid="14846" heatid="19368" lane="9" entrytime="00:01:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="96" reactiontime="+93" swimtime="00:02:15.76" resultid="14847" heatid="19427" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="73" reactiontime="+105" swimtime="00:04:24.14" resultid="14848" heatid="19480" lane="0" entrytime="00:04:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.95" />
                    <SPLIT distance="100" swimtime="00:02:03.10" />
                    <SPLIT distance="150" swimtime="00:03:13.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="76" reactiontime="+125" swimtime="00:09:11.56" resultid="14849" heatid="19695" lane="1" entrytime="00:08:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.03" />
                    <SPLIT distance="100" swimtime="00:02:02.13" />
                    <SPLIT distance="150" swimtime="00:03:10.96" />
                    <SPLIT distance="200" swimtime="00:04:24.90" />
                    <SPLIT distance="250" swimtime="00:05:35.99" />
                    <SPLIT distance="300" swimtime="00:06:48.62" />
                    <SPLIT distance="350" swimtime="00:08:00.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-11-06" firstname="Małgorzata" gender="F" lastname="Wach" nation="POL" athleteid="14888">
              <RESULTS>
                <RESULT eventid="1062" points="248" swimtime="00:00:36.95" resultid="14889" heatid="19279" lane="9" entrytime="00:00:37.00" entrycourse="SCM" />
                <RESULT eventid="1147" reactiontime="+113" status="OTL" swimtime="00:13:55.33" resultid="14890" heatid="19594" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.91" />
                    <SPLIT distance="100" swimtime="00:01:36.16" />
                    <SPLIT distance="150" swimtime="00:02:28.26" />
                    <SPLIT distance="200" swimtime="00:03:20.39" />
                    <SPLIT distance="250" swimtime="00:04:12.46" />
                    <SPLIT distance="300" swimtime="00:05:04.83" />
                    <SPLIT distance="350" swimtime="00:05:57.44" />
                    <SPLIT distance="400" swimtime="00:09:31.42" />
                    <SPLIT distance="450" swimtime="00:10:25.11" />
                    <SPLIT distance="500" swimtime="00:11:18.32" />
                    <SPLIT distance="550" swimtime="00:12:11.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="247" reactiontime="+70" swimtime="00:00:40.86" resultid="14891" heatid="19338" lane="5" entrytime="00:00:41.00" entrycourse="SCM" />
                <RESULT eventid="1256" points="209" reactiontime="+84" swimtime="00:01:25.76" resultid="14892" heatid="19369" lane="7" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="249" reactiontime="+89" swimtime="00:02:56.04" resultid="14893" heatid="19481" lane="3" entrytime="00:03:07.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.53" />
                    <SPLIT distance="100" swimtime="00:01:26.17" />
                    <SPLIT distance="150" swimtime="00:02:12.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-03-22" firstname="Sandra" gender="F" lastname="Wolska" nation="POL" athleteid="14789">
              <RESULTS>
                <RESULT eventid="1062" points="357" reactiontime="+93" swimtime="00:00:32.75" resultid="14790" heatid="19281" lane="5" entrytime="00:00:31.95" entrycourse="SCM" />
                <RESULT eventid="1096" points="310" reactiontime="+90" swimtime="00:02:59.95" resultid="14791" heatid="19307" lane="3" entrytime="00:03:04.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.69" />
                    <SPLIT distance="100" swimtime="00:01:28.47" />
                    <SPLIT distance="150" swimtime="00:02:17.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="350" reactiontime="+90" swimtime="00:03:10.83" resultid="14792" heatid="19358" lane="0" entrytime="00:03:14.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.45" />
                    <SPLIT distance="100" swimtime="00:01:30.60" />
                    <SPLIT distance="150" swimtime="00:02:21.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="178" reactiontime="+98" swimtime="00:03:32.41" resultid="14793" heatid="19412" lane="0" entrytime="00:03:28.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.72" />
                    <SPLIT distance="100" swimtime="00:01:43.11" />
                    <SPLIT distance="150" swimtime="00:02:39.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="372" reactiontime="+94" swimtime="00:01:26.70" resultid="14794" heatid="19431" lane="4" entrytime="00:01:25.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="259" reactiontime="+83" swimtime="00:06:46.70" resultid="14795" heatid="19505" lane="9" entrytime="00:06:24.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.70" />
                    <SPLIT distance="100" swimtime="00:01:42.73" />
                    <SPLIT distance="150" swimtime="00:02:35.33" />
                    <SPLIT distance="200" swimtime="00:03:28.17" />
                    <SPLIT distance="250" swimtime="00:04:19.89" />
                    <SPLIT distance="300" swimtime="00:05:13.55" />
                    <SPLIT distance="350" swimtime="00:06:02.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="380" reactiontime="+92" swimtime="00:00:39.51" resultid="14796" heatid="19544" lane="7" entrytime="00:00:38.23" entrycourse="SCM" />
                <RESULT eventid="1721" points="295" reactiontime="+91" swimtime="00:05:52.19" resultid="14797" heatid="19696" lane="2" entrytime="00:06:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.52" />
                    <SPLIT distance="100" swimtime="00:01:21.66" />
                    <SPLIT distance="150" swimtime="00:02:06.96" />
                    <SPLIT distance="200" swimtime="00:02:52.60" />
                    <SPLIT distance="250" swimtime="00:03:38.58" />
                    <SPLIT distance="300" swimtime="00:04:24.31" />
                    <SPLIT distance="350" swimtime="00:05:10.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-12-10" firstname="Dariusz" gender="M" lastname="Wesołowski" nation="POL" athleteid="14894">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="14895" heatid="19296" lane="6" entrytime="00:00:28.60" entrycourse="SCM" />
                <RESULT eventid="14207" status="DNS" swimtime="00:00:00.00" resultid="14896" heatid="19621" lane="1" entrytime="00:24:30.00" entrycourse="SCM" />
                <RESULT eventid="1273" points="299" reactiontime="+81" swimtime="00:01:07.17" resultid="14897" heatid="19381" lane="2" entrytime="00:01:06.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K14 - Praca nóg w płaszczyźnie pionowej w dół (z wyjątkiem jednego ruchu po starcie i nawrocie) (Time: 12:02)" eventid="14243" reactiontime="+86" status="DSQ" swimtime="00:01:22.36" resultid="14898" heatid="19401" lane="0" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="279" reactiontime="+80" swimtime="00:00:33.33" resultid="14899" heatid="19455" lane="5" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1508" points="262" reactiontime="+88" swimtime="00:02:35.10" resultid="14900" heatid="19490" lane="3" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.17" />
                    <SPLIT distance="100" swimtime="00:01:15.19" />
                    <SPLIT distance="150" swimtime="00:01:55.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-09-25" firstname="Agnieszka" gender="F" lastname="Krupa" nation="POL" athleteid="14806">
              <RESULTS>
                <RESULT eventid="1096" status="DNS" swimtime="00:00:00.00" resultid="14807" heatid="19305" lane="1" />
                <RESULT eventid="1147" reactiontime="+105" status="OTL" swimtime="00:14:21.44" resultid="14808" heatid="19594" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.83" />
                    <SPLIT distance="100" swimtime="00:01:36.21" />
                    <SPLIT distance="150" swimtime="00:02:29.40" />
                    <SPLIT distance="200" swimtime="00:03:22.47" />
                    <SPLIT distance="250" swimtime="00:04:15.70" />
                    <SPLIT distance="300" swimtime="00:05:09.21" />
                    <SPLIT distance="350" swimtime="00:06:03.34" />
                    <SPLIT distance="400" swimtime="00:06:57.73" />
                    <SPLIT distance="450" swimtime="00:07:53.04" />
                    <SPLIT distance="500" swimtime="00:08:48.02" />
                    <SPLIT distance="550" swimtime="00:09:43.16" />
                    <SPLIT distance="600" swimtime="00:10:38.50" />
                    <SPLIT distance="650" swimtime="00:11:35.37" />
                    <SPLIT distance="700" swimtime="00:12:31.51" />
                    <SPLIT distance="750" swimtime="00:13:26.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="186" reactiontime="+101" swimtime="00:01:29.12" resultid="14809" heatid="19368" lane="4" entrytime="00:01:31.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="140" reactiontime="+93" swimtime="00:01:48.90" resultid="14810" heatid="19390" lane="5" entrytime="00:01:50.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" status="DNS" swimtime="00:00:00.00" resultid="14811" heatid="19465" lane="7" />
                <RESULT eventid="1491" points="160" reactiontime="+96" swimtime="00:03:23.84" resultid="14812" heatid="19481" lane="8" entrytime="00:03:26.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.25" />
                    <SPLIT distance="100" swimtime="00:01:36.59" />
                    <SPLIT distance="150" swimtime="00:02:30.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" status="DNS" swimtime="00:00:00.00" resultid="14813" heatid="19538" lane="7" />
                <RESULT eventid="1721" points="167" reactiontime="+94" swimtime="00:07:05.44" resultid="14814" heatid="19695" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.20" />
                    <SPLIT distance="100" swimtime="00:01:38.67" />
                    <SPLIT distance="150" swimtime="00:02:32.03" />
                    <SPLIT distance="200" swimtime="00:03:26.08" />
                    <SPLIT distance="250" swimtime="00:04:20.77" />
                    <SPLIT distance="300" swimtime="00:05:16.07" />
                    <SPLIT distance="350" swimtime="00:06:11.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-07-03" firstname="Jakub" gender="M" lastname="Guzik" nation="POL" athleteid="14267">
              <RESULTS>
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="14268" heatid="19365" lane="9" entrytime="00:02:40.00" />
                <RESULT eventid="14243" points="535" reactiontime="+76" swimtime="00:01:01.95" resultid="14269" heatid="19408" lane="6" entrytime="00:01:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="572" reactiontime="+78" swimtime="00:01:06.96" resultid="14270" heatid="19442" lane="3" entrytime="00:01:09.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="555" reactiontime="+77" swimtime="00:00:30.71" resultid="14271" heatid="19560" lane="0" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-03-19" firstname="Paulina" gender="F" lastname="Kujawa" nation="POL" athleteid="14829">
              <RESULTS>
                <RESULT eventid="1187" points="413" reactiontime="+53" swimtime="00:00:34.47" resultid="14830" heatid="19340" lane="8" entrytime="00:00:36.80" entrycourse="SCM" />
                <RESULT eventid="1457" points="369" reactiontime="+63" swimtime="00:01:16.69" resultid="14831" heatid="19468" lane="2" entrytime="00:01:17.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="354" reactiontime="+67" swimtime="00:02:48.39" resultid="14832" heatid="19528" lane="2" entrytime="00:03:00.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.00" />
                    <SPLIT distance="100" swimtime="00:01:23.09" />
                    <SPLIT distance="150" swimtime="00:02:06.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-09-01" firstname="Grzegorz" gender="M" lastname="Grzybczyk" nation="POL" athleteid="14815">
              <RESULTS>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="14816" heatid="19344" lane="8" entrytime="00:00:54.00" entrycourse="SCM" />
                <RESULT eventid="14243" status="DNS" swimtime="00:00:00.00" resultid="14817" heatid="19398" lane="1" entrytime="00:01:55.00" entrycourse="SCM" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="14818" heatid="19434" lane="5" entrytime="00:02:00.00" entrycourse="SCM" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="14819" heatid="19471" lane="3" entrytime="00:02:04.00" entrycourse="SCM" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="14820" heatid="19516" lane="5" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="14821" heatid="19548" lane="1" entrytime="00:00:56.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-08-23" firstname="Magdalena" gender="F" lastname="Drab" nation="POL" athleteid="14833">
              <RESULTS>
                <RESULT eventid="1062" points="597" reactiontime="+79" swimtime="00:00:27.60" resultid="14834" heatid="19283" lane="3" entrytime="00:00:27.66" entrycourse="SCM" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1096" points="639" reactiontime="+83" swimtime="00:02:21.46" resultid="14835" heatid="19309" lane="4" entrytime="00:02:26.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                    <SPLIT distance="100" swimtime="00:01:08.28" />
                    <SPLIT distance="150" swimtime="00:01:48.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="635" reactiontime="+79" swimtime="00:00:59.23" resultid="14836" heatid="19372" lane="4" entrytime="00:00:58.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="603" reactiontime="+81" swimtime="00:01:07.05" resultid="14837" heatid="19396" lane="4" entrytime="00:01:07.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1491" points="665" reactiontime="+85" swimtime="00:02:06.90" resultid="14838" heatid="19484" lane="4" entrytime="00:02:08.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                    <SPLIT distance="100" swimtime="00:01:01.32" />
                    <SPLIT distance="150" swimtime="00:01:34.53" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1555" points="647" reactiontime="+82" swimtime="00:04:59.97" resultid="14839" heatid="19505" lane="5" entrytime="00:05:04.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                    <SPLIT distance="100" swimtime="00:01:09.15" />
                    <SPLIT distance="150" swimtime="00:01:47.75" />
                    <SPLIT distance="200" swimtime="00:02:25.84" />
                    <SPLIT distance="250" swimtime="00:03:08.13" />
                    <SPLIT distance="300" swimtime="00:03:50.94" />
                    <SPLIT distance="350" swimtime="00:04:26.70" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1664" points="598" reactiontime="+82" swimtime="00:00:33.99" resultid="14840" heatid="19545" lane="4" entrytime="00:00:34.08" entrycourse="SCM" />
                <RESULT eventid="1721" points="630" reactiontime="+86" swimtime="00:04:33.55" resultid="14841" heatid="19698" lane="4" entrytime="00:04:31.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                    <SPLIT distance="100" swimtime="00:01:05.17" />
                    <SPLIT distance="150" swimtime="00:01:40.23" />
                    <SPLIT distance="200" swimtime="00:02:15.40" />
                    <SPLIT distance="250" swimtime="00:02:50.49" />
                    <SPLIT distance="300" swimtime="00:03:25.49" />
                    <SPLIT distance="350" swimtime="00:04:00.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-08-16" firstname="Tomasz" gender="M" lastname="Doniec" nation="POL" athleteid="14782">
              <RESULTS>
                <RESULT eventid="14207" status="DNS" swimtime="00:00:00.00" resultid="14783" heatid="19620" lane="0" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="14784" heatid="19361" lane="2" entrytime="00:03:24.49" entrycourse="SCM" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="14785" heatid="19437" lane="6" entrytime="00:01:28.84" entrycourse="SCM" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="14786" heatid="19488" lane="4" entrytime="00:02:58.00" entrycourse="SCM" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="14787" heatid="19552" lane="1" entrytime="00:00:38.49" entrycourse="SCM" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="14788" heatid="19701" lane="6" entrytime="00:06:31.47" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-02-07" firstname="Bogdan" gender="M" lastname="Szczurek" nation="POL" athleteid="14850">
              <RESULTS>
                <RESULT eventid="1079" points="71" reactiontime="+122" swimtime="00:00:48.90" resultid="14851" heatid="19284" lane="6" entrytime="00:00:52.00" entrycourse="SCM" />
                <RESULT eventid="14207" status="OTL" swimtime="00:00:00.00" resultid="14852" heatid="19620" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.44" />
                    <SPLIT distance="100" swimtime="00:02:08.08" />
                    <SPLIT distance="150" swimtime="00:03:17.39" />
                    <SPLIT distance="200" swimtime="00:04:30.37" />
                    <SPLIT distance="250" swimtime="00:05:43.91" />
                    <SPLIT distance="300" swimtime="00:06:55.86" />
                    <SPLIT distance="350" swimtime="00:08:08.52" />
                    <SPLIT distance="400" swimtime="00:09:25.23" />
                    <SPLIT distance="450" swimtime="00:10:45.17" />
                    <SPLIT distance="500" swimtime="00:11:53.58" />
                    <SPLIT distance="550" swimtime="00:13:07.19" />
                    <SPLIT distance="600" swimtime="00:14:22.31" />
                    <SPLIT distance="650" swimtime="00:15:40.15" />
                    <SPLIT distance="700" swimtime="00:16:53.17" />
                    <SPLIT distance="750" swimtime="00:18:08.63" />
                    <SPLIT distance="800" swimtime="00:19:23.67" />
                    <SPLIT distance="850" swimtime="00:20:41.77" />
                    <SPLIT distance="900" swimtime="00:21:54.11" />
                    <SPLIT distance="950" swimtime="00:23:11.83" />
                    <SPLIT distance="1000" swimtime="00:24:23.84" />
                    <SPLIT distance="1050" swimtime="00:25:43.36" />
                    <SPLIT distance="1100" swimtime="00:26:55.97" />
                    <SPLIT distance="1150" swimtime="00:28:17.21" />
                    <SPLIT distance="1200" swimtime="00:29:28.75" />
                    <SPLIT distance="1250" swimtime="00:30:48.17" />
                    <SPLIT distance="1300" swimtime="00:32:00.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="60" reactiontime="+42" swimtime="00:00:56.52" resultid="14853" heatid="19343" lane="7" entrytime="00:00:59.00" entrycourse="SCM" />
                <RESULT eventid="1273" points="54" reactiontime="+111" swimtime="00:01:58.60" resultid="14854" heatid="19374" lane="7" entrytime="00:02:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="14855" heatid="19471" lane="2" entrytime="00:02:09.00" entrycourse="SCM" />
                <RESULT eventid="1508" points="50" reactiontime="+127" swimtime="00:04:28.10" resultid="14856" heatid="19486" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.65" />
                    <SPLIT distance="100" swimtime="00:02:01.40" />
                    <SPLIT distance="150" swimtime="00:03:12.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="54" reactiontime="+98" swimtime="00:04:39.04" resultid="14857" heatid="19530" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.55" />
                    <SPLIT distance="100" swimtime="00:02:17.34" />
                    <SPLIT distance="150" swimtime="00:04:40.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="51" swimtime="00:09:30.22" resultid="14858" heatid="19699" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.64" />
                    <SPLIT distance="150" swimtime="00:04:37.22" />
                    <SPLIT distance="250" swimtime="00:08:15.34" />
                    <SPLIT distance="300" swimtime="00:09:30.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-05-28" firstname="Marta" gender="F" lastname="Wolska" nation="POL" athleteid="14798">
              <RESULTS>
                <RESULT eventid="1147" reactiontime="+124" status="OTL" swimtime="00:17:37.87" resultid="14799" heatid="19594" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.24" />
                    <SPLIT distance="100" swimtime="00:01:55.73" />
                    <SPLIT distance="150" swimtime="00:03:02.43" />
                    <SPLIT distance="200" swimtime="00:04:07.75" />
                    <SPLIT distance="250" swimtime="00:05:12.89" />
                    <SPLIT distance="300" swimtime="00:06:18.36" />
                    <SPLIT distance="350" swimtime="00:07:28.06" />
                    <SPLIT distance="400" swimtime="00:08:36.13" />
                    <SPLIT distance="450" swimtime="00:09:43.64" />
                    <SPLIT distance="500" swimtime="00:10:51.31" />
                    <SPLIT distance="550" swimtime="00:12:00.12" />
                    <SPLIT distance="600" swimtime="00:13:09.17" />
                    <SPLIT distance="650" swimtime="00:14:17.25" />
                    <SPLIT distance="700" swimtime="00:15:25.75" />
                    <SPLIT distance="750" swimtime="00:16:35.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="113" reactiontime="+80" swimtime="00:00:53.06" resultid="14800" heatid="19337" lane="2" entrytime="00:00:52.00" entrycourse="SCM" />
                <RESULT eventid="14225" points="112" reactiontime="+125" swimtime="00:01:57.50" resultid="14801" heatid="19390" lane="0" entrytime="00:02:08.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="68" reactiontime="+125" swimtime="00:00:59.60" resultid="14802" heatid="19444" lane="5" />
                <RESULT eventid="1457" points="112" reactiontime="+66" swimtime="00:01:53.90" resultid="14803" heatid="19466" lane="8" entrytime="00:01:52.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="108" reactiontime="+78" swimtime="00:04:10.08" resultid="14804" heatid="19527" lane="9" entrytime="00:04:02.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.07" />
                    <SPLIT distance="100" swimtime="00:02:01.94" />
                    <SPLIT distance="150" swimtime="00:03:06.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="116" reactiontime="+113" swimtime="00:00:58.72" resultid="14805" heatid="19539" lane="5" entrytime="00:00:58.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Karolina" gender="F" lastname="Górka" nation="POL" athleteid="14875">
              <RESULTS>
                <RESULT eventid="1062" points="427" reactiontime="+77" swimtime="00:00:30.84" resultid="14876" heatid="19280" lane="4" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1222" points="339" reactiontime="+80" swimtime="00:03:12.95" resultid="14877" heatid="19357" lane="1" entrytime="00:03:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.01" />
                    <SPLIT distance="100" swimtime="00:01:31.52" />
                    <SPLIT distance="150" swimtime="00:02:21.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="348" reactiontime="+79" swimtime="00:01:20.54" resultid="14878" heatid="19392" lane="0" entrytime="00:01:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="383" reactiontime="+74" swimtime="00:01:25.84" resultid="14879" heatid="19430" lane="5" entrytime="00:01:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="297" reactiontime="+73" swimtime="00:02:45.89" resultid="14880" heatid="19482" lane="7" entrytime="00:03:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                    <SPLIT distance="100" swimtime="00:01:17.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="409" reactiontime="+70" swimtime="00:00:38.56" resultid="14881" heatid="19542" lane="3" entrytime="00:00:42.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-08-01" firstname="Paulina" gender="F" lastname="Palmowska - Latuszek" nation="POL" athleteid="14868">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski " eventid="1165" points="384" reactiontime="+82" swimtime="00:21:05.26" resultid="14869" heatid="19624" lane="4" entrytime="00:21:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.97" />
                    <SPLIT distance="100" swimtime="00:01:16.49" />
                    <SPLIT distance="150" swimtime="00:01:58.30" />
                    <SPLIT distance="200" swimtime="00:02:40.15" />
                    <SPLIT distance="250" swimtime="00:03:22.32" />
                    <SPLIT distance="300" swimtime="00:04:04.74" />
                    <SPLIT distance="350" swimtime="00:04:47.15" />
                    <SPLIT distance="400" swimtime="00:05:29.80" />
                    <SPLIT distance="450" swimtime="00:06:12.16" />
                    <SPLIT distance="500" swimtime="00:06:54.29" />
                    <SPLIT distance="550" swimtime="00:07:36.61" />
                    <SPLIT distance="600" swimtime="00:08:19.23" />
                    <SPLIT distance="650" swimtime="00:09:02.09" />
                    <SPLIT distance="700" swimtime="00:09:44.82" />
                    <SPLIT distance="750" swimtime="00:10:27.33" />
                    <SPLIT distance="800" swimtime="00:11:10.29" />
                    <SPLIT distance="850" swimtime="00:11:52.86" />
                    <SPLIT distance="900" swimtime="00:12:35.89" />
                    <SPLIT distance="950" swimtime="00:13:18.68" />
                    <SPLIT distance="1000" swimtime="00:14:01.42" />
                    <SPLIT distance="1050" swimtime="00:14:43.59" />
                    <SPLIT distance="1100" swimtime="00:15:26.35" />
                    <SPLIT distance="1150" swimtime="00:16:09.11" />
                    <SPLIT distance="1200" swimtime="00:16:52.18" />
                    <SPLIT distance="1250" swimtime="00:17:34.90" />
                    <SPLIT distance="1300" swimtime="00:18:17.22" />
                    <SPLIT distance="1350" swimtime="00:18:59.76" />
                    <SPLIT distance="1400" swimtime="00:19:42.54" />
                    <SPLIT distance="1450" swimtime="00:20:24.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="425" reactiontime="+62" swimtime="00:00:34.13" resultid="14870" heatid="19340" lane="4" entrytime="00:00:34.00" entrycourse="SCM" />
                <RESULT eventid="1457" points="416" reactiontime="+67" swimtime="00:01:13.68" resultid="14871" heatid="19468" lane="4" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="387" reactiontime="+69" swimtime="00:02:31.99" resultid="14872" heatid="19484" lane="7" entrytime="00:02:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.44" />
                    <SPLIT distance="100" swimtime="00:01:09.68" />
                    <SPLIT distance="150" swimtime="00:01:50.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="399" reactiontime="+67" swimtime="00:02:41.83" resultid="14873" heatid="19529" lane="2" entrytime="00:02:37.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                    <SPLIT distance="100" swimtime="00:01:17.92" />
                    <SPLIT distance="150" swimtime="00:02:00.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="14874" heatid="19698" lane="2" entrytime="00:05:15.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" name="Wisła 2" number="2">
              <RESULTS>
                <RESULT eventid="1381" points="128" reactiontime="+89" swimtime="00:02:59.13" resultid="14902" heatid="19421" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.52" />
                    <SPLIT distance="100" swimtime="00:01:36.44" />
                    <SPLIT distance="150" swimtime="00:02:10.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14822" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="14859" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="14894" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="14850" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Wisła 4" number="4">
              <RESULTS>
                <RESULT eventid="1548" status="DNS" swimtime="00:00:00.00" resultid="14904" heatid="19499" lane="0">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14815" number="1" />
                    <RELAYPOSITION athleteid="14782" number="2" />
                    <RELAYPOSITION athleteid="14882" number="3" />
                    <RELAYPOSITION athleteid="14894" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" name="Wisła 1" number="1">
              <RESULTS>
                <RESULT eventid="1358" status="DNS" swimtime="00:00:00.00" resultid="14901" heatid="19419" lane="6">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14842" number="1" />
                    <RELAYPOSITION athleteid="14798" number="2" />
                    <RELAYPOSITION athleteid="14806" number="3" />
                    <RELAYPOSITION athleteid="14888" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="Wisła 3" number="3">
              <RESULTS>
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="14903" heatid="19497" lane="2">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14888" number="1" />
                    <RELAYPOSITION athleteid="14829" number="2" />
                    <RELAYPOSITION athleteid="14806" number="3" />
                    <RELAYPOSITION athleteid="14868" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="Wisła 5" number="5">
              <RESULTS>
                <RESULT eventid="1698" status="DNS" swimtime="00:00:00.00" resultid="14905" heatid="19561" lane="5">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14829" number="1" />
                    <RELAYPOSITION athleteid="14798" number="2" />
                    <RELAYPOSITION athleteid="14815" number="3" />
                    <RELAYPOSITION athleteid="14782" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="15864" name="MASTERS Zdzieszowice">
          <CONTACT email="masters.zdzieszowice@gmail.com" name="Jajuga" phone="505127695" />
          <ATHLETES>
            <ATHLETE birthdate="1973-08-18" firstname="Dorota" gender="F" lastname="Woźniak" nation="POL" athleteid="15881">
              <RESULTS>
                <RESULT eventid="1096" points="327" reactiontime="+87" swimtime="00:02:56.74" resultid="15882" heatid="19308" lane="8" entrytime="00:02:59.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.32" />
                    <SPLIT distance="100" swimtime="00:01:22.81" />
                    <SPLIT distance="150" swimtime="00:02:14.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="337" reactiontime="+107" swimtime="00:01:21.36" resultid="15883" heatid="19393" lane="3" entrytime="00:01:23.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="247" reactiontime="+109" swimtime="00:03:10.55" resultid="15884" heatid="19412" lane="5" entrytime="00:03:10.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.61" />
                    <SPLIT distance="100" swimtime="00:01:31.61" />
                    <SPLIT distance="150" swimtime="00:02:21.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="324" reactiontime="+74" swimtime="00:01:20.10" resultid="15885" heatid="19468" lane="0" entrytime="00:01:23.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="328" reactiontime="+77" swimtime="00:02:52.83" resultid="15886" heatid="19528" lane="4" entrytime="00:02:56.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.68" />
                    <SPLIT distance="100" swimtime="00:01:23.92" />
                    <SPLIT distance="150" swimtime="00:02:08.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="290" reactiontime="+114" swimtime="00:05:54.27" resultid="15887" heatid="19697" lane="2" entrytime="00:06:00.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.28" />
                    <SPLIT distance="100" swimtime="00:01:25.67" />
                    <SPLIT distance="150" swimtime="00:02:10.94" />
                    <SPLIT distance="200" swimtime="00:02:56.56" />
                    <SPLIT distance="250" swimtime="00:03:41.70" />
                    <SPLIT distance="300" swimtime="00:04:26.70" />
                    <SPLIT distance="350" swimtime="00:05:11.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-10" firstname="Dawid" gender="M" lastname="Jajuga" nation="POL" athleteid="15895">
              <RESULTS>
                <RESULT eventid="1113" points="487" reactiontime="+84" swimtime="00:02:19.30" resultid="15896" heatid="19318" lane="1" entrytime="00:02:18.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.08" />
                    <SPLIT distance="100" swimtime="00:01:05.83" />
                    <SPLIT distance="150" swimtime="00:01:46.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14189" status="DNS" swimtime="00:00:00.00" resultid="15897" heatid="19617" lane="8" entrytime="00:10:20.00" />
                <RESULT eventid="14243" points="488" reactiontime="+84" swimtime="00:01:03.85" resultid="15898" heatid="19409" lane="2" entrytime="00:01:03.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="428" reactiontime="+80" swimtime="00:02:23.97" resultid="15899" heatid="19418" lane="7" entrytime="00:02:22.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                    <SPLIT distance="100" swimtime="00:01:09.33" />
                    <SPLIT distance="150" swimtime="00:01:48.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="15900" heatid="19463" lane="8" entrytime="00:00:27.05" />
                <RESULT eventid="1578" points="451" reactiontime="+82" swimtime="00:05:07.02" resultid="15901" heatid="19512" lane="7" entrytime="00:05:05.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                    <SPLIT distance="100" swimtime="00:01:10.97" />
                    <SPLIT distance="150" swimtime="00:01:51.77" />
                    <SPLIT distance="200" swimtime="00:02:31.39" />
                    <SPLIT distance="250" swimtime="00:03:15.04" />
                    <SPLIT distance="300" swimtime="00:03:57.95" />
                    <SPLIT distance="350" swimtime="00:04:33.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="470" reactiontime="+70" swimtime="00:01:01.80" resultid="15902" heatid="19525" lane="9" entrytime="00:01:00.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="497" reactiontime="+81" swimtime="00:00:31.86" resultid="15903" heatid="19558" lane="3" entrytime="00:00:32.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-12-10" firstname="Ewelina" gender="F" lastname="Cuch" nation="POL" athleteid="15865">
              <RESULTS>
                <RESULT eventid="1256" points="290" reactiontime="+79" swimtime="00:01:16.86" resultid="15866" heatid="19371" lane="8" entrytime="00:01:14.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="303" reactiontime="+90" swimtime="00:01:24.29" resultid="15867" heatid="19393" lane="8" entrytime="00:01:25.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="267" reactiontime="+101" swimtime="00:02:51.98" resultid="15868" heatid="19482" lane="2" entrytime="00:02:59.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.60" />
                    <SPLIT distance="100" swimtime="00:01:23.23" />
                    <SPLIT distance="150" swimtime="00:02:07.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="226" reactiontime="+96" swimtime="00:07:05.78" resultid="15869" heatid="19503" lane="4" entrytime="00:07:20.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.85" />
                    <SPLIT distance="100" swimtime="00:01:25.02" />
                    <SPLIT distance="150" swimtime="00:02:24.64" />
                    <SPLIT distance="200" swimtime="00:03:23.76" />
                    <SPLIT distance="250" swimtime="00:04:24.27" />
                    <SPLIT distance="300" swimtime="00:05:25.72" />
                    <SPLIT distance="350" swimtime="00:06:16.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="271" reactiontime="+85" swimtime="00:01:24.35" resultid="15870" heatid="19514" lane="5" entrytime="00:01:25.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="266" reactiontime="+91" swimtime="00:06:04.30" resultid="15871" heatid="19697" lane="7" entrytime="00:06:11.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.93" />
                    <SPLIT distance="100" swimtime="00:01:25.47" />
                    <SPLIT distance="150" swimtime="00:02:11.29" />
                    <SPLIT distance="200" swimtime="00:02:57.99" />
                    <SPLIT distance="250" swimtime="00:03:45.11" />
                    <SPLIT distance="300" swimtime="00:04:31.02" />
                    <SPLIT distance="350" swimtime="00:05:17.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-10-02" firstname="Szymon" gender="M" lastname="Paciej" nation="POL" athleteid="15888">
              <RESULTS>
                <RESULT eventid="1113" points="384" reactiontime="+86" swimtime="00:02:30.77" resultid="15889" heatid="19316" lane="4" entrytime="00:02:29.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                    <SPLIT distance="100" swimtime="00:01:11.00" />
                    <SPLIT distance="150" swimtime="00:01:55.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="360" reactiontime="+87" swimtime="00:02:49.26" resultid="15890" heatid="19363" lane="7" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.11" />
                    <SPLIT distance="100" swimtime="00:01:21.91" />
                    <SPLIT distance="150" swimtime="00:02:06.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="280" reactiontime="+87" swimtime="00:02:45.79" resultid="15891" heatid="19417" lane="6" entrytime="00:02:43.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="100" swimtime="00:01:15.58" />
                    <SPLIT distance="150" swimtime="00:01:59.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="328" reactiontime="+83" swimtime="00:01:10.89" resultid="15892" heatid="19477" lane="7" entrytime="00:01:08.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="352" reactiontime="+92" swimtime="00:05:33.41" resultid="15893" heatid="19511" lane="2" entrytime="00:05:30.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                    <SPLIT distance="100" swimtime="00:01:15.69" />
                    <SPLIT distance="150" swimtime="00:01:57.35" />
                    <SPLIT distance="200" swimtime="00:02:39.48" />
                    <SPLIT distance="250" swimtime="00:03:27.20" />
                    <SPLIT distance="300" swimtime="00:04:14.84" />
                    <SPLIT distance="350" swimtime="00:04:55.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="323" reactiontime="+92" swimtime="00:02:33.86" resultid="15894" heatid="19536" lane="0" entrytime="00:02:40.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                    <SPLIT distance="100" swimtime="00:01:13.64" />
                    <SPLIT distance="150" swimtime="00:01:53.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-08" firstname="Przemysław" gender="M" lastname="Osiwała" nation="POL" athleteid="15904">
              <RESULTS>
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="15905" heatid="19313" lane="3" entrytime="00:02:45.87" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="15906" heatid="19362" lane="3" entrytime="00:03:05.67" />
                <RESULT eventid="1341" points="311" reactiontime="+91" swimtime="00:02:40.19" resultid="15907" heatid="19416" lane="5" entrytime="00:02:50.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                    <SPLIT distance="100" swimtime="00:01:16.86" />
                    <SPLIT distance="150" swimtime="00:01:57.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="15908" heatid="19457" lane="4" entrytime="00:00:31.33" />
                <RESULT eventid="1578" points="272" reactiontime="+93" swimtime="00:06:03.42" resultid="15909" heatid="19510" lane="9" entrytime="00:06:05.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                    <SPLIT distance="100" swimtime="00:01:20.60" />
                    <SPLIT distance="150" swimtime="00:02:09.02" />
                    <SPLIT distance="200" swimtime="00:02:57.78" />
                    <SPLIT distance="250" swimtime="00:03:51.01" />
                    <SPLIT distance="300" swimtime="00:04:43.33" />
                    <SPLIT distance="350" swimtime="00:05:24.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="15910" heatid="19522" lane="3" entrytime="00:01:09.22" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="15911" heatid="19555" lane="9" entrytime="00:00:36.55" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-08-23" firstname="Katarzyna" gender="F" lastname="Gniot" nation="POL" athleteid="15872">
              <RESULTS>
                <RESULT eventid="1062" points="241" swimtime="00:00:37.34" resultid="15873" heatid="19278" lane="0" entrytime="00:00:39.76" />
                <RESULT eventid="1096" points="156" reactiontime="+119" swimtime="00:03:46.31" resultid="15874" heatid="19307" lane="4" entrytime="00:03:00.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.42" />
                    <SPLIT distance="100" swimtime="00:01:50.52" />
                    <SPLIT distance="150" swimtime="00:02:54.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="138" reactiontime="+95" swimtime="00:00:49.63" resultid="15875" heatid="19339" lane="0" entrytime="00:00:40.98" />
                <RESULT eventid="1222" points="172" reactiontime="+112" swimtime="00:04:01.77" resultid="15876" heatid="19356" lane="1" entrytime="00:03:50.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.19" />
                    <SPLIT distance="100" swimtime="00:01:54.68" />
                    <SPLIT distance="150" swimtime="00:02:57.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="189" reactiontime="+126" swimtime="00:01:48.64" resultid="15877" heatid="19428" lane="2" entrytime="00:01:56.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="134" reactiontime="+82" swimtime="00:01:47.33" resultid="15878" heatid="19466" lane="6" entrytime="00:01:35.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="139" reactiontime="+83" swimtime="00:03:50.09" resultid="15879" heatid="19526" lane="4" entrytime="00:04:10.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.00" />
                    <SPLIT distance="100" swimtime="00:01:50.58" />
                    <SPLIT distance="150" swimtime="00:02:50.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="217" reactiontime="+106" swimtime="00:00:47.63" resultid="15880" heatid="19540" lane="2" entrytime="00:00:51.23" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="339" reactiontime="+77" swimtime="00:02:06.90" resultid="15912" heatid="19320" lane="4" entrytime="00:02:10.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.13" />
                    <SPLIT distance="100" swimtime="00:01:05.08" />
                    <SPLIT distance="150" swimtime="00:01:38.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15895" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="15872" number="2" reactiontime="+78" />
                    <RELAYPOSITION athleteid="15881" number="3" reactiontime="+99" />
                    <RELAYPOSITION athleteid="15888" number="4" reactiontime="+73" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="373" reactiontime="+74" swimtime="00:02:14.94" resultid="15913" heatid="19563" lane="1" entrytime="00:02:20.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.82" />
                    <SPLIT distance="100" swimtime="00:01:13.03" />
                    <SPLIT distance="150" swimtime="00:01:49.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15881" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="15888" number="2" reactiontime="+76" />
                    <RELAYPOSITION athleteid="15865" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="15895" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="16777" name="Masters Łódź">
          <CONTACT email="sport@masterslodz.pl" internet="http://masterslodz.pl" name="Trudnos Rafał" phone="604184311" />
          <ATHLETES>
            <ATHLETE birthdate="1978-03-01" firstname="Marek" gender="M" lastname="Gurbski" nation="POL" athleteid="16844">
              <RESULTS>
                <RESULT eventid="1079" points="297" reactiontime="+92" swimtime="00:00:30.36" resultid="16845" heatid="19290" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="1205" points="234" reactiontime="+68" swimtime="00:00:36.02" resultid="16846" heatid="19346" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="14243" points="250" reactiontime="+95" swimtime="00:01:19.79" resultid="16847" heatid="19401" lane="8" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="279" reactiontime="+86" swimtime="00:00:33.34" resultid="16848" heatid="19455" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="1681" points="242" reactiontime="+94" swimtime="00:00:40.47" resultid="16849" heatid="19551" lane="5" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-16" firstname="Jakub" gender="M" lastname="Karczmarczyk" nation="POL" athleteid="16855">
              <RESULTS>
                <RESULT eventid="1079" points="343" swimtime="00:00:28.93" resultid="16856" heatid="19285" lane="9" entrytime="00:00:45.00" />
                <RESULT eventid="1113" points="234" reactiontime="+101" swimtime="00:02:57.66" resultid="16857" heatid="19311" lane="6" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.91" />
                    <SPLIT distance="100" swimtime="00:01:22.74" />
                    <SPLIT distance="150" swimtime="00:02:15.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="16858" heatid="19361" lane="1" entrytime="00:03:30.00" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="16859" heatid="19436" lane="2" entrytime="00:01:35.00" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="16860" heatid="19506" lane="5" />
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="16861" heatid="19534" lane="8" entrytime="00:03:15.00" />
                <RESULT eventid="1681" points="268" reactiontime="+96" swimtime="00:00:39.15" resultid="16862" heatid="19549" lane="5" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-02" firstname="Wojciech" gender="M" lastname="Zdzieszyński" nation="POL" athleteid="16850">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="16851" heatid="19299" lane="7" entrytime="00:00:27.00" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="16852" heatid="19381" lane="3" entrytime="00:01:06.00" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="16853" heatid="19455" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="16854" heatid="19555" lane="2" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-16" firstname="Joanna" gender="F" lastname="Wilińska" nation="POL" athleteid="16793">
              <RESULTS>
                <RESULT eventid="1423" points="405" reactiontime="+100" swimtime="00:00:32.94" resultid="16794" heatid="19448" lane="4" entrytime="00:00:32.50" />
                <RESULT eventid="1595" points="406" reactiontime="+101" swimtime="00:01:13.75" resultid="16795" heatid="19515" lane="1" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-06-12" firstname="Igor" gender="M" lastname="Olejarczyk" nation="POL" athleteid="16796">
              <RESULTS>
                <RESULT eventid="1079" points="460" reactiontime="+67" swimtime="00:00:26.24" resultid="16797" heatid="19300" lane="8" entrytime="00:00:26.50" />
                <RESULT eventid="1273" points="437" reactiontime="+75" swimtime="00:00:59.22" resultid="16798" heatid="19385" lane="2" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" status="DNS" swimtime="00:00:00.00" resultid="16799" heatid="19417" lane="9" entrytime="00:02:50.00" />
                <RESULT eventid="1440" points="411" reactiontime="+72" swimtime="00:00:29.31" resultid="16800" heatid="19461" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="1613" points="405" reactiontime="+77" swimtime="00:01:04.98" resultid="16801" heatid="19523" lane="2" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-06-28" firstname="Artur" gender="M" lastname="Frąckowiak" nation="POL" athleteid="16822">
              <RESULTS>
                <RESULT eventid="1079" points="440" reactiontime="+85" swimtime="00:00:26.62" resultid="16823" heatid="19286" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1113" points="417" reactiontime="+84" swimtime="00:02:26.70" resultid="16824" heatid="19315" lane="7" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.60" />
                    <SPLIT distance="100" swimtime="00:01:09.51" />
                    <SPLIT distance="150" swimtime="00:01:53.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="443" reactiontime="+80" swimtime="00:00:58.92" resultid="16825" heatid="19385" lane="9" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="426" reactiontime="+84" swimtime="00:00:28.97" resultid="16826" heatid="19459" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1508" points="420" reactiontime="+86" swimtime="00:02:12.59" resultid="16827" heatid="19494" lane="6" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.16" />
                    <SPLIT distance="100" swimtime="00:01:03.16" />
                    <SPLIT distance="150" swimtime="00:01:37.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="16828" heatid="19706" lane="7" entrytime="00:05:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-09" firstname="Marcin" gender="M" lastname="Strąkowski" nation="POL" athleteid="16814">
              <RESULTS>
                <RESULT eventid="1079" points="331" reactiontime="+94" swimtime="00:00:29.28" resultid="16815" heatid="19296" lane="2" entrytime="00:00:28.60" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="16816" heatid="19381" lane="0" entrytime="00:01:07.80" />
                <RESULT eventid="1681" points="263" reactiontime="+98" swimtime="00:00:39.41" resultid="16817" heatid="19553" lane="2" entrytime="00:00:37.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-04-28" firstname="Kornel" gender="M" lastname="Pintara" nation="POL" athleteid="16808">
              <RESULTS>
                <RESULT eventid="1079" points="450" reactiontime="+79" swimtime="00:00:26.43" resultid="16809" heatid="19295" lane="3" entrytime="00:00:29.00" />
                <RESULT eventid="14243" points="286" reactiontime="+94" swimtime="00:01:16.31" resultid="16810" heatid="19401" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="321" reactiontime="+85" swimtime="00:00:31.83" resultid="16811" heatid="19458" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="1508" points="261" reactiontime="+107" swimtime="00:02:35.38" resultid="16812" heatid="19491" lane="1" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.62" />
                    <SPLIT distance="100" swimtime="00:01:15.59" />
                    <SPLIT distance="150" swimtime="00:01:55.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="261" reactiontime="+88" swimtime="00:00:39.47" resultid="16813" heatid="19550" lane="0" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-15" firstname="Arkadiusz" gender="M" lastname="Olkowicz" nation="POL" athleteid="16835">
              <RESULTS>
                <RESULT eventid="1079" points="286" reactiontime="+83" swimtime="00:00:30.72" resultid="16836" heatid="19292" lane="2" entrytime="00:00:30.10" />
                <RESULT eventid="14189" points="293" reactiontime="+89" swimtime="00:11:07.00" resultid="16837" heatid="19616" lane="6" entrytime="00:11:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.99" />
                    <SPLIT distance="100" swimtime="00:01:16.47" />
                    <SPLIT distance="150" swimtime="00:01:56.46" />
                    <SPLIT distance="200" swimtime="00:02:37.80" />
                    <SPLIT distance="250" swimtime="00:03:19.03" />
                    <SPLIT distance="300" swimtime="00:04:00.77" />
                    <SPLIT distance="350" swimtime="00:04:42.88" />
                    <SPLIT distance="400" swimtime="00:05:25.10" />
                    <SPLIT distance="450" swimtime="00:06:08.12" />
                    <SPLIT distance="500" swimtime="00:06:50.90" />
                    <SPLIT distance="550" swimtime="00:07:33.76" />
                    <SPLIT distance="600" swimtime="00:08:16.75" />
                    <SPLIT distance="650" swimtime="00:09:00.37" />
                    <SPLIT distance="700" swimtime="00:09:43.42" />
                    <SPLIT distance="750" swimtime="00:10:26.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="223" reactiontime="+85" swimtime="00:00:36.60" resultid="16838" heatid="19350" lane="1" entrytime="00:00:32.50" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="16839" heatid="19381" lane="7" entrytime="00:01:06.50" />
                <RESULT eventid="1440" points="305" reactiontime="+82" swimtime="00:00:32.38" resultid="16840" heatid="19458" lane="9" entrytime="00:00:31.10" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="16841" heatid="19492" lane="0" entrytime="00:02:27.70" />
                <RESULT eventid="1647" reactiontime="+51" status="DNS" swimtime="00:00:00.00" resultid="16842" heatid="19534" lane="9" entrytime="00:03:17.70" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="16843" heatid="19703" lane="6" entrytime="00:05:51.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-14" firstname="Damian" gender="M" lastname="Karkusiński" nation="POL" athleteid="16818">
              <RESULTS>
                <RESULT eventid="1079" points="306" reactiontime="+89" swimtime="00:00:30.06" resultid="16819" heatid="19294" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="1205" points="228" reactiontime="+69" swimtime="00:00:36.35" resultid="16820" heatid="19349" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="16821" heatid="19475" lane="5" entrytime="00:01:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-08-10" firstname="Błażej" gender="M" lastname="Dunajczyk" nation="POL" athleteid="16832">
              <RESULTS>
                <RESULT eventid="1079" points="358" reactiontime="+85" swimtime="00:00:28.51" resultid="16833" heatid="19292" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1440" points="293" reactiontime="+94" swimtime="00:00:32.81" resultid="16834" heatid="19457" lane="1" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-02-14" firstname="Jakub" gender="M" lastname="Gryczyński" nation="POL" athleteid="16873">
              <RESULTS>
                <RESULT eventid="1079" points="263" reactiontime="+96" swimtime="00:00:31.59" resultid="16874" heatid="19290" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="14243" status="DNS" swimtime="00:00:00.00" resultid="16875" heatid="19400" lane="8" entrytime="00:01:30.00" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="16876" heatid="19437" lane="1" entrytime="00:01:30.00" />
                <RESULT eventid="1681" points="251" reactiontime="+97" swimtime="00:00:40.00" resultid="16877" heatid="19552" lane="2" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-08-19" firstname="Łukasz" gender="M" lastname="Raj" nation="POL" athleteid="16868">
              <RESULTS>
                <RESULT eventid="1079" points="269" reactiontime="+86" swimtime="00:00:31.38" resultid="16869" heatid="19291" lane="7" entrytime="00:00:31.50" />
                <RESULT eventid="14243" status="DNS" swimtime="00:00:00.00" resultid="16870" heatid="19401" lane="6" entrytime="00:01:24.33" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="16871" heatid="19438" lane="8" entrytime="00:01:27.11" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="16872" heatid="19551" lane="4" entrytime="00:00:39.98" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-11-02" firstname="Ksawery" gender="M" lastname="Wiaderek" nation="POL" athleteid="16863">
              <RESULTS>
                <RESULT eventid="1079" points="433" reactiontime="+87" swimtime="00:00:26.77" resultid="16864" heatid="19301" lane="7" entrytime="00:00:26.00" />
                <RESULT eventid="1205" points="301" reactiontime="+83" swimtime="00:00:33.13" resultid="16865" heatid="19349" lane="1" entrytime="00:00:34.00" />
                <RESULT eventid="1273" points="367" reactiontime="+92" swimtime="00:01:02.74" resultid="16866" heatid="19385" lane="8" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="396" reactiontime="+93" swimtime="00:00:29.67" resultid="16867" heatid="19461" lane="6" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-03-14" firstname="Anna" gender="F" lastname="Ostrowska" nation="POL" athleteid="16829">
              <RESULTS>
                <RESULT eventid="1062" points="427" reactiontime="+88" swimtime="00:00:30.86" resultid="16830" heatid="19282" lane="6" entrytime="00:00:30.20" />
                <RESULT eventid="1256" points="370" reactiontime="+86" swimtime="00:01:10.86" resultid="16831" heatid="19370" lane="7" entrytime="00:01:15.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-09-18" firstname="Konrad" gender="M" lastname="Hasik" nation="POL" athleteid="16878">
              <RESULTS>
                <RESULT eventid="1113" points="447" reactiontime="+86" swimtime="00:02:23.38" resultid="16879" heatid="19314" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.34" />
                    <SPLIT distance="100" swimtime="00:01:07.75" />
                    <SPLIT distance="150" swimtime="00:01:49.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="431" reactiontime="+63" swimtime="00:00:29.40" resultid="16880" heatid="19352" lane="6" entrytime="00:00:29.00" />
                <RESULT eventid="1341" status="DNS" swimtime="00:00:00.00" resultid="16881" heatid="19416" lane="2" entrytime="00:03:00.00" />
                <RESULT eventid="1474" points="449" reactiontime="+64" swimtime="00:01:03.88" resultid="16882" heatid="19478" lane="8" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="16883" heatid="19510" lane="8" entrytime="00:06:00.00" />
                <RESULT eventid="1647" points="386" swimtime="00:02:25.02" resultid="16884" heatid="19535" lane="8" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                    <SPLIT distance="100" swimtime="00:01:10.42" />
                    <SPLIT distance="150" swimtime="00:01:48.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="16885" heatid="19557" lane="0" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-09" firstname="Rafał" gender="M" lastname="Trudnos" nation="POL" athleteid="16802">
              <RESULTS>
                <RESULT eventid="1079" points="392" reactiontime="+80" swimtime="00:00:27.66" resultid="16803" heatid="19299" lane="6" entrytime="00:00:27.00" />
                <RESULT eventid="1239" points="402" reactiontime="+80" swimtime="00:02:43.11" resultid="16804" heatid="19364" lane="8" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.48" />
                    <SPLIT distance="100" swimtime="00:01:17.07" />
                    <SPLIT distance="150" swimtime="00:01:59.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="425" reactiontime="+79" swimtime="00:01:13.93" resultid="16805" heatid="19441" lane="9" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="400" reactiontime="+81" swimtime="00:00:29.57" resultid="16806" heatid="19459" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1681" points="466" reactiontime="+85" swimtime="00:00:32.55" resultid="16807" heatid="19557" lane="2" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1381" points="459" swimtime="00:01:57.28" resultid="16888" heatid="19424" lane="1" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.55" />
                    <SPLIT distance="100" swimtime="00:01:02.26" />
                    <SPLIT distance="150" swimtime="00:01:30.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16878" number="1" />
                    <RELAYPOSITION athleteid="16802" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="16796" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="16863" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1381" points="297" reactiontime="+78" swimtime="00:02:15.58" resultid="16889" heatid="19423" lane="1" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                    <SPLIT distance="100" swimtime="00:01:15.94" />
                    <SPLIT distance="150" swimtime="00:01:45.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16835" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="16855" number="2" reactiontime="+91" />
                    <RELAYPOSITION athleteid="16822" number="3" reactiontime="+65" />
                    <RELAYPOSITION athleteid="16814" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="1381" points="290" reactiontime="+62" swimtime="00:02:16.70" resultid="16890" heatid="19423" lane="9" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.90" />
                    <SPLIT distance="100" swimtime="00:01:15.68" />
                    <SPLIT distance="150" swimtime="00:01:48.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16818" number="1" reactiontime="+62" />
                    <RELAYPOSITION athleteid="16873" number="2" reactiontime="+33" />
                    <RELAYPOSITION athleteid="16808" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="16832" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="6">
              <RESULTS>
                <RESULT eventid="1548" points="460" reactiontime="+67" swimtime="00:01:46.95" resultid="16891" heatid="19502" lane="7" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.59" />
                    <SPLIT distance="100" swimtime="00:00:52.67" />
                    <SPLIT distance="150" swimtime="00:01:19.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16796" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="16878" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="16822" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="16863" number="4" reactiontime="+16" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="7">
              <RESULTS>
                <RESULT eventid="1548" points="375" reactiontime="+87" swimtime="00:01:54.52" resultid="16892" heatid="19502" lane="8" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.02" />
                    <SPLIT distance="100" swimtime="00:00:56.64" />
                    <SPLIT distance="150" swimtime="00:01:26.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16808" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="16802" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="16814" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="16832" number="4" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="8">
              <RESULTS>
                <RESULT eventid="1548" points="328" reactiontime="+83" swimtime="00:01:59.66" resultid="16893" heatid="19501" lane="0" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                    <SPLIT distance="100" swimtime="00:00:59.76" />
                    <SPLIT distance="150" swimtime="00:01:29.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16818" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="16835" number="2" reactiontime="+21" />
                    <RELAYPOSITION athleteid="16844" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="16855" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="474" reactiontime="+83" swimtime="00:01:53.56" resultid="16886" heatid="19322" lane="3" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.40" />
                    <SPLIT distance="100" swimtime="00:00:57.04" />
                    <SPLIT distance="150" swimtime="00:01:27.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16796" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="16829" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="16793" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="16863" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1698" points="480" reactiontime="+69" swimtime="00:02:04.06" resultid="16887" heatid="19564" lane="5" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                    <SPLIT distance="100" swimtime="00:01:01.38" />
                    <SPLIT distance="150" swimtime="00:01:33.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16878" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="16802" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="16793" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="16829" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MASTKRAS" nation="POL" region="LBL" clubid="16225" name="Masterskrasnik">
          <CONTACT city="Krasnik" email="masterskrasnik@gmail.com" internet="www.masterskrasnik.za.pl" name="Michalczyk" phone="601698977" state="LUB" street="Żwirki i Wigury 2" zip="23-200" />
          <ATHLETES>
            <ATHLETE birthdate="1960-09-07" firstname="Andrzej" gender="M" lastname="Cis" nation="POL" athleteid="16226">
              <RESULTS>
                <RESULT eventid="1079" points="278" reactiontime="+74" swimtime="00:00:31.04" resultid="16227" heatid="19290" lane="7" entrytime="00:00:32.10" />
                <RESULT eventid="14189" points="148" reactiontime="+85" swimtime="00:13:56.74" resultid="16228" heatid="19615" lane="3" entrytime="00:14:10.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.52" />
                    <SPLIT distance="100" swimtime="00:01:27.65" />
                    <SPLIT distance="150" swimtime="00:02:17.12" />
                    <SPLIT distance="200" swimtime="00:03:08.22" />
                    <SPLIT distance="250" swimtime="00:04:00.69" />
                    <SPLIT distance="300" swimtime="00:04:54.52" />
                    <SPLIT distance="350" swimtime="00:05:50.16" />
                    <SPLIT distance="400" swimtime="00:06:44.62" />
                    <SPLIT distance="450" swimtime="00:07:38.00" />
                    <SPLIT distance="500" swimtime="00:08:30.40" />
                    <SPLIT distance="550" swimtime="00:09:24.30" />
                    <SPLIT distance="600" swimtime="00:10:17.33" />
                    <SPLIT distance="650" swimtime="00:11:10.54" />
                    <SPLIT distance="700" swimtime="00:12:05.67" />
                    <SPLIT distance="750" swimtime="00:13:04.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="187" reactiontime="+73" swimtime="00:00:38.81" resultid="16229" heatid="19347" lane="1" entrytime="00:00:38.20" />
                <RESULT eventid="1341" points="85" reactiontime="+92" swimtime="00:04:06.30" resultid="16230" heatid="19414" lane="6" entrytime="00:04:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.63" />
                    <SPLIT distance="100" swimtime="00:01:59.50" />
                    <SPLIT distance="150" swimtime="00:03:04.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="16231" heatid="19474" lane="0" entrytime="00:01:26.00" />
                <RESULT eventid="1578" points="134" reactiontime="+73" swimtime="00:07:39.23" resultid="16232" heatid="19508" lane="0" entrytime="00:07:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.00" />
                    <SPLIT distance="100" swimtime="00:01:55.31" />
                    <SPLIT distance="150" swimtime="00:02:54.53" />
                    <SPLIT distance="200" swimtime="00:03:55.29" />
                    <SPLIT distance="250" swimtime="00:05:00.52" />
                    <SPLIT distance="300" swimtime="00:06:04.08" />
                    <SPLIT distance="350" swimtime="00:06:55.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="92" reactiontime="+80" swimtime="00:01:46.38" resultid="16233" heatid="19518" lane="6" entrytime="00:01:38.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="16234" heatid="19705" lane="3" entrytime="00:05:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-11-05" firstname="Krzysztof" gender="M" lastname="Samonek" nation="POL" athleteid="16243">
              <RESULTS>
                <RESULT eventid="1079" points="94" swimtime="00:00:44.47" resultid="16244" heatid="19286" lane="9" entrytime="00:00:40.20" />
                <RESULT eventid="1113" points="101" reactiontime="+108" swimtime="00:03:55.35" resultid="16245" heatid="19310" lane="6" entrytime="00:04:04.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.54" />
                    <SPLIT distance="100" swimtime="00:01:51.89" />
                    <SPLIT distance="150" swimtime="00:03:03.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="112" reactiontime="+72" swimtime="00:00:45.97" resultid="16246" heatid="19345" lane="9" entrytime="00:00:48.35" />
                <RESULT eventid="14243" points="116" reactiontime="+113" swimtime="00:01:43.12" resultid="16247" heatid="19398" lane="5" entrytime="00:01:49.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="95" reactiontime="+90" swimtime="00:01:47.10" resultid="16248" heatid="19472" lane="0" entrytime="00:01:51.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="16249" heatid="19507" lane="3" entrytime="00:08:40.30" />
                <RESULT eventid="1647" points="102" reactiontime="+85" swimtime="00:03:45.78" resultid="16250" heatid="19532" lane="3" entrytime="00:04:03.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.34" />
                    <SPLIT distance="100" swimtime="00:02:52.63" />
                    <SPLIT distance="150" swimtime="00:03:45.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-09" firstname="Jerzy" gender="M" lastname="Michalczyk" nation="POL" athleteid="16251">
              <RESULTS>
                <RESULT eventid="1079" points="98" reactiontime="+102" swimtime="00:00:43.89" resultid="16252" heatid="19285" lane="1" entrytime="00:00:45.00" />
                <RESULT eventid="1205" points="77" reactiontime="+95" swimtime="00:00:52.20" resultid="16253" heatid="19344" lane="0" entrytime="00:00:55.00" />
                <RESULT eventid="1273" points="104" reactiontime="+97" swimtime="00:01:35.53" resultid="16254" heatid="19374" lane="5" entrytime="00:01:45.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="105" reactiontime="+95" swimtime="00:01:57.70" resultid="16255" heatid="19435" lane="8" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="81" reactiontime="+99" swimtime="00:00:50.28" resultid="16256" heatid="19451" lane="7" entrytime="00:00:55.00" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="16257" heatid="19517" lane="6" entrytime="00:01:58.30" />
                <RESULT eventid="1681" points="119" reactiontime="+96" swimtime="00:00:51.29" resultid="16258" heatid="19548" lane="0" entrytime="00:00:58.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-08-17" firstname="Jacek" gender="M" lastname="Janik" nation="POL" athleteid="16235">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="16236" heatid="19288" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="16237" heatid="19360" lane="6" entrytime="00:03:54.47" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="16238" heatid="19377" lane="6" entrytime="00:01:20.00" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="16239" heatid="19436" lane="9" entrytime="00:01:44.00" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="16240" heatid="19488" lane="9" entrytime="00:03:10.00" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="16241" heatid="19550" lane="6" entrytime="00:00:44.00" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="16242" heatid="19700" lane="0" entrytime="00:07:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="18592" name="MIŁEK TRIATHLON TEAM">
          <ATHLETES>
            <ATHLETE birthdate="1987-12-13" firstname="Mateusz" gender="M" lastname="Miłek" nation="POL" athleteid="18583">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="18584" heatid="19300" lane="0" entrytime="00:00:26.50" />
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="18585" heatid="19316" lane="2" entrytime="00:02:30.00" />
                <RESULT eventid="1205" points="409" reactiontime="+74" swimtime="00:00:29.92" resultid="18586" heatid="19352" lane="1" entrytime="00:00:29.50" />
                <RESULT eventid="1341" points="328" reactiontime="+83" swimtime="00:02:37.35" resultid="18587" heatid="19417" lane="3" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                    <SPLIT distance="100" swimtime="00:01:13.50" />
                    <SPLIT distance="150" swimtime="00:01:55.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="465" reactiontime="+78" swimtime="00:00:28.12" resultid="18588" heatid="19462" lane="0" entrytime="00:00:27.80" />
                <RESULT eventid="1474" points="341" reactiontime="+76" swimtime="00:01:10.02" resultid="18589" heatid="19477" lane="6" entrytime="00:01:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="18590" heatid="19524" lane="8" entrytime="00:01:04.50" />
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="18591" heatid="19537" lane="0" entrytime="00:02:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00308" nation="POL" region="PDK" clubid="16524" name="MKP Bobry Dębica">
          <CONTACT name="GOGACZ" phone="506694816" />
          <ATHLETES>
            <ATHLETE birthdate="1976-10-28" firstname="Sebastian" gender="M" lastname="Gogacz" nation="POL" athleteid="16525">
              <RESULTS>
                <RESULT eventid="14189" points="362" reactiontime="+93" status="EXH" swimtime="00:10:22.14" resultid="16526" heatid="19617" lane="0" entrytime="00:10:22.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                    <SPLIT distance="100" swimtime="00:01:14.00" />
                    <SPLIT distance="150" swimtime="00:01:53.40" />
                    <SPLIT distance="200" swimtime="00:02:32.53" />
                    <SPLIT distance="250" swimtime="00:03:11.96" />
                    <SPLIT distance="300" swimtime="00:03:51.36" />
                    <SPLIT distance="350" swimtime="00:04:30.54" />
                    <SPLIT distance="400" swimtime="00:05:09.87" />
                    <SPLIT distance="450" swimtime="00:05:49.45" />
                    <SPLIT distance="500" swimtime="00:06:27.93" />
                    <SPLIT distance="550" swimtime="00:07:06.70" />
                    <SPLIT distance="600" swimtime="00:07:45.67" />
                    <SPLIT distance="650" swimtime="00:08:24.77" />
                    <SPLIT distance="700" swimtime="00:09:03.85" />
                    <SPLIT distance="750" swimtime="00:09:42.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14207" points="367" reactiontime="+84" swimtime="00:19:44.30" resultid="16527" heatid="19623" lane="0" entrytime="00:20:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.26" />
                    <SPLIT distance="100" swimtime="00:01:12.62" />
                    <SPLIT distance="200" swimtime="00:02:30.25" />
                    <SPLIT distance="250" swimtime="00:03:09.72" />
                    <SPLIT distance="300" swimtime="00:03:48.97" />
                    <SPLIT distance="350" swimtime="00:04:28.02" />
                    <SPLIT distance="400" swimtime="00:05:07.23" />
                    <SPLIT distance="450" swimtime="00:05:47.19" />
                    <SPLIT distance="500" swimtime="00:06:26.43" />
                    <SPLIT distance="550" swimtime="00:07:05.93" />
                    <SPLIT distance="600" swimtime="00:07:45.54" />
                    <SPLIT distance="650" swimtime="00:08:24.64" />
                    <SPLIT distance="700" swimtime="00:09:04.50" />
                    <SPLIT distance="750" swimtime="00:09:43.76" />
                    <SPLIT distance="800" swimtime="00:10:23.59" />
                    <SPLIT distance="850" swimtime="00:11:03.20" />
                    <SPLIT distance="900" swimtime="00:11:43.13" />
                    <SPLIT distance="950" swimtime="00:12:23.51" />
                    <SPLIT distance="1000" swimtime="00:13:03.58" />
                    <SPLIT distance="1050" swimtime="00:13:43.05" />
                    <SPLIT distance="1100" swimtime="00:14:23.12" />
                    <SPLIT distance="1150" swimtime="00:15:03.14" />
                    <SPLIT distance="1200" swimtime="00:15:43.77" />
                    <SPLIT distance="1250" swimtime="00:16:24.22" />
                    <SPLIT distance="1300" swimtime="00:17:05.08" />
                    <SPLIT distance="1350" swimtime="00:17:45.17" />
                    <SPLIT distance="1400" swimtime="00:18:24.98" />
                    <SPLIT distance="1450" swimtime="00:19:04.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="372" reactiontime="+93" swimtime="00:02:30.92" resultid="16528" heatid="19417" lane="4" entrytime="00:02:34.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                    <SPLIT distance="100" swimtime="00:01:12.84" />
                    <SPLIT distance="150" swimtime="00:01:52.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="336" reactiontime="+93" swimtime="00:05:38.42" resultid="16529" heatid="19510" lane="6" entrytime="00:05:59.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.30" />
                    <SPLIT distance="100" swimtime="00:01:12.77" />
                    <SPLIT distance="150" swimtime="00:02:00.73" />
                    <SPLIT distance="200" swimtime="00:02:47.23" />
                    <SPLIT distance="250" swimtime="00:03:33.58" />
                    <SPLIT distance="300" swimtime="00:04:19.93" />
                    <SPLIT distance="350" swimtime="00:05:00.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-11-09" firstname="Elżbieta" gender="F" lastname="Nowak-Bereś" nation="POL" license="500308600162" athleteid="16530">
              <RESULTS>
                <RESULT eventid="1062" points="137" swimtime="00:00:45.02" resultid="16531" heatid="19278" lane="9" entrytime="00:00:39.99" />
                <RESULT eventid="1096" points="125" reactiontime="+100" swimtime="00:04:03.57" resultid="16532" heatid="19305" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:01.75" />
                    <SPLIT distance="100" swimtime="00:03:10.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="143" reactiontime="+107" swimtime="00:01:37.27" resultid="16533" heatid="19368" lane="7" entrytime="00:01:36.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="142" reactiontime="+97" swimtime="00:01:48.56" resultid="16534" heatid="19390" lane="6" entrytime="00:01:56.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="144" reactiontime="+98" swimtime="00:00:46.51" resultid="16535" heatid="19445" lane="3" entrytime="00:00:47.80" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="16536" heatid="19481" lane="9" entrytime="00:03:30.96" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MKPSZC" nation="POL" region="SZ" clubid="15769" name="MKP Szczecin">
          <CONTACT email="windmuhle@wp.pl" name="Kowalczyk Piotr" phone="509758055" />
          <ATHLETES>
            <ATHLETE birthdate="1935-08-21" firstname="Stefania" gender="F" lastname="Noetzel" nation="POL" athleteid="15790">
              <RESULTS>
                <RESULT eventid="1222" points="86" swimtime="00:05:04.65" resultid="15791" heatid="19355" lane="2" entrytime="00:04:59.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.29" />
                    <SPLIT distance="100" swimtime="00:03:49.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="76" swimtime="00:02:27.17" resultid="15792" heatid="19427" lane="5" entrytime="00:02:20.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="76" swimtime="00:01:07.45" resultid="15793" heatid="19539" lane="7" entrytime="00:01:06.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-12" firstname="Zbigniew" gender="M" lastname="Szozda" nation="POL" athleteid="15783">
              <RESULTS>
                <RESULT eventid="1239" points="232" reactiontime="+105" swimtime="00:03:16.00" resultid="15784" heatid="19361" lane="5" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.95" />
                    <SPLIT distance="100" swimtime="00:01:33.70" />
                    <SPLIT distance="150" swimtime="00:02:24.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="262" reactiontime="+104" swimtime="00:01:18.53" resultid="15785" heatid="19402" lane="0" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="252" reactiontime="+99" swimtime="00:01:27.95" resultid="15786" heatid="19438" lane="7" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="219" reactiontime="+82" swimtime="00:01:21.10" resultid="15787" heatid="19474" lane="6" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="180" reactiontime="+110" swimtime="00:01:25.10" resultid="15788" heatid="19519" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="265" reactiontime="+106" swimtime="00:00:39.28" resultid="15789" heatid="19551" lane="3" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-02-06" firstname="Lech" gender="M" lastname="Orecki" nation="POL" athleteid="15770">
              <RESULTS>
                <RESULT comment="O4 - Start wykonany przed sygnłem (przedwczesny start) (Time: 15:32)" eventid="1079" reactiontime="+52" status="DSQ" swimtime="00:00:30.23" resultid="15771" heatid="19291" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="14207" points="270" reactiontime="+116" swimtime="00:21:50.62" resultid="15772" heatid="19622" lane="0" entrytime="00:22:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.60" />
                    <SPLIT distance="100" swimtime="00:01:20.58" />
                    <SPLIT distance="150" swimtime="00:02:04.13" />
                    <SPLIT distance="200" swimtime="00:02:48.81" />
                    <SPLIT distance="250" swimtime="00:03:33.87" />
                    <SPLIT distance="300" swimtime="00:04:18.07" />
                    <SPLIT distance="350" swimtime="00:05:02.39" />
                    <SPLIT distance="400" swimtime="00:05:47.01" />
                    <SPLIT distance="450" swimtime="00:06:31.40" />
                    <SPLIT distance="500" swimtime="00:07:15.92" />
                    <SPLIT distance="550" swimtime="00:08:00.55" />
                    <SPLIT distance="600" swimtime="00:08:45.57" />
                    <SPLIT distance="650" swimtime="00:10:14.36" />
                    <SPLIT distance="700" swimtime="00:10:59.83" />
                    <SPLIT distance="750" swimtime="00:11:43.91" />
                    <SPLIT distance="800" swimtime="00:12:27.39" />
                    <SPLIT distance="850" swimtime="00:13:12.21" />
                    <SPLIT distance="900" swimtime="00:13:55.97" />
                    <SPLIT distance="950" swimtime="00:14:39.87" />
                    <SPLIT distance="1000" swimtime="00:15:24.01" />
                    <SPLIT distance="1050" swimtime="00:16:07.31" />
                    <SPLIT distance="1100" swimtime="00:16:50.89" />
                    <SPLIT distance="1150" swimtime="00:17:34.79" />
                    <SPLIT distance="1200" swimtime="00:18:17.59" />
                    <SPLIT distance="1250" swimtime="00:19:00.92" />
                    <SPLIT distance="1300" swimtime="00:19:45.39" />
                    <SPLIT distance="1350" swimtime="00:20:29.82" />
                    <SPLIT distance="1400" swimtime="00:21:12.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="15773" heatid="19345" lane="4" entrytime="00:00:42.00" />
                <RESULT eventid="1273" points="298" reactiontime="+89" swimtime="00:01:07.22" resultid="15774" heatid="19381" lane="9" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="15775" heatid="19472" lane="1" entrytime="00:01:50.00" />
                <RESULT eventid="1508" points="283" reactiontime="+98" swimtime="00:02:31.34" resultid="15776" heatid="19491" lane="5" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.98" />
                    <SPLIT distance="100" swimtime="00:01:12.46" />
                    <SPLIT distance="150" swimtime="00:01:52.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="171" reactiontime="+91" swimtime="00:03:10.18" resultid="15777" heatid="19533" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.64" />
                    <SPLIT distance="100" swimtime="00:01:34.27" />
                    <SPLIT distance="150" swimtime="00:02:23.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="15778" heatid="19704" lane="7" entrytime="00:05:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-10-02" firstname="Jadwiga" gender="F" lastname="Weber" nation="POL" athleteid="15779">
              <RESULTS>
                <RESULT eventid="1187" points="238" reactiontime="+83" swimtime="00:00:41.40" resultid="15780" heatid="19338" lane="7" entrytime="00:00:43.00" />
                <RESULT eventid="1457" points="227" reactiontime="+89" swimtime="00:01:30.16" resultid="15781" heatid="19467" lane="0" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="240" reactiontime="+86" swimtime="00:03:11.81" resultid="15782" heatid="19528" lane="9" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.85" />
                    <SPLIT distance="100" swimtime="00:01:32.67" />
                    <SPLIT distance="150" swimtime="00:02:22.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-08-10" firstname="Małgorzata" gender="F" lastname="Serbin" nation="POL" athleteid="15794">
              <RESULTS>
                <RESULT eventid="1147" points="387" reactiontime="+85" swimtime="00:10:57.47" resultid="15795" heatid="19596" lane="2" entrytime="00:10:51.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.88" />
                    <SPLIT distance="100" swimtime="00:01:15.13" />
                    <SPLIT distance="150" swimtime="00:01:55.60" />
                    <SPLIT distance="200" swimtime="00:02:36.46" />
                    <SPLIT distance="250" swimtime="00:03:17.49" />
                    <SPLIT distance="300" swimtime="00:03:58.55" />
                    <SPLIT distance="350" swimtime="00:04:39.83" />
                    <SPLIT distance="400" swimtime="00:05:21.53" />
                    <SPLIT distance="450" swimtime="00:06:03.40" />
                    <SPLIT distance="500" swimtime="00:06:45.34" />
                    <SPLIT distance="550" swimtime="00:07:27.15" />
                    <SPLIT distance="600" swimtime="00:08:09.06" />
                    <SPLIT distance="650" swimtime="00:08:50.96" />
                    <SPLIT distance="700" swimtime="00:09:33.48" />
                    <SPLIT distance="750" swimtime="00:10:16.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="401" reactiontime="+82" swimtime="00:01:09.03" resultid="15796" heatid="19371" lane="6" entrytime="00:01:10.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="424" reactiontime="+79" swimtime="00:02:27.44" resultid="15797" heatid="19484" lane="8" entrytime="00:02:31.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.96" />
                    <SPLIT distance="100" swimtime="00:01:11.30" />
                    <SPLIT distance="150" swimtime="00:01:49.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="292" reactiontime="+82" swimtime="00:02:59.52" resultid="15798" heatid="19528" lane="6" entrytime="00:02:59.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.12" />
                    <SPLIT distance="100" swimtime="00:01:28.26" />
                    <SPLIT distance="150" swimtime="00:02:14.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="415" reactiontime="+88" swimtime="00:05:14.36" resultid="15799" heatid="19698" lane="1" entrytime="00:05:17.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                    <SPLIT distance="100" swimtime="00:01:13.97" />
                    <SPLIT distance="150" swimtime="00:01:53.51" />
                    <SPLIT distance="200" swimtime="00:02:33.47" />
                    <SPLIT distance="250" swimtime="00:03:13.77" />
                    <SPLIT distance="300" swimtime="00:03:54.27" />
                    <SPLIT distance="350" swimtime="00:04:34.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06611" nation="POL" region="SLA" clubid="18327" name="MKP Wodnik 29 Tychy">
          <CONTACT city="Tychy" email="marekmrozw29@gmail.com" internet="www.wodnik29.pl" name="Mróz Marek" phone="782-985-239" state="SLA" street="Damrota 170" zip="43-100" />
          <ATHLETES>
            <ATHLETE birthdate="1947-05-09" firstname="Stanisław" gender="M" lastname="Zieliński" nation="POL" athleteid="18328">
              <RESULTS>
                <RESULT eventid="1079" points="130" reactiontime="+88" swimtime="00:00:39.97" resultid="18329" heatid="19287" lane="6" entrytime="00:00:36.96" />
                <RESULT eventid="14189" points="115" reactiontime="+87" swimtime="00:15:11.49" resultid="18330" heatid="19615" lane="8" entrytime="00:16:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.78" />
                    <SPLIT distance="100" swimtime="00:01:43.29" />
                    <SPLIT distance="150" swimtime="00:02:40.74" />
                    <SPLIT distance="200" swimtime="00:03:37.60" />
                    <SPLIT distance="250" swimtime="00:04:35.25" />
                    <SPLIT distance="300" swimtime="00:05:33.28" />
                    <SPLIT distance="350" swimtime="00:06:31.21" />
                    <SPLIT distance="400" swimtime="00:07:30.02" />
                    <SPLIT distance="450" swimtime="00:08:28.48" />
                    <SPLIT distance="500" swimtime="00:09:26.96" />
                    <SPLIT distance="550" swimtime="00:10:26.66" />
                    <SPLIT distance="600" swimtime="00:11:25.64" />
                    <SPLIT distance="650" swimtime="00:12:23.63" />
                    <SPLIT distance="700" swimtime="00:13:21.36" />
                    <SPLIT distance="750" swimtime="00:14:18.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="124" reactiontime="+96" swimtime="00:01:30.01" resultid="18331" heatid="19377" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="18332" heatid="19487" lane="2" entrytime="00:03:15.00" />
                <RESULT eventid="1681" points="152" reactiontime="+71" swimtime="00:00:47.22" resultid="18333" heatid="19549" lane="0" entrytime="00:00:48.71" />
                <RESULT eventid="1744" points="116" swimtime="00:07:14.98" resultid="18334" heatid="19700" lane="6" entrytime="00:07:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.24" />
                    <SPLIT distance="100" swimtime="00:01:41.76" />
                    <SPLIT distance="150" swimtime="00:02:38.11" />
                    <SPLIT distance="200" swimtime="00:03:33.84" />
                    <SPLIT distance="250" swimtime="00:04:30.48" />
                    <SPLIT distance="300" swimtime="00:05:27.37" />
                    <SPLIT distance="350" swimtime="00:06:23.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-07-13" firstname="Szymon" gender="M" lastname="Warwas" nation="POL" license="106611700009" athleteid="18335">
              <RESULTS>
                <RESULT eventid="1079" points="580" reactiontime="+66" swimtime="00:00:24.29" resultid="18336" heatid="19304" lane="7" entrytime="00:00:23.80" />
                <RESULT eventid="14189" reactiontime="+70" status="OTL" swimtime="00:10:41.03" resultid="18337" heatid="19618" lane="8" entrytime="00:09:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.85" />
                    <SPLIT distance="100" swimtime="00:01:08.05" />
                    <SPLIT distance="150" swimtime="00:01:44.69" />
                    <SPLIT distance="200" swimtime="00:02:22.48" />
                    <SPLIT distance="250" swimtime="00:03:01.84" />
                    <SPLIT distance="300" swimtime="00:03:41.71" />
                    <SPLIT distance="350" swimtime="00:04:22.31" />
                    <SPLIT distance="400" swimtime="00:05:03.21" />
                    <SPLIT distance="450" swimtime="00:05:44.87" />
                    <SPLIT distance="500" swimtime="00:06:27.26" />
                    <SPLIT distance="550" swimtime="00:07:09.37" />
                    <SPLIT distance="650" swimtime="00:09:17.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="461" swimtime="00:00:28.76" resultid="18338" heatid="19353" lane="2" entrytime="00:00:27.20" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="18339" heatid="19388" lane="6" entrytime="00:00:53.50" />
                <RESULT eventid="14243" status="DNS" swimtime="00:00:00.00" resultid="18340" heatid="19409" lane="4" entrytime="00:01:01.50" />
                <RESULT eventid="1440" points="551" reactiontime="+67" swimtime="00:00:26.59" resultid="18341" heatid="19464" lane="7" entrytime="00:00:25.80" />
                <RESULT eventid="1474" points="451" reactiontime="+72" swimtime="00:01:03.78" resultid="18342" heatid="19478" lane="4" entrytime="00:00:59.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00816" nation="POL" region="SZ" clubid="18021" name="MKS Neptun Stargard">
          <CONTACT city="Stargard" email="prezes@mksneptun.pl" internet="www.mksneptun.pl" name="Miedzyszkolny Klub Sportowy &quot;Neptun&quot;" phone="602731410" state="ZACHO" street="Os. Zachód B 15" zip="73-110" />
          <ATHLETES>
            <ATHLETE birthdate="1994-09-30" firstname="Mateusz" gender="M" lastname="Drozd" nation="POL" athleteid="18050">
              <RESULTS>
                <RESULT eventid="1079" points="572" reactiontime="+77" swimtime="00:00:24.40" resultid="18051" heatid="19304" lane="1" entrytime="00:00:23.82" />
                <RESULT eventid="1113" points="548" reactiontime="+73" swimtime="00:02:13.95" resultid="18052" heatid="19318" lane="6" entrytime="00:02:12.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.90" />
                    <SPLIT distance="100" swimtime="00:01:02.57" />
                    <SPLIT distance="150" swimtime="00:01:42.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="545" reactiontime="+70" swimtime="00:01:01.56" resultid="18053" heatid="19410" lane="7" entrytime="00:00:59.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="18054" heatid="19496" lane="3" entrytime="00:01:56.90" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="18055" heatid="19512" lane="5" entrytime="00:04:40.24" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="18056" heatid="19559" lane="8" entrytime="00:00:31.94" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-02-20" firstname="Mariusz" gender="M" lastname="Chrzan" nation="POL" athleteid="18045">
              <RESULTS>
                <RESULT eventid="1113" points="394" reactiontime="+79" swimtime="00:02:29.45" resultid="18046" heatid="19316" lane="7" entrytime="00:02:30.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.51" />
                    <SPLIT distance="100" swimtime="00:01:08.75" />
                    <SPLIT distance="150" swimtime="00:01:53.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="430" reactiontime="+83" swimtime="00:01:06.59" resultid="18047" heatid="19406" lane="2" entrytime="00:01:09.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="427" reactiontime="+79" swimtime="00:02:11.92" resultid="18048" heatid="19494" lane="2" entrytime="00:02:12.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.40" />
                    <SPLIT distance="100" swimtime="00:01:03.05" />
                    <SPLIT distance="150" swimtime="00:01:37.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="382" reactiontime="+78" swimtime="00:01:06.24" resultid="18049" heatid="19522" lane="8" entrytime="00:01:10.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-05-10" firstname="Bartosz" gender="M" lastname="Pabich" nation="POL" athleteid="18057">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="18058" heatid="19302" lane="4" entrytime="00:00:25.03" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="18059" heatid="19388" lane="3" entrytime="00:00:52.94" />
                <RESULT eventid="1341" status="DNS" swimtime="00:00:00.00" resultid="18060" heatid="19418" lane="5" entrytime="00:02:12.09" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="18061" heatid="19464" lane="6" entrytime="00:00:25.63" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="18062" heatid="19496" lane="5" entrytime="00:01:56.09" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="18063" heatid="19525" lane="3" entrytime="00:00:58.24" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02711" nation="POL" region="SLA" clubid="18593" name="MOS Dąbrowa Górnicza">
          <CONTACT name="Waliczek Mariusz" />
          <ATHLETES>
            <ATHLETE birthdate="1997-10-22" firstname="Anna" gender="F" lastname="Teresko" nation="POL" license="102711100021" athleteid="18599">
              <RESULTS>
                <RESULT eventid="1187" points="538" reactiontime="+65" swimtime="00:00:31.56" resultid="18600" heatid="19341" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1324" points="487" reactiontime="+85" swimtime="00:02:32.00" resultid="18601" heatid="19412" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                    <SPLIT distance="100" swimtime="00:01:11.17" />
                    <SPLIT distance="150" swimtime="00:01:51.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="529" reactiontime="+73" swimtime="00:01:08.02" resultid="18602" heatid="19469" lane="4" entrytime="00:01:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="601" reactiontime="+83" swimtime="00:02:11.23" resultid="18603" heatid="19484" lane="5" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                    <SPLIT distance="100" swimtime="00:01:04.43" />
                    <SPLIT distance="150" swimtime="00:01:38.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" status="DNS" swimtime="00:00:00.00" resultid="18604" heatid="19505" lane="4" entrytime="00:04:59.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-10-21" firstname="Patryk" gender="M" lastname="Droś" nation="POL" license="102711200122" athleteid="18594">
              <RESULTS>
                <RESULT eventid="1239" points="563" reactiontime="+72" swimtime="00:02:25.83" resultid="18595" heatid="19365" lane="4" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.73" />
                    <SPLIT distance="100" swimtime="00:01:08.54" />
                    <SPLIT distance="150" swimtime="00:01:46.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="603" reactiontime="+65" swimtime="00:00:53.19" resultid="18596" heatid="19388" lane="7" entrytime="00:00:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="611" reactiontime="+69" swimtime="00:01:05.51" resultid="18597" heatid="19443" lane="4" entrytime="00:01:02.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="609" reactiontime="+74" swimtime="00:01:57.20" resultid="18598" heatid="19496" lane="4" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.73" />
                    <SPLIT distance="100" swimtime="00:00:56.66" />
                    <SPLIT distance="150" swimtime="00:01:27.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-06-01" firstname="Dawid" gender="M" lastname="Nowodworski" nation="POL" license="102711200028" athleteid="18605">
              <RESULTS>
                <RESULT eventid="1205" points="569" reactiontime="+84" swimtime="00:00:26.80" resultid="18606" heatid="19352" lane="3" entrytime="00:00:28.50" />
                <RESULT eventid="14243" points="640" reactiontime="+77" swimtime="00:00:58.36" resultid="18607" heatid="19410" lane="4" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="18608" heatid="19443" lane="6" entrytime="00:01:05.00" />
                <RESULT eventid="1440" points="631" reactiontime="+69" swimtime="00:00:25.41" resultid="18609" heatid="19464" lane="8" entrytime="00:00:26.00" />
                <RESULT eventid="1474" points="548" reactiontime="+76" swimtime="00:00:59.75" resultid="18610" heatid="19478" lane="5" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-03-23" firstname="Bernard" gender="M" lastname="Filek" nation="POL" athleteid="18611">
              <RESULTS>
                <RESULT eventid="1079" points="517" reactiontime="+74" swimtime="00:00:25.23" resultid="18612" heatid="19303" lane="6" entrytime="00:00:24.50" />
                <RESULT eventid="14189" reactiontime="+82" status="OTL" swimtime="00:10:28.88" resultid="18613" heatid="19618" lane="2" entrytime="00:09:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.55" />
                    <SPLIT distance="100" swimtime="00:01:06.42" />
                    <SPLIT distance="150" swimtime="00:01:41.96" />
                    <SPLIT distance="200" swimtime="00:02:18.36" />
                    <SPLIT distance="250" swimtime="00:02:55.00" />
                    <SPLIT distance="300" swimtime="00:03:32.76" />
                    <SPLIT distance="350" swimtime="00:04:12.23" />
                    <SPLIT distance="400" swimtime="00:04:53.01" />
                    <SPLIT distance="500" swimtime="00:06:59.36" />
                    <SPLIT distance="550" swimtime="00:07:41.76" />
                    <SPLIT distance="600" swimtime="00:08:24.60" />
                    <SPLIT distance="750" swimtime="00:09:49.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="18614" heatid="19352" lane="4" entrytime="00:00:28.50" />
                <RESULT eventid="1341" points="362" reactiontime="+72" swimtime="00:02:32.21" resultid="18615" heatid="19418" lane="9" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.83" />
                    <SPLIT distance="100" swimtime="00:01:10.93" />
                    <SPLIT distance="150" swimtime="00:01:51.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="579" reactiontime="+77" swimtime="00:00:26.15" resultid="18616" heatid="19464" lane="1" entrytime="00:00:26.00" />
                <RESULT eventid="1474" points="438" reactiontime="+64" swimtime="00:01:04.41" resultid="18617" heatid="19478" lane="7" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="18618" heatid="19537" lane="3" entrytime="00:02:20.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="14355" name="MOSiR Ostrowiec Św.">
          <CONTACT name="Różalski Józef" />
          <ATHLETES>
            <ATHLETE birthdate="1945-03-28" firstname="Józef" gender="M" lastname="Różalski" nation="POL" license="501012700001" athleteid="14356">
              <RESULTS>
                <RESULT eventid="1079" points="225" reactiontime="+88" swimtime="00:00:33.28" resultid="14357" heatid="19288" lane="5" entrytime="00:00:34.80" />
                <RESULT eventid="1113" points="137" reactiontime="+89" swimtime="00:03:32.36" resultid="14358" heatid="19311" lane="8" entrytime="00:03:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.58" />
                    <SPLIT distance="100" swimtime="00:01:45.35" />
                    <SPLIT distance="150" swimtime="00:02:48.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="127" reactiontime="+91" swimtime="00:03:58.99" resultid="14359" heatid="19360" lane="7" entrytime="00:04:04.00" />
                <RESULT eventid="14243" points="160" reactiontime="+91" swimtime="00:01:32.65" resultid="14360" heatid="19399" lane="6" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="211" reactiontime="+85" swimtime="00:00:36.61" resultid="14361" heatid="19453" lane="7" entrytime="00:00:37.00" />
                <RESULT eventid="1578" points="117" reactiontime="+94" swimtime="00:08:01.39" resultid="14362" heatid="19508" lane="9" entrytime="00:08:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.61" />
                    <SPLIT distance="100" swimtime="00:01:55.44" />
                    <SPLIT distance="150" swimtime="00:02:59.82" />
                    <SPLIT distance="200" swimtime="00:04:06.43" />
                    <SPLIT distance="250" swimtime="00:05:11.54" />
                    <SPLIT distance="300" swimtime="00:06:17.28" />
                    <SPLIT distance="350" swimtime="00:07:09.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="134" reactiontime="+98" swimtime="00:01:33.79" resultid="14363" heatid="19518" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="190" reactiontime="+99" swimtime="00:00:43.91" resultid="14364" heatid="19549" lane="2" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOTYL" nation="POL" region="PDK" clubid="15053" name="MOTYL MOSiR STALOWA WOLA">
          <CONTACT city="Stalowa Wola" email="lorkowska@wp.pl" name="Jarosław Niedbałowski" phone="600831914" state="PODK" street="Hutnicza 15" zip="37-450" />
          <ATHLETES>
            <ATHLETE birthdate="1967-04-17" firstname="Maria" gender="F" lastname="Petecka" nation="POL" athleteid="15063">
              <RESULTS>
                <RESULT eventid="1062" points="269" reactiontime="+94" swimtime="00:00:35.98" resultid="15064" heatid="19279" lane="7" entrytime="00:00:36.00" />
                <RESULT eventid="1096" points="244" reactiontime="+97" swimtime="00:03:14.82" resultid="15065" heatid="19306" lane="5" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.72" />
                    <SPLIT distance="100" swimtime="00:01:33.98" />
                    <SPLIT distance="150" swimtime="00:02:28.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="255" reactiontime="+96" swimtime="00:03:32.19" resultid="15066" heatid="19356" lane="4" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.91" />
                    <SPLIT distance="100" swimtime="00:01:43.26" />
                    <SPLIT distance="150" swimtime="00:02:38.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="254" reactiontime="+96" swimtime="00:01:29.45" resultid="15067" heatid="19392" lane="7" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="245" reactiontime="+95" swimtime="00:01:39.57" resultid="15068" heatid="19429" lane="2" entrytime="00:01:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="244" reactiontime="+94" swimtime="00:00:39.00" resultid="15069" heatid="19446" lane="7" entrytime="00:00:40.00" />
                <RESULT eventid="1595" points="182" reactiontime="+101" swimtime="00:01:36.28" resultid="15070" heatid="19513" lane="5" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="251" reactiontime="+96" swimtime="00:00:45.40" resultid="15071" heatid="19541" lane="2" entrytime="00:00:46.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-14" firstname="Arkadiusz" gender="M" lastname="Berwecki" nation="POL" athleteid="15054">
              <RESULTS>
                <RESULT eventid="1079" points="444" reactiontime="+73" swimtime="00:00:26.54" resultid="15055" heatid="19293" lane="7" entrytime="00:00:29.99" />
                <RESULT eventid="1113" points="485" reactiontime="+77" swimtime="00:02:19.45" resultid="15056" heatid="19318" lane="8" entrytime="00:02:19.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.55" />
                    <SPLIT distance="100" swimtime="00:01:07.85" />
                    <SPLIT distance="150" swimtime="00:01:46.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="483" reactiontime="+82" swimtime="00:00:57.25" resultid="15057" heatid="19387" lane="2" entrytime="00:00:56.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="435" reactiontime="+90" swimtime="00:02:23.25" resultid="15058" heatid="19418" lane="1" entrytime="00:02:24.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                    <SPLIT distance="100" swimtime="00:01:09.05" />
                    <SPLIT distance="150" swimtime="00:01:46.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="473" reactiontime="+79" swimtime="00:00:27.96" resultid="15059" heatid="19462" lane="3" entrytime="00:00:27.49" />
                <RESULT eventid="1508" points="498" reactiontime="+80" swimtime="00:02:05.29" resultid="15060" heatid="19495" lane="6" entrytime="00:02:05.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.66" />
                    <SPLIT distance="100" swimtime="00:01:01.82" />
                    <SPLIT distance="150" swimtime="00:01:33.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="481" reactiontime="+76" swimtime="00:01:01.35" resultid="15061" heatid="19525" lane="8" entrytime="00:01:00.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="466" reactiontime="+89" swimtime="00:04:33.69" resultid="15062" heatid="19708" lane="1" entrytime="00:04:31.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.78" />
                    <SPLIT distance="100" swimtime="00:01:04.46" />
                    <SPLIT distance="150" swimtime="00:01:39.01" />
                    <SPLIT distance="200" swimtime="00:02:14.17" />
                    <SPLIT distance="250" swimtime="00:02:49.48" />
                    <SPLIT distance="300" swimtime="00:03:24.94" />
                    <SPLIT distance="350" swimtime="00:04:00.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="SLO" clubid="15197" name="MPK Prievidza">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1966-01-01" firstname="Petr" gender="M" lastname="Soukup" nation="SLO" athleteid="15209">
              <RESULTS>
                <RESULT eventid="1079" points="361" reactiontime="+87" swimtime="00:00:28.43" resultid="15210" heatid="19298" lane="0" entrytime="00:00:27.80" />
                <RESULT eventid="1273" points="340" reactiontime="+92" swimtime="00:01:04.33" resultid="15211" heatid="19383" lane="7" entrytime="00:01:02.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="366" reactiontime="+92" swimtime="00:02:18.85" resultid="15212" heatid="19493" lane="2" entrytime="00:02:17.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.85" />
                    <SPLIT distance="100" swimtime="00:01:07.57" />
                    <SPLIT distance="150" swimtime="00:01:43.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="291" reactiontime="+92" swimtime="00:01:12.53" resultid="15213" heatid="19521" lane="2" entrytime="00:01:12.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Nina" gender="F" lastname="Hlatká" nation="SLO" athleteid="15198">
              <RESULTS>
                <RESULT eventid="1062" points="345" reactiontime="+93" swimtime="00:00:33.13" resultid="15199" heatid="19280" lane="1" entrytime="00:00:33.80" />
                <RESULT eventid="1256" points="327" reactiontime="+90" swimtime="00:01:13.85" resultid="15200" heatid="19371" lane="9" entrytime="00:01:14.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="250" reactiontime="+89" swimtime="00:00:38.69" resultid="15201" heatid="19446" lane="2" entrytime="00:00:39.40" />
                <RESULT eventid="1664" points="251" reactiontime="+94" swimtime="00:00:45.39" resultid="15202" heatid="19541" lane="0" entrytime="00:00:47.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-01" firstname="Mária" gender="F" lastname="Hausnerová" nation="SLO" athleteid="15203">
              <RESULTS>
                <RESULT eventid="1062" points="231" reactiontime="+90" swimtime="00:00:37.85" resultid="15204" heatid="19278" lane="5" entrytime="00:00:37.90" />
                <RESULT eventid="1187" points="178" reactiontime="+82" swimtime="00:00:45.56" resultid="15205" heatid="19338" lane="9" entrytime="00:00:46.70" />
                <RESULT eventid="1256" points="209" reactiontime="+94" swimtime="00:01:25.72" resultid="15206" heatid="19368" lane="5" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="182" reactiontime="+71" swimtime="00:01:37.03" resultid="15207" heatid="19466" lane="7" entrytime="00:01:40.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="173" reactiontime="+51" swimtime="00:03:33.66" resultid="15208" heatid="19527" lane="1" entrytime="00:03:40.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.25" />
                    <SPLIT distance="100" swimtime="00:01:44.57" />
                    <SPLIT distance="150" swimtime="00:02:39.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="004/03" nation="POL" region="LBL" clubid="14287" name="MUKS Lider Chełm">
          <ATHLETES>
            <ATHLETE birthdate="1941-10-11" firstname="Janusz" gender="M" lastname="Golik" nation="POL" license="100403700118" athleteid="14288">
              <RESULTS>
                <RESULT eventid="1239" points="108" reactiontime="+128" swimtime="00:04:12.50" resultid="14289" heatid="19360" lane="1" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.88" />
                    <SPLIT distance="100" swimtime="00:02:05.89" />
                    <SPLIT distance="150" swimtime="00:03:11.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="49" reactiontime="+132" swimtime="00:04:55.58" resultid="14290" heatid="19414" lane="0" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.26" />
                    <SPLIT distance="100" swimtime="00:02:19.85" />
                    <SPLIT distance="150" swimtime="00:03:38.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="130" reactiontime="+107" swimtime="00:01:49.65" resultid="14291" heatid="19436" lane="0" entrytime="00:01:43.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="79" reactiontime="+114" swimtime="00:00:50.66" resultid="14292" heatid="19451" lane="6" entrytime="00:00:47.50" />
                <RESULT eventid="1613" points="71" reactiontime="+119" swimtime="00:01:56.01" resultid="14293" heatid="19517" lane="4" entrytime="00:01:54.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="162" reactiontime="+124" swimtime="00:00:46.31" resultid="14294" heatid="19550" lane="2" entrytime="00:00:44.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NABAIJI" nation="POL" clubid="16584" name="Nabaiji Team Decathlon">
          <CONTACT city="Warszawa" email="filip.wojciechowski@decathlon.com" name="Filip Wojciechowski" phone="731981998" street="Ostrobramska 97" zip="04-118" />
          <ATHLETES>
            <ATHLETE birthdate="1994-01-01" firstname="Paweł" gender="M" lastname="Bednarczyk" nation="POL" athleteid="16618">
              <RESULTS>
                <RESULT eventid="1079" points="592" reactiontime="+77" swimtime="00:00:24.12" resultid="16619" heatid="19304" lane="6" entrytime="00:00:23.69" entrycourse="SCM" />
                <RESULT eventid="14189" reactiontime="+80" status="OTL" swimtime="00:10:02.93" resultid="16620" heatid="19618" lane="5" entrytime="00:09:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.00" />
                    <SPLIT distance="100" swimtime="00:01:05.01" />
                    <SPLIT distance="150" swimtime="00:01:40.10" />
                    <SPLIT distance="200" swimtime="00:02:15.80" />
                    <SPLIT distance="250" swimtime="00:02:51.76" />
                    <SPLIT distance="300" swimtime="00:03:28.81" />
                    <SPLIT distance="350" swimtime="00:04:06.66" />
                    <SPLIT distance="400" swimtime="00:04:45.31" />
                    <SPLIT distance="450" swimtime="00:05:24.46" />
                    <SPLIT distance="500" swimtime="00:06:03.94" />
                    <SPLIT distance="550" swimtime="00:06:44.04" />
                    <SPLIT distance="600" swimtime="00:07:24.20" />
                    <SPLIT distance="650" swimtime="00:08:04.66" />
                    <SPLIT distance="700" swimtime="00:08:45.25" />
                    <SPLIT distance="750" swimtime="00:09:24.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="608" reactiontime="+79" swimtime="00:00:53.02" resultid="16621" heatid="19388" lane="4" entrytime="00:00:52.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="564" reactiontime="+79" swimtime="00:01:00.85" resultid="16622" heatid="19410" lane="1" entrytime="00:01:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="627" reactiontime="+73" swimtime="00:00:25.47" resultid="16623" heatid="19464" lane="5" entrytime="00:00:25.00" entrycourse="SCM" />
                <RESULT eventid="1508" points="538" reactiontime="+79" swimtime="00:02:02.11" resultid="16624" heatid="19496" lane="8" entrytime="00:02:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.19" />
                    <SPLIT distance="150" swimtime="00:01:30.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="597" reactiontime="+77" swimtime="00:00:57.07" resultid="16625" heatid="19525" lane="4" entrytime="00:00:57.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="16626" heatid="19708" lane="7" entrytime="00:04:30.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-03-31" firstname="Agnieszka" gender="F" lastname="Dusza-Sabadasz" nation="POL" athleteid="16611">
              <RESULTS>
                <RESULT eventid="1062" points="211" reactiontime="+94" swimtime="00:00:38.98" resultid="16612" heatid="19277" lane="7" entrytime="00:00:43.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-11-04" firstname="Tomasz" gender="M" lastname="Sabadasz" nation="POL" athleteid="16585">
              <RESULTS>
                <RESULT eventid="1079" points="240" reactiontime="+88" swimtime="00:00:32.59" resultid="16586" heatid="19290" lane="8" entrytime="00:00:32.96" entrycourse="SCM" />
                <RESULT eventid="1113" points="184" reactiontime="+88" swimtime="00:03:12.60" resultid="16587" heatid="19311" lane="5" entrytime="00:03:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.83" />
                    <SPLIT distance="100" swimtime="00:01:34.82" />
                    <SPLIT distance="150" swimtime="00:02:30.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="221" reactiontime="+89" swimtime="00:01:14.33" resultid="16588" heatid="19377" lane="1" entrytime="00:01:22.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="193" reactiontime="+87" swimtime="00:01:27.03" resultid="16589" heatid="19400" lane="4" entrytime="00:01:26.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="197" reactiontime="+90" swimtime="00:00:37.46" resultid="16590" heatid="19454" lane="0" entrytime="00:00:36.17" entrycourse="SCM" />
                <RESULT eventid="1508" points="184" reactiontime="+80" swimtime="00:02:54.61" resultid="16591" heatid="19489" lane="9" entrytime="00:02:57.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.12" />
                    <SPLIT distance="100" swimtime="00:01:23.81" />
                    <SPLIT distance="150" swimtime="00:02:10.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Martyna" gender="F" lastname="Górajewska" nation="POL" athleteid="16592">
              <RESULTS>
                <RESULT eventid="1062" points="372" reactiontime="+90" swimtime="00:00:32.29" resultid="16593" heatid="19282" lane="2" entrytime="00:00:30.30" entrycourse="SCM" />
                <RESULT eventid="14225" points="332" reactiontime="+83" swimtime="00:01:21.78" resultid="16594" heatid="19394" lane="7" entrytime="00:01:19.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="293" reactiontime="+84" swimtime="00:02:46.77" resultid="16595" heatid="19484" lane="9" entrytime="00:02:35.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.30" />
                    <SPLIT distance="100" swimtime="00:01:17.81" />
                    <SPLIT distance="150" swimtime="00:02:01.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="335" reactiontime="+92" swimtime="00:00:41.22" resultid="16596" heatid="19543" lane="1" entrytime="00:00:40.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-01" firstname="Maciej" gender="M" lastname="Jekiełek" nation="POL" athleteid="16629">
              <RESULTS>
                <RESULT eventid="1079" points="455" reactiontime="+87" swimtime="00:00:26.34" resultid="16630" heatid="19300" lane="5" entrytime="00:00:26.00" entrycourse="SCM" />
                <RESULT eventid="14189" reactiontime="+86" status="OTL" swimtime="00:11:04.78" resultid="16631" heatid="19618" lane="9" entrytime="00:10:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="250" swimtime="00:03:04.57" />
                    <SPLIT distance="300" swimtime="00:03:46.49" />
                    <SPLIT distance="350" swimtime="00:04:28.65" />
                    <SPLIT distance="400" swimtime="00:05:12.27" />
                    <SPLIT distance="450" swimtime="00:05:55.28" />
                    <SPLIT distance="500" swimtime="00:06:39.40" />
                    <SPLIT distance="550" swimtime="00:07:24.42" />
                    <SPLIT distance="600" swimtime="00:08:09.97" />
                    <SPLIT distance="650" swimtime="00:08:55.13" />
                    <SPLIT distance="700" swimtime="00:09:38.32" />
                    <SPLIT distance="750" swimtime="00:10:21.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="364" reactiontime="+83" swimtime="00:01:10.44" resultid="16632" heatid="19404" lane="8" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="400" reactiontime="+94" swimtime="00:02:14.78" resultid="16633" heatid="19493" lane="4" entrytime="00:02:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                    <SPLIT distance="100" swimtime="00:01:05.93" />
                    <SPLIT distance="150" swimtime="00:01:40.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="16634" heatid="19707" lane="3" entrytime="00:04:40.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-04-13" firstname="Aleksander" gender="M" lastname="Ziemiński" nation="POL" athleteid="16627">
              <RESULTS>
                <RESULT eventid="1079" points="190" reactiontime="+101" swimtime="00:00:35.19" resultid="16628" heatid="19287" lane="3" entrytime="00:00:36.02" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-08-24" firstname="Aleksandra" gender="F" lastname="Czechowicz" nation="POL" athleteid="16635">
              <RESULTS>
                <RESULT eventid="1062" status="DNS" swimtime="00:00:00.00" resultid="16636" heatid="19276" lane="2" entrytime="00:00:50.00" entrycourse="SCM" />
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="16637" heatid="19369" lane="3" entrytime="00:01:20.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-01" firstname="Rafał" gender="M" lastname="Liszewski" nation="POL" athleteid="16613">
              <RESULTS>
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="16614" heatid="19314" lane="6" entrytime="00:02:40.00" entrycourse="SCM" />
                <RESULT eventid="14243" status="DNS" swimtime="00:00:00.00" resultid="16615" heatid="19404" lane="0" entrytime="00:01:15.00" entrycourse="SCM" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="16616" heatid="19439" lane="4" entrytime="00:01:20.00" entrycourse="SCM" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="16617" heatid="19558" lane="8" entrytime="00:00:33.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Magdalena" gender="F" lastname="Sproska" nation="POL" athleteid="16606">
              <RESULTS>
                <RESULT eventid="1187" points="430" reactiontime="+86" swimtime="00:00:33.99" resultid="16607" heatid="19340" lane="5" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="14225" points="492" reactiontime="+86" swimtime="00:01:11.77" resultid="16608" heatid="19395" lane="2" entrytime="00:01:14.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="441" reactiontime="+76" swimtime="00:00:32.02" resultid="16609" heatid="19448" lane="6" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1664" points="454" reactiontime="+77" swimtime="00:00:37.24" resultid="16610" heatid="19543" lane="7" entrytime="00:00:40.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-10-02" firstname="Agnieszka" gender="F" lastname="Kos" nation="POL" athleteid="16602">
              <RESULTS>
                <RESULT eventid="1256" points="230" reactiontime="+93" swimtime="00:01:23.02" resultid="16603" heatid="19369" lane="5" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="191" reactiontime="+95" swimtime="00:03:12.19" resultid="16604" heatid="19482" lane="4" entrytime="00:02:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                    <SPLIT distance="100" swimtime="00:01:29.46" />
                    <SPLIT distance="150" swimtime="00:02:21.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="179" reactiontime="+101" swimtime="00:06:55.83" resultid="16605" heatid="19698" lane="8" entrytime="00:05:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.13" />
                    <SPLIT distance="100" swimtime="00:01:30.41" />
                    <SPLIT distance="200" swimtime="00:04:11.10" />
                    <SPLIT distance="250" swimtime="00:05:06.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-05-17" firstname="Zuzanna" gender="F" lastname="Kacalska" nation="POL" athleteid="16597">
              <RESULTS>
                <RESULT eventid="1062" points="402" reactiontime="+88" swimtime="00:00:31.48" resultid="16598" heatid="19281" lane="2" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1256" points="393" reactiontime="+90" swimtime="00:01:09.48" resultid="16599" heatid="19370" lane="1" entrytime="00:01:17.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="364" reactiontime="+85" swimtime="00:01:19.30" resultid="16600" heatid="19391" lane="6" entrytime="00:01:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="396" reactiontime="+85" swimtime="00:02:30.82" resultid="16601" heatid="19483" lane="3" entrytime="00:02:42.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                    <SPLIT distance="100" swimtime="00:01:12.13" />
                    <SPLIT distance="150" swimtime="00:01:51.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" status="DNS" swimtime="00:00:00.00" resultid="16640" heatid="19423" lane="2" entrytime="00:02:05.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16585" number="1" />
                    <RELAYPOSITION athleteid="16613" number="2" />
                    <RELAYPOSITION athleteid="16618" number="3" />
                    <RELAYPOSITION athleteid="16629" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" points="321" reactiontime="+90" swimtime="00:02:00.54" resultid="16641" heatid="19501" lane="3" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.09" />
                    <SPLIT distance="100" swimtime="00:01:03.69" />
                    <SPLIT distance="150" swimtime="00:01:36.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16627" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="16613" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="16629" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="16618" number="4" reactiontime="+62" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="99" agetotalmin="80" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1358" status="DNS" swimtime="00:00:00.00" resultid="16638" heatid="19420" lane="4" entrytime="00:02:17.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16597" number="1" />
                    <RELAYPOSITION athleteid="16592" number="2" />
                    <RELAYPOSITION athleteid="16606" number="3" />
                    <RELAYPOSITION athleteid="16602" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1525" points="380" reactiontime="+85" swimtime="00:02:10.10" resultid="16639" heatid="19498" lane="4" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.70" />
                    <SPLIT distance="100" swimtime="00:01:09.45" />
                    <SPLIT distance="150" swimtime="00:01:40.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16597" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="16602" number="2" reactiontime="+72" />
                    <RELAYPOSITION athleteid="16606" number="3" reactiontime="-1" />
                    <RELAYPOSITION athleteid="16592" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="330" reactiontime="+86" swimtime="00:02:08.15" resultid="16642" heatid="19321" lane="9" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.86" />
                    <SPLIT distance="100" swimtime="00:01:11.10" />
                    <SPLIT distance="150" swimtime="00:01:42.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16611" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="16613" number="2" reactiontime="+12" />
                    <RELAYPOSITION athleteid="16597" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="16629" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" status="DNS" swimtime="00:00:00.00" resultid="16643" heatid="19563" lane="9" entrytime="00:02:25.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16597" number="1" />
                    <RELAYPOSITION athleteid="16613" number="2" />
                    <RELAYPOSITION athleteid="16629" number="3" />
                    <RELAYPOSITION athleteid="16611" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="99" agetotalmin="80" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1130" points="383" reactiontime="+88" swimtime="00:02:01.90" resultid="16644" heatid="19322" lane="6" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                    <SPLIT distance="100" swimtime="00:01:08.78" />
                    <SPLIT distance="150" swimtime="00:01:37.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16592" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="16627" number="2" reactiontime="+45" />
                    <RELAYPOSITION athleteid="16606" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="16618" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="430" reactiontime="+74" swimtime="00:02:08.69" resultid="16645" heatid="19564" lane="6" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                    <SPLIT distance="100" swimtime="00:01:12.11" />
                    <SPLIT distance="150" swimtime="00:01:37.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16606" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="16592" number="2" reactiontime="+27" />
                    <RELAYPOSITION athleteid="16618" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="16627" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="CZE" clubid="18488" name="Neptun Masters Praha">
          <ATHLETES>
            <ATHLETE birthdate="1992-09-22" firstname="Denis" gender="M" lastname="Bushkov" nation="CZE" athleteid="18497">
              <RESULTS>
                <RESULT eventid="1113" points="415" reactiontime="+81" swimtime="00:02:26.93" resultid="18498" heatid="19313" lane="5" entrytime="00:02:45.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.65" />
                    <SPLIT distance="100" swimtime="00:01:08.55" />
                    <SPLIT distance="150" swimtime="00:01:51.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14189" points="476" reactiontime="+88" swimtime="00:09:27.77" resultid="18499" heatid="19618" lane="1" entrytime="00:09:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.47" />
                    <SPLIT distance="100" swimtime="00:01:06.02" />
                    <SPLIT distance="150" swimtime="00:01:41.07" />
                    <SPLIT distance="200" swimtime="00:02:16.65" />
                    <SPLIT distance="250" swimtime="00:02:52.53" />
                    <SPLIT distance="300" swimtime="00:03:28.75" />
                    <SPLIT distance="350" swimtime="00:04:05.23" />
                    <SPLIT distance="400" swimtime="00:04:41.16" />
                    <SPLIT distance="450" swimtime="00:05:17.13" />
                    <SPLIT distance="500" swimtime="00:05:53.20" />
                    <SPLIT distance="550" swimtime="00:06:29.07" />
                    <SPLIT distance="600" swimtime="00:07:05.50" />
                    <SPLIT distance="650" swimtime="00:07:41.61" />
                    <SPLIT distance="700" swimtime="00:08:17.97" />
                    <SPLIT distance="750" swimtime="00:08:54.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="342" reactiontime="+90" swimtime="00:02:35.23" resultid="18501" heatid="19417" lane="1" entrytime="00:02:45.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                    <SPLIT distance="100" swimtime="00:01:15.10" />
                    <SPLIT distance="150" swimtime="00:01:56.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="467" reactiontime="+85" swimtime="00:02:08.06" resultid="18502" heatid="19494" lane="3" entrytime="00:02:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.44" />
                    <SPLIT distance="100" swimtime="00:01:01.89" />
                    <SPLIT distance="150" swimtime="00:01:35.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="415" reactiontime="+85" swimtime="00:05:15.63" resultid="18503" heatid="19510" lane="4" entrytime="00:05:50.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                    <SPLIT distance="100" swimtime="00:01:12.70" />
                    <SPLIT distance="150" swimtime="00:01:53.81" />
                    <SPLIT distance="200" swimtime="00:02:34.55" />
                    <SPLIT distance="250" swimtime="00:03:19.51" />
                    <SPLIT distance="300" swimtime="00:04:05.33" />
                    <SPLIT distance="350" swimtime="00:04:41.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="355" swimtime="00:01:07.89" resultid="18504" heatid="19523" lane="0" entrytime="00:01:08.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="464" reactiontime="+82" swimtime="00:04:34.09" resultid="18505" heatid="19707" lane="7" entrytime="00:04:45.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                    <SPLIT distance="100" swimtime="00:01:05.25" />
                    <SPLIT distance="150" swimtime="00:01:39.30" />
                    <SPLIT distance="200" swimtime="00:02:13.80" />
                    <SPLIT distance="250" swimtime="00:02:48.73" />
                    <SPLIT distance="300" swimtime="00:03:24.08" />
                    <SPLIT distance="350" swimtime="00:03:59.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="410" swimtime="00:01:07.66" resultid="18518" heatid="19406" lane="0" entrytime="00:01:10.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-05-16" firstname="Hana" gender="F" lastname="Bohuslávková " nation="CZE" athleteid="18513">
              <RESULTS>
                <RESULT eventid="1096" points="412" reactiontime="+74" swimtime="00:02:43.66" resultid="18514" heatid="19309" lane="9" entrytime="00:02:43.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                    <SPLIT distance="100" swimtime="00:01:16.44" />
                    <SPLIT distance="150" swimtime="00:02:02.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="466" reactiontime="+85" swimtime="00:02:53.52" resultid="18515" heatid="19358" lane="5" entrytime="00:02:55.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                    <SPLIT distance="100" swimtime="00:01:23.18" />
                    <SPLIT distance="150" swimtime="00:02:07.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="472" reactiontime="+80" swimtime="00:01:20.08" resultid="18516" heatid="19432" lane="5" entrytime="00:01:17.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="440" reactiontime="+77" swimtime="00:00:37.63" resultid="18517" heatid="19545" lane="8" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-03-04" firstname="Tomáš" gender="M" lastname="Vonšovský " nation="CZE" athleteid="18506">
              <RESULTS>
                <RESULT eventid="1079" points="385" reactiontime="+79" swimtime="00:00:27.83" resultid="18507" heatid="19298" lane="2" entrytime="00:00:27.51" />
                <RESULT eventid="1205" points="346" reactiontime="+68" swimtime="00:00:31.65" resultid="18508" heatid="19350" lane="5" entrytime="00:00:31.20" />
                <RESULT eventid="14243" points="361" reactiontime="+77" swimtime="00:01:10.59" resultid="18509" heatid="19407" lane="1" entrytime="00:01:08.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="385" reactiontime="+72" swimtime="00:00:29.95" resultid="18510" heatid="19460" lane="8" entrytime="00:00:29.73" />
                <RESULT eventid="1613" points="370" reactiontime="+82" swimtime="00:01:06.97" resultid="18511" heatid="19523" lane="6" entrytime="00:01:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="362" reactiontime="+72" swimtime="00:00:35.42" resultid="18512" heatid="19554" lane="5" entrytime="00:00:36.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-08" firstname="Tomáš" gender="M" lastname="Mudruňka " nation="CZE" athleteid="18490">
              <RESULTS>
                <RESULT eventid="1079" points="379" reactiontime="+80" swimtime="00:00:27.98" resultid="18491" heatid="19296" lane="1" entrytime="00:00:28.90" />
                <RESULT eventid="1239" points="482" reactiontime="+73" swimtime="00:02:33.61" resultid="18492" heatid="19364" lane="5" entrytime="00:02:40.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="100" swimtime="00:01:13.30" />
                    <SPLIT distance="150" swimtime="00:01:53.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="342" reactiontime="+73" swimtime="00:01:11.90" resultid="18493" heatid="19407" lane="6" entrytime="00:01:08.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="538" reactiontime="+74" swimtime="00:01:08.37" resultid="18494" heatid="19442" lane="1" entrytime="00:01:10.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="18495" heatid="19458" lane="0" entrytime="00:00:31.10" />
                <RESULT eventid="1681" points="559" reactiontime="+65" swimtime="00:00:30.65" resultid="18496" heatid="19559" lane="6" entrytime="00:00:31.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NTT" nation="POL" region="MAL" clubid="15440" name="Neptun Team Tarnow">
          <CONTACT city="Tarnow" email="neptunteam.pl" internet="neptunteamtw@gmail.com" name="Dymiter" phone="792436359" state="MALOP" street="Parkowa" zip="33-100" />
          <ATHLETES>
            <ATHLETE birthdate="1986-06-23" firstname="Mateusz" gender="M" lastname="Dymiter" nation="POL" athleteid="15441">
              <RESULTS>
                <RESULT eventid="1079" points="388" reactiontime="+87" swimtime="00:00:27.76" resultid="15442" heatid="19294" lane="5" entrytime="00:00:29.00" entrycourse="SCM" />
                <RESULT eventid="1113" points="388" reactiontime="+104" swimtime="00:02:30.20" resultid="15443" heatid="19318" lane="5" entrytime="00:01:19.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.69" />
                    <SPLIT distance="100" swimtime="00:01:10.88" />
                    <SPLIT distance="150" swimtime="00:01:53.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="368" reactiontime="+92" swimtime="00:02:48.01" resultid="15444" heatid="19365" lane="3" entrytime="00:02:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                    <SPLIT distance="100" swimtime="00:01:18.67" />
                    <SPLIT distance="150" swimtime="00:02:02.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="383" reactiontime="+87" swimtime="00:01:09.26" resultid="15445" heatid="19405" lane="8" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="15446" heatid="19458" lane="8" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1578" points="363" reactiontime="+92" swimtime="00:05:30.05" resultid="15447" heatid="19511" lane="1" entrytime="00:05:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                    <SPLIT distance="100" swimtime="00:01:08.64" />
                    <SPLIT distance="150" swimtime="00:01:53.55" />
                    <SPLIT distance="200" swimtime="00:02:38.14" />
                    <SPLIT distance="250" swimtime="00:03:24.85" />
                    <SPLIT distance="300" swimtime="00:04:10.77" />
                    <SPLIT distance="350" swimtime="00:04:51.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="15448" heatid="19522" lane="9" entrytime="00:01:11.00" entrycourse="SCM" />
                <RESULT eventid="1744" points="363" reactiontime="+89" swimtime="00:04:57.45" resultid="15449" heatid="19707" lane="6" entrytime="00:04:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                    <SPLIT distance="100" swimtime="00:01:07.68" />
                    <SPLIT distance="150" swimtime="00:01:45.30" />
                    <SPLIT distance="200" swimtime="00:02:24.96" />
                    <SPLIT distance="250" swimtime="00:03:03.03" />
                    <SPLIT distance="300" swimtime="00:03:41.66" />
                    <SPLIT distance="350" swimtime="00:04:21.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-11-23" firstname="Dawid" gender="M" lastname="Wiklański" nation="POL" athleteid="15455">
              <RESULTS>
                <RESULT eventid="1079" points="177" reactiontime="+113" swimtime="00:00:36.05" resultid="15456" heatid="19288" lane="6" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1273" points="125" reactiontime="+113" swimtime="00:01:29.65" resultid="15457" heatid="19375" lane="1" entrytime="00:01:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="148" reactiontime="+119" swimtime="00:01:45.01" resultid="15458" heatid="19434" lane="2" entrytime="00:02:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="167" reactiontime="+94" swimtime="00:00:45.82" resultid="15459" heatid="19548" lane="4" entrytime="00:00:50.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-11-16" firstname="Filip" gender="M" lastname="Gawłowski" nation="POL" athleteid="15450">
              <RESULTS>
                <RESULT eventid="1079" points="169" reactiontime="+97" swimtime="00:00:36.63" resultid="15451" heatid="19286" lane="0" entrytime="00:00:40.00" entrycourse="SCM" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="15452" heatid="19375" lane="6" entrytime="00:01:35.00" entrycourse="SCM" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="15453" heatid="19434" lane="6" entrytime="00:02:05.00" entrycourse="SCM" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="15454" heatid="19548" lane="3" entrytime="00:00:52.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="14261" name="Niezrzeszeni">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1961-01-18" firstname="Wojciech" gender="M" lastname="Warchoł" nation="POL" athleteid="14921">
              <RESULTS>
                <RESULT eventid="1079" points="382" reactiontime="+83" swimtime="00:00:27.92" resultid="14922" heatid="19295" lane="9" entrytime="00:00:29.00" />
                <RESULT eventid="1273" points="368" reactiontime="+85" swimtime="00:01:02.69" resultid="14923" heatid="19381" lane="6" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="361" reactiontime="+86" swimtime="00:01:10.60" resultid="14924" heatid="19402" lane="4" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-04-04" firstname="Karolina" gender="F" lastname="Szkudlarek" nation="POL" athleteid="14610">
              <RESULTS>
                <RESULT eventid="1062" points="442" reactiontime="+85" swimtime="00:00:30.50" resultid="14611" heatid="19282" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1187" points="364" reactiontime="+83" swimtime="00:00:35.95" resultid="14612" heatid="19340" lane="1" entrytime="00:00:36.00" />
                <RESULT eventid="1256" points="423" reactiontime="+86" swimtime="00:01:07.79" resultid="14613" heatid="19371" lane="5" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="307" reactiontime="+89" swimtime="00:00:36.12" resultid="14614" heatid="19448" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="1457" points="373" reactiontime="+77" swimtime="00:01:16.42" resultid="14615" heatid="19467" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-07-15" firstname="Alina" gender="F" lastname="Piekarska " nation="POL" athleteid="14663">
              <RESULTS>
                <RESULT comment="K14 - Praca nóg w płaszczyźnie pionowej w dół (z wyjątkiem jednego ruchu po starcie i nawrocie) (Time: 10:42), K-15" eventid="1664" status="DSQ" swimtime="00:02:28.45" resultid="14664" heatid="19539" lane="9" entrytime="00:02:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-06-06" firstname="Jolanta" gender="F" lastname="Lipińska" nation="POL" athleteid="15025">
              <RESULTS>
                <RESULT eventid="1222" points="43" reactiontime="+110" swimtime="00:06:23.20" resultid="15026" heatid="19355" lane="1" entrytime="00:06:05.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:27.34" />
                    <SPLIT distance="100" swimtime="00:03:06.00" />
                    <SPLIT distance="150" swimtime="00:04:47.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="25" reactiontime="+107" swimtime="00:03:13.04" resultid="15027" heatid="19389" lane="4" entrytime="00:03:11.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:35.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="36" reactiontime="+120" swimtime="00:03:08.62" resultid="15028" heatid="19427" lane="2" entrytime="00:02:53.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="21" reactiontime="+131" swimtime="00:06:35.98" resultid="15029" heatid="19479" lane="5" entrytime="00:06:10.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:31.68" />
                    <SPLIT distance="100" swimtime="00:03:14.46" />
                    <SPLIT distance="150" swimtime="00:04:56.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="30" reactiontime="+81" swimtime="00:06:21.67" resultid="15030" heatid="19526" lane="7" entrytime="00:06:19.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:31.81" />
                    <SPLIT distance="100" swimtime="00:03:09.23" />
                    <SPLIT distance="150" swimtime="00:04:46.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="43" reactiontime="+115" swimtime="00:01:21.19" resultid="15031" heatid="19539" lane="0" entrytime="00:01:19.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-07-22" firstname="Ireneusz" gender="M" lastname="Stachurski" nation="POL" athleteid="14283">
              <RESULTS>
                <RESULT eventid="1079" points="183" reactiontime="+101" swimtime="00:00:35.63" resultid="14284" heatid="19288" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="1508" points="184" reactiontime="+113" swimtime="00:02:54.46" resultid="14285" heatid="19488" lane="5" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.57" />
                    <SPLIT distance="100" swimtime="00:01:22.47" />
                    <SPLIT distance="150" swimtime="00:02:09.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="167" reactiontime="+123" swimtime="00:06:25.27" resultid="14286" heatid="19701" lane="1" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.22" />
                    <SPLIT distance="100" swimtime="00:01:26.28" />
                    <SPLIT distance="150" swimtime="00:02:15.90" />
                    <SPLIT distance="200" swimtime="00:03:06.18" />
                    <SPLIT distance="250" swimtime="00:03:57.43" />
                    <SPLIT distance="300" swimtime="00:04:48.72" />
                    <SPLIT distance="350" swimtime="00:05:37.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-11-29" firstname="Edward" gender="M" lastname="Dziekoński" nation="POL" athleteid="17282">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="17283" heatid="19285" lane="5" entrytime="00:00:42.00" />
                <RESULT eventid="14189" status="DNS" swimtime="00:00:00.00" resultid="17284" heatid="19615" lane="7" entrytime="00:15:02.00" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="17285" heatid="19344" lane="2" entrytime="00:00:51.00" />
                <RESULT eventid="14243" status="DNS" swimtime="00:00:00.00" resultid="17286" heatid="19398" lane="4" entrytime="00:01:49.00" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="17287" heatid="19452" lane="8" entrytime="00:00:44.00" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="17288" heatid="19487" lane="1" entrytime="00:03:29.50" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="17289" heatid="19517" lane="3" entrytime="00:01:58.00" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="17290" heatid="19700" lane="7" entrytime="00:07:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1941-11-21" firstname="Zbigniew" gender="M" lastname="Dymecki" nation="POL" athleteid="14925">
              <RESULTS>
                <RESULT eventid="1113" reactiontime="+106" status="DNF" swimtime="00:00:00.00" resultid="14926" heatid="19310" lane="8" entrytime="00:04:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.65" />
                    <SPLIT distance="100" swimtime="00:02:15.08" />
                    <SPLIT distance="150" swimtime="00:03:17.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14189" status="DNS" swimtime="00:00:00.00" resultid="14927" heatid="19614" lane="3" entrytime="00:18:59.00" />
                <RESULT eventid="1239" points="73" reactiontime="+110" swimtime="00:04:48.08" resultid="14928" heatid="19360" lane="9" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.31" />
                    <SPLIT distance="100" swimtime="00:02:16.19" />
                    <SPLIT distance="150" swimtime="00:03:32.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="69" reactiontime="+111" swimtime="00:02:02.31" resultid="14929" heatid="19398" lane="0" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.21" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K10 - Dłonie przeniesione poza linię bioder (z wyjątkiem pierwszego ruchu ramon po starcie i nawrotach (Time: 16:39)" eventid="1406" reactiontime="+111" status="DSQ" swimtime="00:02:11.77" resultid="14930" heatid="19434" lane="7" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="71" reactiontime="+135" swimtime="00:03:58.94" resultid="14931" heatid="19486" lane="3" entrytime="00:04:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.05" />
                    <SPLIT distance="100" swimtime="00:01:50.73" />
                    <SPLIT distance="150" swimtime="00:02:54.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="44" reactiontime="+132" swimtime="00:04:58.34" resultid="14932" heatid="19531" lane="2" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.99" />
                    <SPLIT distance="100" swimtime="00:02:27.81" />
                    <SPLIT distance="150" swimtime="00:03:43.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="71" reactiontime="+120" swimtime="00:08:31.91" resultid="14933" heatid="19699" lane="3" entrytime="00:08:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.21" />
                    <SPLIT distance="100" swimtime="00:01:57.94" />
                    <SPLIT distance="150" swimtime="00:03:03.99" />
                    <SPLIT distance="200" swimtime="00:04:10.25" />
                    <SPLIT distance="250" swimtime="00:05:20.07" />
                    <SPLIT distance="300" swimtime="00:06:24.32" />
                    <SPLIT distance="350" swimtime="00:07:29.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-11-19" firstname="Judyta" gender="F" lastname="Sołtyk" nation="POL" athleteid="14280">
              <RESULTS>
                <RESULT eventid="1062" points="377" reactiontime="+91" swimtime="00:00:32.16" resultid="14281" heatid="19281" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1096" points="379" reactiontime="+92" swimtime="00:02:48.32" resultid="14282" heatid="19308" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                    <SPLIT distance="100" swimtime="00:01:18.52" />
                    <SPLIT distance="150" swimtime="00:02:08.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-03-06" firstname="Andrzej" gender="M" lastname="Pawlak" nation="POL" athleteid="16699">
              <RESULTS>
                <RESULT eventid="1079" points="203" reactiontime="+102" swimtime="00:00:34.46" resultid="16700" heatid="19289" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1205" points="143" reactiontime="+80" swimtime="00:00:42.40" resultid="16701" heatid="19347" lane="0" entrytime="00:00:39.00" />
                <RESULT eventid="14243" status="DNS" swimtime="00:00:00.00" resultid="16702" heatid="19400" lane="0" entrytime="00:01:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-07-23" firstname="Jakub" gender="M" lastname="Jeznach" nation="POL" athleteid="16141">
              <RESULTS>
                <RESULT eventid="14243" points="85" reactiontime="+85" swimtime="00:01:54.36" resultid="16142" heatid="19399" lane="7" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="79" reactiontime="+93" swimtime="00:00:50.63" resultid="16143" heatid="19451" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="1681" points="124" reactiontime="+79" swimtime="00:00:50.52" resultid="16144" heatid="19550" lane="9" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-12-20" firstname="Arkadiusz" gender="M" lastname="Aptewicz" nation="POL" athleteid="16212">
              <RESULTS>
                <RESULT eventid="1113" points="579" reactiontime="+76" swimtime="00:02:11.46" resultid="16213" heatid="19318" lane="2" entrytime="00:02:14.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.35" />
                    <SPLIT distance="100" swimtime="00:01:03.39" />
                    <SPLIT distance="150" swimtime="00:01:40.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="615" reactiontime="+77" swimtime="00:02:21.59" resultid="16214" heatid="19365" lane="5" entrytime="00:02:21.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                    <SPLIT distance="100" swimtime="00:01:07.60" />
                    <SPLIT distance="150" swimtime="00:01:44.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="589" reactiontime="+80" swimtime="00:01:06.31" resultid="16215" heatid="19443" lane="3" entrytime="00:01:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="591" reactiontime="+80" swimtime="00:04:40.60" resultid="16216" heatid="19512" lane="3" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.96" />
                    <SPLIT distance="100" swimtime="00:01:04.92" />
                    <SPLIT distance="150" swimtime="00:01:43.81" />
                    <SPLIT distance="200" swimtime="00:02:21.72" />
                    <SPLIT distance="250" swimtime="00:02:59.00" />
                    <SPLIT distance="300" swimtime="00:03:37.14" />
                    <SPLIT distance="350" swimtime="00:04:09.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="569" reactiontime="+67" swimtime="00:00:30.47" resultid="16217" heatid="19560" lane="7" entrytime="00:00:30.50" />
                <RESULT eventid="1744" points="615" reactiontime="+79" swimtime="00:04:09.52" resultid="16218" heatid="19708" lane="4" entrytime="00:04:17.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.36" />
                    <SPLIT distance="100" swimtime="00:00:59.48" />
                    <SPLIT distance="150" swimtime="00:01:31.12" />
                    <SPLIT distance="200" swimtime="00:02:03.00" />
                    <SPLIT distance="250" swimtime="00:02:34.68" />
                    <SPLIT distance="300" swimtime="00:03:06.77" />
                    <SPLIT distance="350" swimtime="00:03:38.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-07-11" firstname="Paweł" gender="M" lastname="Adamowicz" nation="POL" athleteid="14617">
              <RESULTS>
                <RESULT eventid="1079" reactiontime="+100" status="DNS" swimtime="00:00:00.00" resultid="14618" heatid="19286" lane="2" entrytime="00:00:39.39" />
                <RESULT eventid="14243" status="DNS" swimtime="00:00:00.00" resultid="14619" heatid="19397" lane="2" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="14620" heatid="19436" lane="8" entrytime="00:01:42.42" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="14621" heatid="19550" lane="7" entrytime="00:00:44.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-11-28" firstname="Przemysław" gender="M" lastname="Szczypiński" nation="POL" athleteid="18346">
              <RESULTS>
                <RESULT eventid="1113" points="303" reactiontime="+70" swimtime="00:02:43.20" resultid="18347" heatid="19315" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                    <SPLIT distance="100" swimtime="00:01:13.33" />
                    <SPLIT distance="150" swimtime="00:02:03.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="320" reactiontime="+69" swimtime="00:01:13.52" resultid="18348" heatid="19403" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="353" reactiontime="+67" swimtime="00:00:30.84" resultid="18349" heatid="19461" lane="9" entrytime="00:00:29.00" />
                <RESULT eventid="1578" points="291" reactiontime="+73" swimtime="00:05:55.14" resultid="18350" heatid="19510" lane="7" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.63" />
                    <SPLIT distance="100" swimtime="00:01:18.98" />
                    <SPLIT distance="150" swimtime="00:02:54.78" />
                    <SPLIT distance="200" swimtime="00:03:44.76" />
                    <SPLIT distance="250" swimtime="00:04:35.28" />
                    <SPLIT distance="300" swimtime="00:05:17.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-05-13" firstname="Maciej" gender="M" lastname="Dąbrowski" nation="POL" athleteid="16136">
              <RESULTS>
                <RESULT eventid="1205" points="238" reactiontime="+75" swimtime="00:00:35.83" resultid="16137" heatid="19348" lane="6" entrytime="00:00:35.90" />
                <RESULT eventid="14243" status="DNS" swimtime="00:00:00.00" resultid="16138" heatid="19403" lane="9" entrytime="00:01:17.70" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="16139" heatid="19455" lane="0" entrytime="00:00:34.70" />
                <RESULT eventid="1474" points="230" reactiontime="+81" swimtime="00:01:19.73" resultid="16140" heatid="19475" lane="7" entrytime="00:01:16.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-09-08" firstname="Igor" gender="M" lastname="Zalewski" nation="POL" athleteid="16265">
              <RESULTS>
                <RESULT eventid="1113" points="410" reactiontime="+76" swimtime="00:02:27.55" resultid="16266" heatid="19316" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.19" />
                    <SPLIT distance="100" swimtime="00:01:10.08" />
                    <SPLIT distance="150" swimtime="00:01:54.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14207" points="396" reactiontime="+80" swimtime="00:19:14.22" resultid="16267" heatid="19623" lane="6" entrytime="00:19:27.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                    <SPLIT distance="100" swimtime="00:01:08.86" />
                    <SPLIT distance="150" swimtime="00:01:46.62" />
                    <SPLIT distance="200" swimtime="00:02:24.40" />
                    <SPLIT distance="250" swimtime="00:03:02.65" />
                    <SPLIT distance="300" swimtime="00:03:41.07" />
                    <SPLIT distance="350" swimtime="00:04:19.91" />
                    <SPLIT distance="400" swimtime="00:04:58.78" />
                    <SPLIT distance="450" swimtime="00:05:38.33" />
                    <SPLIT distance="500" swimtime="00:06:17.66" />
                    <SPLIT distance="550" swimtime="00:06:56.79" />
                    <SPLIT distance="600" swimtime="00:07:36.19" />
                    <SPLIT distance="650" swimtime="00:08:15.48" />
                    <SPLIT distance="700" swimtime="00:08:54.81" />
                    <SPLIT distance="750" swimtime="00:09:34.08" />
                    <SPLIT distance="800" swimtime="00:10:13.37" />
                    <SPLIT distance="850" swimtime="00:10:52.41" />
                    <SPLIT distance="900" swimtime="00:11:31.22" />
                    <SPLIT distance="950" swimtime="00:12:10.01" />
                    <SPLIT distance="1000" swimtime="00:12:48.43" />
                    <SPLIT distance="1050" swimtime="00:13:27.19" />
                    <SPLIT distance="1100" swimtime="00:14:05.95" />
                    <SPLIT distance="1150" swimtime="00:14:45.02" />
                    <SPLIT distance="1200" swimtime="00:15:24.04" />
                    <SPLIT distance="1250" swimtime="00:16:02.89" />
                    <SPLIT distance="1300" swimtime="00:16:41.79" />
                    <SPLIT distance="1350" swimtime="00:17:20.18" />
                    <SPLIT distance="1400" swimtime="00:17:59.08" />
                    <SPLIT distance="1450" swimtime="00:18:37.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="454" reactiontime="+79" swimtime="00:00:58.47" resultid="16268" heatid="19383" lane="3" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="436" reactiontime="+77" swimtime="00:01:06.29" resultid="16269" heatid="19407" lane="4" entrytime="00:01:07.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="434" reactiontime="+74" swimtime="00:02:11.16" resultid="16270" heatid="19494" lane="7" entrytime="00:02:12.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.24" />
                    <SPLIT distance="100" swimtime="00:01:02.31" />
                    <SPLIT distance="150" swimtime="00:01:36.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="398" reactiontime="+75" swimtime="00:05:20.00" resultid="16271" heatid="19512" lane="8" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                    <SPLIT distance="100" swimtime="00:01:11.31" />
                    <SPLIT distance="150" swimtime="00:01:53.86" />
                    <SPLIT distance="200" swimtime="00:02:34.59" />
                    <SPLIT distance="250" swimtime="00:03:22.58" />
                    <SPLIT distance="300" swimtime="00:04:08.49" />
                    <SPLIT distance="350" swimtime="00:04:45.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="410" reactiontime="+72" swimtime="00:01:04.67" resultid="16272" heatid="19524" lane="1" entrytime="00:01:03.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="16273" heatid="19707" lane="9" entrytime="00:04:51.44" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-07-31" firstname="Piotr" gender="M" lastname="Krogulec" nation="POL" athleteid="17291">
              <RESULTS>
                <RESULT eventid="1079" points="431" reactiontime="+72" swimtime="00:00:26.81" resultid="17292" heatid="19294" lane="0" entrytime="00:00:29.50" />
                <RESULT eventid="1113" points="398" reactiontime="+89" swimtime="00:02:29.02" resultid="17293" heatid="19314" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.58" />
                    <SPLIT distance="100" swimtime="00:01:06.92" />
                    <SPLIT distance="150" swimtime="00:01:51.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="17294" heatid="19350" lane="0" entrytime="00:00:33.00" />
                <RESULT eventid="14243" status="DNS" swimtime="00:00:00.00" resultid="17295" heatid="19405" lane="0" entrytime="00:01:13.00" />
                <RESULT eventid="1440" points="425" reactiontime="+74" swimtime="00:00:28.98" resultid="17296" heatid="19457" lane="0" entrytime="00:00:32.00" />
                <RESULT eventid="1474" points="401" reactiontime="+75" swimtime="00:01:06.32" resultid="17297" heatid="19475" lane="3" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="379" reactiontime="+72" swimtime="00:02:25.96" resultid="17298" heatid="19535" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                    <SPLIT distance="100" swimtime="00:01:10.28" />
                    <SPLIT distance="150" swimtime="00:01:48.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="17299" heatid="19705" lane="0" entrytime="00:05:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-09-23" firstname="Paweł" gender="M" lastname="Wrona" nation="POL" athleteid="18543">
              <RESULTS>
                <RESULT eventid="1647" points="425" reactiontime="+64" swimtime="00:02:20.41" resultid="18544" heatid="19537" lane="6" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.98" />
                    <SPLIT distance="100" swimtime="00:01:05.54" />
                    <SPLIT distance="150" swimtime="00:01:42.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-02-01" firstname="Jolanta" gender="F" lastname="Zawadzka" nation="POL" athleteid="14622">
              <RESULTS>
                <RESULT eventid="1096" points="207" reactiontime="+97" swimtime="00:03:25.87" resultid="14623" heatid="19306" lane="7" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.46" />
                    <SPLIT distance="100" swimtime="00:01:38.08" />
                    <SPLIT distance="150" swimtime="00:02:35.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="239" reactiontime="+86" swimtime="00:01:31.20" resultid="14624" heatid="19392" lane="9" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="246" reactiontime="+97" swimtime="00:01:39.42" resultid="14625" heatid="19429" lane="0" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="233" reactiontime="+93" swimtime="00:00:39.62" resultid="14626" heatid="19446" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1664" points="283" reactiontime="+93" swimtime="00:00:43.59" resultid="14627" heatid="19541" lane="4" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-07-22" firstname="Magdalena" gender="F" lastname="Antonijczuk- Krzyśków" nation="POL" athleteid="16998">
              <RESULTS>
                <RESULT eventid="1062" status="DNS" swimtime="00:00:00.00" resultid="16999" heatid="19278" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1187" points="258" reactiontime="+66" swimtime="00:00:40.31" resultid="17000" heatid="19339" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1457" status="DNS" swimtime="00:00:00.00" resultid="17001" heatid="19466" lane="5" entrytime="00:01:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-05-22" firstname="Piotr" gender="M" lastname="Krzyśków" nation="POL" athleteid="17002">
              <RESULTS>
                <RESULT eventid="1079" points="502" reactiontime="+77" swimtime="00:00:25.48" resultid="17003" heatid="19300" lane="7" entrytime="00:00:26.30" />
                <RESULT eventid="1273" points="468" reactiontime="+77" swimtime="00:00:57.88" resultid="17004" heatid="19384" lane="4" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="17005" heatid="19462" lane="9" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-05-24" firstname="Ryszadard" gender="M" lastname="Łukowski" nation="POL" athleteid="16093">
              <RESULTS>
                <RESULT eventid="1341" points="102" reactiontime="+95" swimtime="00:03:51.93" resultid="16094" heatid="19415" lane="9" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.20" />
                    <SPLIT distance="100" swimtime="00:01:48.61" />
                    <SPLIT distance="150" swimtime="00:02:50.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="182" reactiontime="+93" swimtime="00:00:38.41" resultid="16095" heatid="19452" lane="9" entrytime="00:00:45.00" />
                <RESULT eventid="1613" points="114" reactiontime="+104" swimtime="00:01:38.99" resultid="16096" heatid="19518" lane="1" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-04-24" firstname="Igor" gender="M" lastname="Okarmus" nation="POL" athleteid="14365">
              <RESULTS>
                <RESULT eventid="14207" points="319" reactiontime="+120" swimtime="00:20:40.23" resultid="14366" heatid="19623" lane="1" entrytime="00:20:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                    <SPLIT distance="100" swimtime="00:01:12.27" />
                    <SPLIT distance="150" swimtime="00:01:51.52" />
                    <SPLIT distance="200" swimtime="00:02:31.06" />
                    <SPLIT distance="250" swimtime="00:03:10.88" />
                    <SPLIT distance="300" swimtime="00:03:50.66" />
                    <SPLIT distance="350" swimtime="00:04:30.89" />
                    <SPLIT distance="400" swimtime="00:05:10.72" />
                    <SPLIT distance="450" swimtime="00:05:52.52" />
                    <SPLIT distance="500" swimtime="00:06:33.65" />
                    <SPLIT distance="550" swimtime="00:07:14.75" />
                    <SPLIT distance="600" swimtime="00:07:56.91" />
                    <SPLIT distance="650" swimtime="00:08:38.92" />
                    <SPLIT distance="700" swimtime="00:09:21.73" />
                    <SPLIT distance="750" swimtime="00:10:04.31" />
                    <SPLIT distance="800" swimtime="00:10:46.80" />
                    <SPLIT distance="850" swimtime="00:11:29.10" />
                    <SPLIT distance="900" swimtime="00:12:11.81" />
                    <SPLIT distance="950" swimtime="00:12:54.50" />
                    <SPLIT distance="1000" swimtime="00:13:37.00" />
                    <SPLIT distance="1050" swimtime="00:14:20.02" />
                    <SPLIT distance="1100" swimtime="00:15:02.75" />
                    <SPLIT distance="1150" swimtime="00:15:45.13" />
                    <SPLIT distance="1200" swimtime="00:16:27.75" />
                    <SPLIT distance="1250" swimtime="00:17:10.57" />
                    <SPLIT distance="1300" swimtime="00:17:53.09" />
                    <SPLIT distance="1350" swimtime="00:18:34.96" />
                    <SPLIT distance="1400" swimtime="00:19:17.18" />
                    <SPLIT distance="1450" swimtime="00:19:59.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-05-15" firstname="Łukasz" gender="M" lastname="Chmiel" nation="POL" athleteid="15047">
              <RESULTS>
                <RESULT eventid="1205" points="580" reactiontime="+67" swimtime="00:00:26.63" resultid="15048" heatid="19353" lane="5" entrytime="00:00:26.00" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="15049" heatid="19373" lane="5" />
                <RESULT eventid="14243" points="647" reactiontime="+71" swimtime="00:00:58.15" resultid="15050" heatid="19397" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="573" reactiontime="+74" swimtime="00:01:06.93" resultid="15051" heatid="19442" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="640" reactiontime="+70" swimtime="00:00:25.29" resultid="15052" heatid="19450" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-12-30" firstname="Krzysztof" gender="M" lastname="Krzak" nation="POL" athleteid="14634">
              <RESULTS>
                <RESULT eventid="1113" status="WDR" swimtime="00:00:00.00" resultid="14635" entrytime="00:02:44.87" />
                <RESULT eventid="14207" points="332" reactiontime="+107" swimtime="00:20:24.44" resultid="14636" heatid="19622" lane="4" entrytime="00:21:01.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.37" />
                    <SPLIT distance="100" swimtime="00:01:14.30" />
                    <SPLIT distance="150" swimtime="00:01:54.11" />
                    <SPLIT distance="200" swimtime="00:02:34.35" />
                    <SPLIT distance="250" swimtime="00:03:13.77" />
                    <SPLIT distance="300" swimtime="00:03:54.13" />
                    <SPLIT distance="350" swimtime="00:04:34.29" />
                    <SPLIT distance="400" swimtime="00:05:14.97" />
                    <SPLIT distance="450" swimtime="00:05:55.25" />
                    <SPLIT distance="500" swimtime="00:06:36.15" />
                    <SPLIT distance="550" swimtime="00:07:17.30" />
                    <SPLIT distance="600" swimtime="00:07:58.64" />
                    <SPLIT distance="650" swimtime="00:08:39.97" />
                    <SPLIT distance="700" swimtime="00:09:21.14" />
                    <SPLIT distance="750" swimtime="00:10:03.28" />
                    <SPLIT distance="800" swimtime="00:10:45.11" />
                    <SPLIT distance="850" swimtime="00:11:26.99" />
                    <SPLIT distance="900" swimtime="00:12:08.95" />
                    <SPLIT distance="950" swimtime="00:12:51.19" />
                    <SPLIT distance="1000" swimtime="00:13:33.18" />
                    <SPLIT distance="1050" swimtime="00:14:14.73" />
                    <SPLIT distance="1100" swimtime="00:14:56.60" />
                    <SPLIT distance="1150" swimtime="00:15:38.35" />
                    <SPLIT distance="1200" swimtime="00:16:20.46" />
                    <SPLIT distance="1250" swimtime="00:17:02.16" />
                    <SPLIT distance="1300" swimtime="00:17:43.47" />
                    <SPLIT distance="1350" swimtime="00:18:24.47" />
                    <SPLIT distance="1400" swimtime="00:19:05.57" />
                    <SPLIT distance="1450" swimtime="00:19:46.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="WDR" swimtime="00:00:00.00" resultid="14637" entrytime="00:00:35.41" />
                <RESULT eventid="14243" status="WDR" swimtime="00:00:00.00" resultid="14638" entrytime="00:01:13.08" />
                <RESULT eventid="1474" points="305" swimtime="00:01:12.61" resultid="14639" heatid="19475" lane="8" entrytime="00:01:17.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="331" reactiontime="+100" swimtime="00:05:40.38" resultid="14640" heatid="19510" lane="2" entrytime="00:05:59.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.45" />
                    <SPLIT distance="100" swimtime="00:01:21.02" />
                    <SPLIT distance="150" swimtime="00:02:05.30" />
                    <SPLIT distance="200" swimtime="00:02:47.47" />
                    <SPLIT distance="250" swimtime="00:03:34.58" />
                    <SPLIT distance="300" swimtime="00:04:23.86" />
                    <SPLIT distance="350" swimtime="00:05:03.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="306" reactiontime="+84" swimtime="00:02:36.70" resultid="14641" heatid="19535" lane="5" entrytime="00:02:43.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                    <SPLIT distance="100" swimtime="00:01:16.94" />
                    <SPLIT distance="150" swimtime="00:01:58.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="346" reactiontime="+105" swimtime="00:05:02.23" resultid="14642" heatid="19705" lane="4" entrytime="00:05:09.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.97" />
                    <SPLIT distance="100" swimtime="00:01:11.66" />
                    <SPLIT distance="150" swimtime="00:01:49.38" />
                    <SPLIT distance="200" swimtime="00:02:27.67" />
                    <SPLIT distance="250" swimtime="00:03:06.34" />
                    <SPLIT distance="300" swimtime="00:03:45.02" />
                    <SPLIT distance="350" swimtime="00:04:24.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-03-25" firstname="Jacek" gender="M" lastname="Kwiatkowski" nation="POL" athleteid="14665">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="14666" heatid="19289" lane="8" entrytime="00:00:33.52" />
                <RESULT eventid="14207" status="DNS" swimtime="00:00:00.00" resultid="14667" heatid="19621" lane="0" entrytime="00:24:51.00" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="14668" heatid="19508" lane="7" entrytime="00:07:10.00" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="14669" heatid="19702" lane="3" entrytime="00:06:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-18" firstname="Emil" gender="M" lastname="Strumiński" nation="POL" athleteid="14606">
              <RESULTS>
                <RESULT eventid="1079" points="432" reactiontime="+79" swimtime="00:00:26.80" resultid="14607" heatid="19299" lane="4" entrytime="00:00:26.80" />
                <RESULT eventid="1273" points="456" reactiontime="+80" swimtime="00:00:58.37" resultid="14608" heatid="19386" lane="0" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="14609" heatid="19460" lane="9" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-09-07" firstname="Tomasz" gender="M" lastname="Biadoń" nation="POL" athleteid="15972">
              <RESULTS>
                <RESULT eventid="1079" points="548" reactiontime="+73" swimtime="00:00:24.75" resultid="15973" heatid="19302" lane="5" entrytime="00:00:25.10" />
                <RESULT eventid="1273" points="508" reactiontime="+67" swimtime="00:00:56.30" resultid="15974" heatid="19386" lane="9" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="433" reactiontime="+67" swimtime="00:01:06.48" resultid="15975" heatid="19406" lane="8" entrytime="00:01:10.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="15976" heatid="19463" lane="2" entrytime="00:00:27.00" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="15977" heatid="19511" lane="3" entrytime="00:05:30.00" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="15978" heatid="19524" lane="2" entrytime="00:01:03.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-06-08" firstname="Wiesław" gender="M" lastname="Ciekliński" nation="POL" athleteid="18632">
              <RESULTS>
                <RESULT eventid="1079" points="258" reactiontime="+83" swimtime="00:00:31.80" resultid="18633" heatid="19290" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="14207" points="191" reactiontime="+106" swimtime="00:24:32.48" resultid="18634" heatid="19621" lane="7" entrytime="00:24:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.74" />
                    <SPLIT distance="200" swimtime="00:03:04.67" />
                    <SPLIT distance="250" swimtime="00:03:53.43" />
                    <SPLIT distance="300" swimtime="00:08:52.02" />
                    <SPLIT distance="350" swimtime="00:09:41.92" />
                    <SPLIT distance="400" swimtime="00:10:31.68" />
                    <SPLIT distance="450" swimtime="00:13:51.61" />
                    <SPLIT distance="500" swimtime="00:15:31.02" />
                    <SPLIT distance="550" swimtime="00:17:59.92" />
                    <SPLIT distance="600" swimtime="00:18:50.53" />
                    <SPLIT distance="650" swimtime="00:21:21.45" />
                    <SPLIT distance="700" swimtime="00:22:10.81" />
                    <SPLIT distance="750" swimtime="00:22:59.97" />
                    <SPLIT distance="1450" swimtime="00:23:48.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="236" reactiontime="+96" swimtime="00:01:12.62" resultid="18635" heatid="19379" lane="1" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="137" reactiontime="+92" swimtime="00:01:37.50" resultid="18636" heatid="19400" lane="6" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="18637" heatid="19453" lane="8" entrytime="00:00:38.00" />
                <RESULT eventid="1508" points="207" reactiontime="+92" swimtime="00:02:47.86" resultid="18638" heatid="19489" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.04" />
                    <SPLIT distance="100" swimtime="00:01:19.91" />
                    <SPLIT distance="150" swimtime="00:02:05.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="188" reactiontime="+103" swimtime="00:06:10.36" resultid="18639" heatid="19703" lane="0" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.68" />
                    <SPLIT distance="100" swimtime="00:02:16.07" />
                    <SPLIT distance="150" swimtime="00:03:03.93" />
                    <SPLIT distance="200" swimtime="00:03:51.42" />
                    <SPLIT distance="250" swimtime="00:04:39.52" />
                    <SPLIT distance="300" swimtime="00:05:27.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-16" firstname="Bartosz" gender="M" lastname="Rauczyński" nation="POL" athleteid="15043">
              <RESULTS>
                <RESULT eventid="1079" points="362" reactiontime="+87" swimtime="00:00:28.42" resultid="15044" heatid="19297" lane="1" entrytime="00:00:28.00" />
                <RESULT eventid="1341" points="279" reactiontime="+92" swimtime="00:02:46.09" resultid="15045" heatid="19416" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                    <SPLIT distance="100" swimtime="00:01:17.03" />
                    <SPLIT distance="150" swimtime="00:02:01.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="408" reactiontime="+93" swimtime="00:00:29.38" resultid="15046" heatid="19460" lane="3" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-11-14" firstname="Aleksandra" gender="F" lastname="Matraszek" nation="POL" athleteid="16537">
              <RESULTS>
                <RESULT eventid="1062" points="392" reactiontime="+89" swimtime="00:00:31.75" resultid="16538" heatid="19282" lane="7" entrytime="00:00:30.50" />
                <RESULT eventid="1096" points="297" reactiontime="+88" swimtime="00:03:02.53" resultid="16539" heatid="19308" lane="9" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.40" />
                    <SPLIT distance="100" swimtime="00:01:29.05" />
                    <SPLIT distance="150" swimtime="00:02:18.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="365" reactiontime="+91" swimtime="00:01:11.20" resultid="16540" heatid="19371" lane="3" entrytime="00:01:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="347" reactiontime="+97" swimtime="00:01:20.59" resultid="16541" heatid="19393" lane="2" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="348" reactiontime="+97" swimtime="00:01:28.62" resultid="16542" heatid="19431" lane="2" entrytime="00:01:27.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="315" reactiontime="+93" swimtime="00:02:42.68" resultid="16543" heatid="19483" lane="7" entrytime="00:02:45.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                    <SPLIT distance="100" swimtime="00:01:16.84" />
                    <SPLIT distance="150" swimtime="00:01:59.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="388" reactiontime="+94" swimtime="00:00:39.25" resultid="16544" heatid="19544" lane="3" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-07-18" firstname="Adrianna" gender="F" lastname="Buraczyńska" nation="POL" athleteid="16963">
              <RESULTS>
                <RESULT eventid="1147" status="DNS" swimtime="00:00:00.00" resultid="16964" heatid="19596" lane="1" entrytime="00:11:00.00" />
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="16965" heatid="19341" lane="1" entrytime="00:00:33.00" />
                <RESULT eventid="14225" status="DNS" swimtime="00:00:00.00" resultid="16966" heatid="19394" lane="4" entrytime="00:01:15.00" />
                <RESULT eventid="1457" points="462" reactiontime="+77" swimtime="00:01:11.18" resultid="16967" heatid="19469" lane="0" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="432" reactiontime="+80" swimtime="00:02:37.66" resultid="16968" heatid="19529" lane="3" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                    <SPLIT distance="100" swimtime="00:01:17.22" />
                    <SPLIT distance="150" swimtime="00:01:58.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-02-17" firstname="Piotr" gender="M" lastname="Kister" nation="POL" athleteid="14670">
              <RESULTS>
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="14671" heatid="19363" lane="6" entrytime="00:02:59.00" />
                <RESULT eventid="1341" points="272" reactiontime="+90" swimtime="00:02:47.49" resultid="14672" heatid="19417" lane="2" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                    <SPLIT distance="100" swimtime="00:01:14.78" />
                    <SPLIT distance="150" swimtime="00:01:58.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="295" reactiontime="+92" swimtime="00:01:23.49" resultid="14673" heatid="19440" lane="1" entrytime="00:01:19.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="333" reactiontime="+87" swimtime="00:00:31.43" resultid="14674" heatid="19458" lane="3" entrytime="00:00:30.99" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="14675" heatid="19522" lane="0" entrytime="00:01:11.00" />
                <RESULT eventid="1681" points="313" swimtime="00:00:37.15" resultid="14676" heatid="19555" lane="0" entrytime="00:00:36.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-03-16" firstname="Paweł" gender="M" lastname="Borkowski" nation="POL" athleteid="17138">
              <RESULTS>
                <RESULT eventid="1273" points="428" reactiontime="+96" swimtime="00:00:59.61" resultid="17139" heatid="19384" lane="7" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="388" reactiontime="+81" swimtime="00:02:16.16" resultid="17140" heatid="19493" lane="9" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.92" />
                    <SPLIT distance="100" swimtime="00:01:06.12" />
                    <SPLIT distance="150" swimtime="00:01:41.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-01-01" firstname="Mateusz" gender="M" lastname="Kwaśniewski" nation="POL" athleteid="14445">
              <RESULTS>
                <RESULT eventid="1079" points="534" reactiontime="+79" swimtime="00:00:24.96" resultid="14446" heatid="19303" lane="0" entrytime="00:00:25.00" />
                <RESULT eventid="14189" points="427" reactiontime="+75" swimtime="00:09:48.54" resultid="14447" heatid="19617" lane="6" entrytime="00:10:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.00" />
                    <SPLIT distance="100" swimtime="00:01:41.78" />
                    <SPLIT distance="200" swimtime="00:02:18.20" />
                    <SPLIT distance="250" swimtime="00:02:54.70" />
                    <SPLIT distance="300" swimtime="00:03:31.43" />
                    <SPLIT distance="350" swimtime="00:04:08.56" />
                    <SPLIT distance="400" swimtime="00:04:45.49" />
                    <SPLIT distance="450" swimtime="00:05:22.83" />
                    <SPLIT distance="500" swimtime="00:06:00.21" />
                    <SPLIT distance="550" swimtime="00:06:37.86" />
                    <SPLIT distance="600" swimtime="00:07:15.41" />
                    <SPLIT distance="650" swimtime="00:07:53.94" />
                    <SPLIT distance="700" swimtime="00:08:32.49" />
                    <SPLIT distance="750" swimtime="00:09:12.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="556" reactiontime="+77" swimtime="00:00:54.62" resultid="14448" heatid="19387" lane="3" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="532" reactiontime="+78" swimtime="00:00:26.89" resultid="14449" heatid="19463" lane="1" entrytime="00:00:27.00" />
                <RESULT eventid="1508" points="509" reactiontime="+78" swimtime="00:02:04.45" resultid="14450" heatid="19496" lane="2" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.28" />
                    <SPLIT distance="100" swimtime="00:00:58.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-04-25" firstname="Adriana" gender="F" lastname="Hofman" nation="POL" athleteid="15022">
              <RESULTS>
                <RESULT eventid="1388" points="509" reactiontime="+77" swimtime="00:01:18.06" resultid="15023" heatid="19432" lane="6" entrytime="00:01:20.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="513" reactiontime="+75" swimtime="00:00:35.76" resultid="15024" heatid="19545" lane="6" entrytime="00:00:35.75" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-05-18" firstname="Marcin" gender="M" lastname="Klimkowski" nation="POL" athleteid="15032">
              <RESULTS>
                <RESULT eventid="1474" points="16" swimtime="00:03:11.75" resultid="15033" heatid="19470" lane="2" entrytime="00:04:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:33.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="9" swimtime="00:07:50.10" resultid="15034" heatid="19486" lane="8" entrytime="00:08:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:45.83" />
                    <SPLIT distance="100" swimtime="00:03:47.99" />
                    <SPLIT distance="150" swimtime="00:05:52.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="18" swimtime="00:06:41.22" resultid="15035" heatid="19531" lane="8" entrytime="00:08:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:35.95" />
                    <SPLIT distance="100" swimtime="00:03:18.25" />
                    <SPLIT distance="150" swimtime="00:05:00.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="8" swimtime="00:02:01.68" resultid="15036" heatid="19547" lane="2" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-05-09" firstname="Łukasz" gender="M" lastname="Amanowicz" nation="POL" athleteid="14720">
              <RESULTS>
                <RESULT eventid="1079" points="266" reactiontime="+101" swimtime="00:00:31.48" resultid="14721" heatid="19286" lane="5" entrytime="00:00:38.00" />
                <RESULT eventid="1273" points="197" reactiontime="+96" swimtime="00:01:17.15" resultid="14722" heatid="19376" lane="9" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="148" swimtime="00:01:45.12" resultid="14723" heatid="19435" lane="0" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="179" reactiontime="+97" swimtime="00:00:44.75" resultid="14724" heatid="19548" lane="6" entrytime="00:00:53.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-08-29" firstname="Leszek" gender="M" lastname="Zawadzki" nation="POL" athleteid="14628">
              <RESULTS>
                <RESULT eventid="1079" points="289" reactiontime="+105" swimtime="00:00:30.62" resultid="14629" heatid="19297" lane="9" entrytime="00:00:28.05" />
                <RESULT eventid="14207" reactiontime="+137" status="OTL" swimtime="00:22:23.37" resultid="14630" heatid="19621" lane="5" entrytime="00:23:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                    <SPLIT distance="100" swimtime="00:01:13.66" />
                    <SPLIT distance="150" swimtime="00:01:55.53" />
                    <SPLIT distance="200" swimtime="00:02:39.20" />
                    <SPLIT distance="250" swimtime="00:03:22.69" />
                    <SPLIT distance="300" swimtime="00:04:06.34" />
                    <SPLIT distance="350" swimtime="00:04:49.91" />
                    <SPLIT distance="400" swimtime="00:05:33.63" />
                    <SPLIT distance="450" swimtime="00:06:17.71" />
                    <SPLIT distance="500" swimtime="00:07:03.06" />
                    <SPLIT distance="550" swimtime="00:07:46.96" />
                    <SPLIT distance="600" swimtime="00:08:31.54" />
                    <SPLIT distance="650" swimtime="00:09:16.08" />
                    <SPLIT distance="700" swimtime="00:10:00.79" />
                    <SPLIT distance="750" swimtime="00:10:47.06" />
                    <SPLIT distance="800" swimtime="00:11:31.70" />
                    <SPLIT distance="850" swimtime="00:12:16.94" />
                    <SPLIT distance="900" swimtime="00:13:02.33" />
                    <SPLIT distance="950" swimtime="00:13:47.71" />
                    <SPLIT distance="1000" swimtime="00:14:34.38" />
                    <SPLIT distance="1050" swimtime="00:15:20.23" />
                    <SPLIT distance="1100" swimtime="00:16:05.38" />
                    <SPLIT distance="1150" swimtime="00:16:54.28" />
                    <SPLIT distance="1200" swimtime="00:17:42.01" />
                    <SPLIT distance="1250" swimtime="00:18:29.32" />
                    <SPLIT distance="1300" swimtime="00:19:16.80" />
                    <SPLIT distance="1350" swimtime="00:20:03.65" />
                    <SPLIT distance="1400" swimtime="00:20:50.76" />
                    <SPLIT distance="1450" swimtime="00:21:39.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="270" reactiontime="+104" swimtime="00:01:09.47" resultid="14631" heatid="19384" lane="0" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="286" reactiontime="+110" swimtime="00:02:30.74" resultid="14632" heatid="19493" lane="5" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                    <SPLIT distance="100" swimtime="00:01:08.92" />
                    <SPLIT distance="150" swimtime="00:01:49.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="260" swimtime="00:05:32.50" resultid="14633" heatid="19705" lane="6" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                    <SPLIT distance="100" swimtime="00:01:12.35" />
                    <SPLIT distance="150" swimtime="00:01:51.88" />
                    <SPLIT distance="200" swimtime="00:02:33.35" />
                    <SPLIT distance="250" swimtime="00:03:16.79" />
                    <SPLIT distance="300" swimtime="00:04:02.66" />
                    <SPLIT distance="350" swimtime="00:04:48.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-06-20" firstname="Zbigniew" gender="M" lastname="Kapara" nation="POL" athleteid="15192">
              <RESULTS>
                <RESULT eventid="1273" points="189" reactiontime="+94" swimtime="00:01:18.21" resultid="15193" heatid="19378" lane="0" entrytime="00:01:17.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="127" reactiontime="+110" swimtime="00:01:39.92" resultid="15194" heatid="19397" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="133" reactiontime="+92" swimtime="00:00:42.69" resultid="15195" heatid="19450" lane="7" />
                <RESULT eventid="1508" points="130" reactiontime="+94" swimtime="00:03:15.95" resultid="15196" heatid="19487" lane="0" entrytime="00:03:39.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.41" />
                    <SPLIT distance="100" swimtime="00:01:28.32" />
                    <SPLIT distance="150" swimtime="00:02:19.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-03-11" firstname="Anna" gender="F" lastname="Głowiak" nation="POL" athleteid="14677">
              <RESULTS>
                <RESULT eventid="1062" points="375" reactiontime="+77" swimtime="00:00:32.22" resultid="14678" heatid="19279" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1187" points="272" swimtime="00:00:39.58" resultid="14679" heatid="19338" lane="1" entrytime="00:00:43.00" />
                <RESULT eventid="14225" points="299" reactiontime="+74" swimtime="00:01:24.72" resultid="14680" heatid="19392" lane="5" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="318" reactiontime="+79" swimtime="00:01:31.29" resultid="14681" heatid="19429" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="302" reactiontime="+79" swimtime="00:02:44.96" resultid="14682" heatid="19482" lane="5" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                    <SPLIT distance="100" swimtime="00:01:16.58" />
                    <SPLIT distance="150" swimtime="00:02:00.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="320" reactiontime="+76" swimtime="00:00:41.83" resultid="14683" heatid="19541" lane="3" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-09-23" firstname="Patrycja" gender="F" lastname="Sołtysiak" nation="POL" athleteid="15845">
              <RESULTS>
                <RESULT eventid="1222" points="410" reactiontime="+86" swimtime="00:03:01.01" resultid="15846" heatid="19358" lane="7" entrytime="00:03:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.74" />
                    <SPLIT distance="100" swimtime="00:01:26.49" />
                    <SPLIT distance="150" swimtime="00:02:14.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="422" reactiontime="+89" swimtime="00:01:23.11" resultid="15847" heatid="19432" lane="7" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="331" reactiontime="+81" swimtime="00:01:19.53" resultid="15848" heatid="19467" lane="4" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" status="DNS" swimtime="00:00:00.00" resultid="15849" heatid="19545" lane="1" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-08-13" firstname="Dmytro" gender="M" lastname="Bielskyi" nation="POL" athleteid="14276">
              <RESULTS>
                <RESULT eventid="1239" points="300" reactiontime="+100" swimtime="00:02:59.74" resultid="14277" heatid="19363" lane="1" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                    <SPLIT distance="100" swimtime="00:01:24.49" />
                    <SPLIT distance="150" swimtime="00:02:12.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="338" reactiontime="+91" swimtime="00:01:19.80" resultid="14278" heatid="19439" lane="5" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="336" reactiontime="+89" swimtime="00:00:36.29" resultid="14279" heatid="19555" lane="1" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-03-29" firstname="Mateusz" gender="M" lastname="Burzawa" nation="POL" athleteid="15013">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="15014" heatid="19301" lane="2" entrytime="00:00:26.00" />
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="15015" heatid="19318" lane="0" entrytime="00:02:20.00" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="15016" heatid="19351" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1239" points="451" reactiontime="+79" swimtime="00:02:36.96" resultid="15017" heatid="19364" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.55" />
                    <SPLIT distance="100" swimtime="00:01:15.71" />
                    <SPLIT distance="150" swimtime="00:01:55.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="15018" heatid="19441" lane="3" entrytime="00:01:13.00" />
                <RESULT eventid="1474" points="413" reactiontime="+66" swimtime="00:01:05.68" resultid="15019" heatid="19477" lane="5" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="15020" heatid="19537" lane="2" entrytime="00:02:25.00" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="15021" heatid="19558" lane="4" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-16" firstname="Wojciech" gender="M" lastname="Zmiejko" nation="POL" athleteid="14906">
              <RESULTS>
                <RESULT eventid="1079" points="384" reactiontime="+82" swimtime="00:00:27.87" resultid="14907" heatid="19297" lane="4" entrytime="00:00:27.95" />
                <RESULT eventid="1113" points="346" reactiontime="+90" swimtime="00:02:36.03" resultid="14908" heatid="19315" lane="1" entrytime="00:02:37.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                    <SPLIT distance="100" swimtime="00:01:13.16" />
                    <SPLIT distance="150" swimtime="00:02:00.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="380" reactiontime="+87" swimtime="00:01:02.04" resultid="14909" heatid="19383" lane="6" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="357" reactiontime="+90" swimtime="00:01:10.89" resultid="14910" heatid="19405" lane="4" entrytime="00:01:11.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="369" reactiontime="+90" swimtime="00:00:30.38" resultid="14911" heatid="19459" lane="0" entrytime="00:00:30.60" />
                <RESULT eventid="1474" points="283" reactiontime="+74" swimtime="00:01:14.49" resultid="14912" heatid="19475" lane="2" entrytime="00:01:15.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="343" reactiontime="+92" swimtime="00:01:08.66" resultid="14913" heatid="19522" lane="6" entrytime="00:01:09.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="262" reactiontime="+79" swimtime="00:02:45.00" resultid="14914" heatid="19535" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.56" />
                    <SPLIT distance="100" swimtime="00:01:20.61" />
                    <SPLIT distance="150" swimtime="00:02:02.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-02-12" firstname="Krzysztod" gender="M" lastname="Drózd" nation="POL" athleteid="14601">
              <RESULTS>
                <RESULT eventid="1205" points="315" reactiontime="+88" swimtime="00:00:32.63" resultid="14602" heatid="19349" lane="0" entrytime="00:00:34.00" />
                <RESULT eventid="1273" points="376" reactiontime="+77" swimtime="00:01:02.24" resultid="14603" heatid="19383" lane="4" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="320" reactiontime="+68" swimtime="00:01:11.50" resultid="14604" heatid="19470" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="14605" heatid="19491" lane="6" entrytime="00:02:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-06-28" firstname="Bolewław" gender="M" lastname="Czyż" nation="POL" athleteid="17141">
              <RESULTS>
                <RESULT eventid="1341" points="65" reactiontime="+118" swimtime="00:04:29.23" resultid="17142" heatid="19414" lane="2" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.59" />
                    <SPLIT distance="100" swimtime="00:02:12.08" />
                    <SPLIT distance="150" swimtime="00:03:21.96" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K16 - Niejednoczesne dotknięcie ściany dłońmi przy nawrocie lub na zakończenie wyścigu (Time: 20:45)" eventid="1578" reactiontime="+111" status="DSQ" swimtime="00:08:41.66" resultid="17143" heatid="19507" lane="4" entrytime="00:08:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.47" />
                    <SPLIT distance="100" swimtime="00:02:08.06" />
                    <SPLIT distance="150" swimtime="00:03:13.74" />
                    <SPLIT distance="200" swimtime="00:04:19.76" />
                    <SPLIT distance="250" swimtime="00:05:31.22" />
                    <SPLIT distance="300" swimtime="00:06:41.23" />
                    <SPLIT distance="350" swimtime="00:07:41.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-02-18" firstname="Kazimierz" gender="M" lastname="Sinicki" nation="POL" athleteid="14272">
              <RESULTS>
                <RESULT eventid="1079" points="321" reactiontime="+81" swimtime="00:00:29.57" resultid="14273" heatid="19292" lane="7" entrytime="00:00:30.21" />
                <RESULT eventid="1273" points="280" reactiontime="+84" swimtime="00:01:08.65" resultid="14274" heatid="19380" lane="6" entrytime="00:01:08.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="251" reactiontime="+84" swimtime="00:00:34.52" resultid="14275" heatid="19454" lane="9" entrytime="00:00:36.21" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-12-31" firstname="Piotr" gender="M" lastname="Żuczek" nation="POL" athleteid="18954">
              <RESULTS>
                <RESULT eventid="1239" points="430" reactiontime="+87" swimtime="00:02:39.56" resultid="18955" heatid="19365" lane="2" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.69" />
                    <SPLIT distance="100" swimtime="00:01:14.50" />
                    <SPLIT distance="150" swimtime="00:01:55.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="490" reactiontime="+77" swimtime="00:01:10.53" resultid="18956" heatid="19442" lane="6" entrytime="00:01:09.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="399" reactiontime="+63" swimtime="00:01:06.41" resultid="18957" heatid="19478" lane="9" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="351" reactiontime="+71" swimtime="00:02:29.72" resultid="18958" heatid="19536" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.95" />
                    <SPLIT distance="100" swimtime="00:01:12.83" />
                    <SPLIT distance="150" swimtime="00:01:51.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="487" reactiontime="+79" swimtime="00:00:32.08" resultid="18959" heatid="19559" lane="3" entrytime="00:00:31.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-08-26" firstname="Adrian" gender="M" lastname="Kozioł" nation="POL" athleteid="16221">
              <RESULTS>
                <RESULT eventid="1079" points="395" reactiontime="+81" swimtime="00:00:27.60" resultid="16222" heatid="19296" lane="3" entrytime="00:00:28.50" />
                <RESULT eventid="1440" points="395" reactiontime="+82" swimtime="00:00:29.71" resultid="16223" heatid="19458" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="1508" points="275" reactiontime="+81" swimtime="00:02:32.76" resultid="16224" heatid="19491" lane="8" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                    <SPLIT distance="100" swimtime="00:01:10.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-05-20" firstname="Łukasz" gender="M" lastname="Popławski" nation="POL" athleteid="16259">
              <RESULTS>
                <RESULT eventid="14207" reactiontime="+78" status="OTL" swimtime="00:20:06.65" resultid="16260" heatid="19623" lane="8" entrytime="00:20:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                    <SPLIT distance="100" swimtime="00:01:11.30" />
                    <SPLIT distance="200" swimtime="00:02:29.66" />
                    <SPLIT distance="250" swimtime="00:03:10.32" />
                    <SPLIT distance="300" swimtime="00:03:51.17" />
                    <SPLIT distance="350" swimtime="00:04:31.77" />
                    <SPLIT distance="400" swimtime="00:05:13.62" />
                    <SPLIT distance="450" swimtime="00:05:54.33" />
                    <SPLIT distance="550" swimtime="00:07:15.73" />
                    <SPLIT distance="650" swimtime="00:08:36.53" />
                    <SPLIT distance="700" swimtime="00:09:16.71" />
                    <SPLIT distance="750" swimtime="00:09:57.62" />
                    <SPLIT distance="850" swimtime="00:11:20.12" />
                    <SPLIT distance="950" swimtime="00:12:40.94" />
                    <SPLIT distance="1000" swimtime="00:13:21.82" />
                    <SPLIT distance="1050" swimtime="00:14:02.94" />
                    <SPLIT distance="1150" swimtime="00:15:25.43" />
                    <SPLIT distance="1200" swimtime="00:16:07.15" />
                    <SPLIT distance="1250" swimtime="00:16:47.59" />
                    <SPLIT distance="1300" swimtime="00:17:28.23" />
                    <SPLIT distance="1350" swimtime="00:18:08.67" />
                    <SPLIT distance="1400" swimtime="00:18:49.48" />
                    <SPLIT distance="1450" swimtime="00:19:28.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="426" reactiontime="+77" swimtime="00:02:40.06" resultid="16261" heatid="19365" lane="8" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                    <SPLIT distance="100" swimtime="00:01:16.10" />
                    <SPLIT distance="150" swimtime="00:01:57.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="425" reactiontime="+80" swimtime="00:01:13.94" resultid="16262" heatid="19441" lane="2" entrytime="00:01:13.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="393" reactiontime="+76" swimtime="00:05:21.45" resultid="16263" heatid="19512" lane="9" entrytime="00:05:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                    <SPLIT distance="100" swimtime="00:01:11.27" />
                    <SPLIT distance="150" swimtime="00:01:55.84" />
                    <SPLIT distance="200" swimtime="00:02:39.22" />
                    <SPLIT distance="250" swimtime="00:03:23.01" />
                    <SPLIT distance="300" swimtime="00:04:07.27" />
                    <SPLIT distance="350" swimtime="00:04:45.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="406" reactiontime="+80" swimtime="00:00:34.09" resultid="16264" heatid="19557" lane="7" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-10-28" firstname="Robert" gender="M" lastname="Drzazga" nation="POL" athleteid="14262">
              <RESULTS>
                <RESULT eventid="1273" points="283" reactiontime="+83" swimtime="00:01:08.41" resultid="14263" heatid="19378" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="235" reactiontime="+87" swimtime="00:01:21.48" resultid="14264" heatid="19399" lane="4" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="266" reactiontime="+86" swimtime="00:00:33.86" resultid="14265" heatid="19454" lane="7" entrytime="00:00:35.50" />
                <RESULT eventid="1508" points="266" reactiontime="+88" swimtime="00:02:34.47" resultid="14266" heatid="19489" lane="0" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                    <SPLIT distance="100" swimtime="00:01:12.53" />
                    <SPLIT distance="150" swimtime="00:01:53.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-27" firstname="Marta" gender="F" lastname="Sołtysiak" nation="POL" athleteid="15840">
              <RESULTS>
                <RESULT eventid="1187" points="289" reactiontime="+77" swimtime="00:00:38.82" resultid="15841" heatid="19338" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="1256" points="298" reactiontime="+100" swimtime="00:01:16.16" resultid="15842" heatid="19369" lane="2" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="266" reactiontime="+76" swimtime="00:01:25.48" resultid="15843" heatid="19466" lane="4" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" status="DNS" swimtime="00:00:00.00" resultid="15844" heatid="19527" lane="5" entrytime="00:03:15.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="UKR" clubid="18471" name="Niezrzeszeni UKR">
          <ATHLETES>
            <ATHLETE birthdate="1980-11-16" firstname="Yurii" gender="M" lastname="VASHCHUK" nation="POL" athleteid="17135">
              <RESULTS>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="17136" heatid="19457" lane="8" entrytime="00:00:32.00" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="17137" heatid="19558" lane="2" entrytime="00:00:32.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="UKR" clubid="17658" name="No Stars">
          <CONTACT city="Chernigiv" email="nostarsswimming@gmail.com" name="Kutueva Olga" phone="+38 050 4651785" street="Rokossovskiy str 17A/36" zip="14000" />
          <ATHLETES>
            <ATHLETE birthdate="1970-05-27" firstname="Oleksandr" gender="M" lastname="Zubets" nation="UKR" athleteid="17668">
              <RESULTS>
                <RESULT eventid="1079" points="426" reactiontime="+77" swimtime="00:00:26.91" resultid="17669" heatid="19299" lane="3" entrytime="00:00:27.00" />
                <RESULT eventid="1113" points="300" reactiontime="+75" swimtime="00:02:43.59" resultid="17670" heatid="19314" lane="7" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                    <SPLIT distance="100" swimtime="00:01:12.20" />
                    <SPLIT distance="150" swimtime="00:02:03.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="444" reactiontime="+71" swimtime="00:00:58.88" resultid="17671" heatid="19384" lane="8" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="389" reactiontime="+76" swimtime="00:01:08.90" resultid="17672" heatid="19404" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="410" reactiontime="+69" swimtime="00:00:29.33" resultid="17673" heatid="19460" lane="5" entrytime="00:00:29.00" />
                <RESULT eventid="1508" points="383" reactiontime="+63" swimtime="00:02:16.74" resultid="17674" heatid="19492" lane="9" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.36" />
                    <SPLIT distance="100" swimtime="00:01:04.43" />
                    <SPLIT distance="150" swimtime="00:01:41.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="358" reactiontime="+72" swimtime="00:01:07.65" resultid="17675" heatid="19521" lane="5" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="17676" heatid="19552" lane="7" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-05" firstname="Sergii" gender="M" lastname="Mezherytskyi" nation="UKR" athleteid="17677">
              <RESULTS>
                <RESULT eventid="1079" points="390" reactiontime="+81" swimtime="00:00:27.73" resultid="17678" heatid="19299" lane="5" entrytime="00:00:26.80" />
                <RESULT eventid="1113" points="310" reactiontime="+85" swimtime="00:02:41.90" resultid="17679" heatid="19314" lane="1" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                    <SPLIT distance="100" swimtime="00:01:18.39" />
                    <SPLIT distance="150" swimtime="00:02:04.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="402" reactiontime="+77" swimtime="00:01:00.89" resultid="17680" heatid="19384" lane="6" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="349" reactiontime="+84" swimtime="00:00:30.94" resultid="17681" heatid="19459" lane="1" entrytime="00:00:30.50" />
                <RESULT eventid="1508" points="314" reactiontime="+79" swimtime="00:02:26.13" resultid="17682" heatid="19491" lane="4" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                    <SPLIT distance="100" swimtime="00:01:11.33" />
                    <SPLIT distance="150" swimtime="00:01:49.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="311" reactiontime="+80" swimtime="00:01:10.90" resultid="17683" heatid="19521" lane="3" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ORS OPOLE" nation="POL" region="OPO" clubid="15434" name="ORS Opole">
          <CONTACT name="Stanek" street="Wojciech" />
          <ATHLETES>
            <ATHLETE birthdate="1992-01-01" firstname="Wojciech" gender="M" lastname="Stanek" nation="POL" athleteid="15435">
              <RESULTS>
                <RESULT comment="O4 - Start wykonany przed sygnłem (przedwczesny start) (Time: 16:29)" eventid="1113" reactiontime="+62" status="DSQ" swimtime="00:02:36.83" resultid="15436" heatid="19313" lane="7" entrytime="00:02:48.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.92" />
                    <SPLIT distance="100" swimtime="00:01:16.07" />
                    <SPLIT distance="150" swimtime="00:02:00.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="15437" heatid="19380" lane="9" entrytime="00:01:09.50" />
                <RESULT eventid="1578" points="346" reactiontime="+84" swimtime="00:05:35.19" resultid="15438" heatid="19509" lane="5" entrytime="00:06:08.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.83" />
                    <SPLIT distance="100" swimtime="00:01:20.56" />
                    <SPLIT distance="150" swimtime="00:02:03.62" />
                    <SPLIT distance="200" swimtime="00:02:46.01" />
                    <SPLIT distance="250" swimtime="00:03:33.31" />
                    <SPLIT distance="300" swimtime="00:04:19.75" />
                    <SPLIT distance="350" swimtime="00:04:58.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="15439" heatid="19705" lane="7" entrytime="00:05:12.40" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="SLA" clubid="15312" name="Park Wodny Tarnowskie Góry Masters" shortname="Park Wodny Tarnowskie Góry Mas">
          <CONTACT city="Tarnowskie Góry" email="swimman@o2.pl" name="Pąchalski Tomasz" phone="600-365-944" state="SLA" street="Obwodnica 8" zip="42-600" />
          <ATHLETES>
            <ATHLETE birthdate="1966-12-12" firstname="Barbara" gender="F" lastname="Czichy" nation="POL" athleteid="15352">
              <RESULTS>
                <RESULT eventid="1388" points="148" reactiontime="+112" swimtime="00:01:57.72" resultid="15353" heatid="19427" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="162" reactiontime="+110" swimtime="00:00:52.48" resultid="15354" heatid="19538" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-28" firstname="Michał" gender="M" lastname="Grzybczyk" nation="POL" athleteid="15342">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="15343" heatid="19289" lane="0" entrytime="00:00:34.00" />
                <RESULT eventid="1273" reactiontime="+137" status="DNS" swimtime="00:00:00.00" resultid="15344" heatid="19374" lane="0" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-04-14" firstname="Katarzyna" gender="F" lastname="Sowa" nation="POL" athleteid="15340">
              <RESULTS>
                <RESULT eventid="1721" points="205" reactiontime="+81" swimtime="00:06:37.43" resultid="15341" heatid="19696" lane="7" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.79" />
                    <SPLIT distance="100" swimtime="00:01:30.46" />
                    <SPLIT distance="150" swimtime="00:02:20.65" />
                    <SPLIT distance="200" swimtime="00:03:11.71" />
                    <SPLIT distance="250" swimtime="00:04:02.73" />
                    <SPLIT distance="300" swimtime="00:04:54.86" />
                    <SPLIT distance="350" swimtime="00:05:47.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-21" firstname="Marta" gender="F" lastname="Ginko" nation="POL" athleteid="15364" />
            <ATHLETE birthdate="1975-08-09" firstname="Sonia" gender="F" lastname="Borkowska" nation="POL" athleteid="15345">
              <RESULTS>
                <RESULT eventid="1062" points="378" reactiontime="+78" swimtime="00:00:32.13" resultid="15346" heatid="19280" lane="5" entrytime="00:00:33.15" />
                <RESULT eventid="1256" points="332" reactiontime="+77" swimtime="00:01:13.51" resultid="15347" heatid="19370" lane="6" entrytime="00:01:15.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="277" reactiontime="+73" swimtime="00:01:26.92" resultid="15348" heatid="19391" lane="4" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="276" reactiontime="+80" swimtime="00:00:37.44" resultid="15349" heatid="19446" lane="8" entrytime="00:00:40.10" />
                <RESULT eventid="1491" points="282" reactiontime="+86" swimtime="00:02:48.89" resultid="15350" heatid="19482" lane="6" entrytime="00:02:55.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                    <SPLIT distance="100" swimtime="00:01:18.89" />
                    <SPLIT distance="150" swimtime="00:02:04.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="315" reactiontime="+81" swimtime="00:00:42.07" resultid="15351" heatid="19542" lane="6" entrytime="00:00:42.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-08-07" firstname="Mirosław" gender="M" lastname="Gondek" nation="POL" athleteid="15360">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="15361" heatid="19287" lane="0" entrytime="00:00:38.00" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="15362" heatid="19377" lane="2" entrytime="00:01:20.00" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="15363" heatid="19452" lane="2" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-10-03" firstname="Tomasz" gender="M" lastname="Pąchalski" nation="POL" athleteid="19748" />
            <ATHLETE birthdate="1977-10-10" firstname="Krzysztof" gender="M" lastname="Dyr" nation="POL" athleteid="15355">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="15356" heatid="19284" lane="9" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="15357" heatid="19546" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-07-26" firstname="Marta" gender="F" lastname="Oracz" nation="POL" athleteid="15337">
              <RESULTS>
                <RESULT eventid="1147" status="DNF" swimtime="00:00:00.00" resultid="15338" heatid="19595" lane="0" entrytime="00:15:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.79" />
                    <SPLIT distance="100" swimtime="00:01:32.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="240" reactiontime="+95" swimtime="00:06:16.94" resultid="15339" heatid="19696" lane="0" entrytime="00:07:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.04" />
                    <SPLIT distance="100" swimtime="00:01:31.47" />
                    <SPLIT distance="150" swimtime="00:02:21.13" />
                    <SPLIT distance="200" swimtime="00:03:08.31" />
                    <SPLIT distance="250" swimtime="00:03:56.51" />
                    <SPLIT distance="300" swimtime="00:04:44.01" />
                    <SPLIT distance="350" swimtime="00:05:31.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-02-27" firstname="Rafał" gender="M" lastname="Domeracki" nation="POL" athleteid="15332">
              <RESULTS>
                <RESULT eventid="14207" reactiontime="+92" status="OTL" swimtime="00:21:51.47" resultid="15333" heatid="19622" lane="5" entrytime="00:21:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.45" />
                    <SPLIT distance="100" swimtime="00:01:20.16" />
                    <SPLIT distance="150" swimtime="00:02:01.94" />
                    <SPLIT distance="200" swimtime="00:02:45.97" />
                    <SPLIT distance="250" swimtime="00:03:28.27" />
                    <SPLIT distance="300" swimtime="00:04:12.99" />
                    <SPLIT distance="350" swimtime="00:04:56.06" />
                    <SPLIT distance="400" swimtime="00:05:39.54" />
                    <SPLIT distance="450" swimtime="00:06:22.89" />
                    <SPLIT distance="500" swimtime="00:07:06.01" />
                    <SPLIT distance="550" swimtime="00:07:50.11" />
                    <SPLIT distance="600" swimtime="00:08:35.07" />
                    <SPLIT distance="650" swimtime="00:09:18.26" />
                    <SPLIT distance="700" swimtime="00:10:03.44" />
                    <SPLIT distance="750" swimtime="00:10:48.65" />
                    <SPLIT distance="800" swimtime="00:11:32.34" />
                    <SPLIT distance="850" swimtime="00:12:16.09" />
                    <SPLIT distance="900" swimtime="00:13:00.15" />
                    <SPLIT distance="950" swimtime="00:13:43.94" />
                    <SPLIT distance="1000" swimtime="00:14:29.34" />
                    <SPLIT distance="1050" swimtime="00:15:13.59" />
                    <SPLIT distance="1100" swimtime="00:15:58.02" />
                    <SPLIT distance="1150" swimtime="00:16:42.38" />
                    <SPLIT distance="1200" swimtime="00:17:26.74" />
                    <SPLIT distance="1250" swimtime="00:18:12.07" />
                    <SPLIT distance="1300" swimtime="00:18:57.06" />
                    <SPLIT distance="1350" swimtime="00:19:40.73" />
                    <SPLIT distance="1400" swimtime="00:20:24.82" />
                    <SPLIT distance="1450" swimtime="00:21:08.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="248" reactiontime="+89" swimtime="00:01:11.51" resultid="15334" heatid="19378" lane="3" entrytime="00:01:14.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="278" reactiontime="+113" swimtime="00:02:32.15" resultid="15335" heatid="19491" lane="2" entrytime="00:02:31.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                    <SPLIT distance="100" swimtime="00:01:14.59" />
                    <SPLIT distance="150" swimtime="00:01:53.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="289" reactiontime="+96" swimtime="00:05:21.00" resultid="15336" heatid="19704" lane="2" entrytime="00:05:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                    <SPLIT distance="100" swimtime="00:01:16.79" />
                    <SPLIT distance="150" swimtime="00:01:57.16" />
                    <SPLIT distance="200" swimtime="00:02:38.58" />
                    <SPLIT distance="250" swimtime="00:03:19.39" />
                    <SPLIT distance="300" swimtime="00:04:00.84" />
                    <SPLIT distance="350" swimtime="00:04:41.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-09-09" firstname="Anna" gender="F" lastname="Chmiel" nation="POL" athleteid="15358">
              <RESULTS>
                <RESULT eventid="1256" points="213" reactiontime="+132" swimtime="00:01:25.24" resultid="15359" heatid="19366" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" status="DNS" swimtime="00:00:00.00" resultid="15369" heatid="19499" lane="1">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15342" number="1" />
                    <RELAYPOSITION athleteid="15360" number="2" />
                    <RELAYPOSITION athleteid="15355" number="3" />
                    <RELAYPOSITION athleteid="15332" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT comment="S4 - Przedwczesna zmiana sztafetowa (stopy pływaka utraciły kontakt z platformą startową słupka zanim poprzedzający go pływak dotkną ściany) (Time: 19:30), Na pierwszej zmianie" eventid="1525" reactiontime="+141" status="DSQ" swimtime="00:02:24.21" resultid="15367" heatid="19497" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.04" />
                    <SPLIT distance="100" swimtime="00:01:15.91" />
                    <SPLIT distance="150" swimtime="00:01:52.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15358" number="1" reactiontime="+141" />
                    <RELAYPOSITION athleteid="15340" number="2" reactiontime="-23" status="DSQ" />
                    <RELAYPOSITION athleteid="15337" number="3" reactiontime="+73" status="DSQ" />
                    <RELAYPOSITION athleteid="15345" number="4" reactiontime="+50" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1358" points="145" reactiontime="+83" swimtime="00:03:16.34" resultid="15368" heatid="19419" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.01" />
                    <SPLIT distance="100" swimtime="00:01:51.32" />
                    <SPLIT distance="150" swimtime="00:02:39.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15364" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="15352" number="2" reactiontime="+94" />
                    <RELAYPOSITION athleteid="15337" number="3" reactiontime="+73" />
                    <RELAYPOSITION athleteid="15358" number="4" reactiontime="+72" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1698" status="DNS" swimtime="00:00:00.00" resultid="15365" heatid="19561" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15340" number="1" />
                    <RELAYPOSITION athleteid="15332" number="2" />
                    <RELAYPOSITION athleteid="15360" number="3" />
                    <RELAYPOSITION athleteid="15345" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1130" status="DNS" swimtime="00:00:00.00" resultid="15366" heatid="19319" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15345" number="1" />
                    <RELAYPOSITION athleteid="15337" number="2" />
                    <RELAYPOSITION athleteid="15360" number="3" />
                    <RELAYPOSITION athleteid="15332" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="PAŁAC" nation="POL" region="SLA" clubid="15989" name="Pałac Katowice Masters">
          <CONTACT name="Bucholz" phone="606135860" />
          <ATHLETES>
            <ATHLETE birthdate="1973-11-08" firstname="Piotr" gender="M" lastname="Przebindowski" nation="POL" athleteid="15994" />
            <ATHLETE birthdate="1972-01-26" firstname="Tomasz" gender="M" lastname="Bucholz" nation="POL" athleteid="15990">
              <RESULTS>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="15991" heatid="19492" lane="5" entrytime="00:02:23.00" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="15992" heatid="19705" lane="9" entrytime="00:05:17.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-05-02" firstname="Mateusz" gender="M" lastname="Matysiewicz" nation="POL" athleteid="15995" />
            <ATHLETE birthdate="1973-08-28" firstname="jacek" gender="M" lastname="Kobylczak" nation="POL" athleteid="15993" />
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" status="DNS" swimtime="00:00:00.00" resultid="15996" heatid="19501" lane="9" entrytime="00:02:03.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15993" number="1" />
                    <RELAYPOSITION athleteid="15995" number="2" />
                    <RELAYPOSITION athleteid="15994" number="3" />
                    <RELAYPOSITION athleteid="15990" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" points="293" reactiontime="+62" swimtime="00:02:16.12" resultid="15997" heatid="19422" lane="5" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                    <SPLIT distance="100" swimtime="00:00:55.65" />
                    <SPLIT distance="150" swimtime="00:01:47.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15994" number="1" reactiontime="+62" />
                    <RELAYPOSITION athleteid="15995" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="15990" number="3" />
                    <RELAYPOSITION athleteid="15993" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="107" nation="SVK" clubid="15914" name="PKM Turčianski raci">
          <CONTACT city="Vrútky" email="chrapco@gmail.com" name="Branislav Turanský" phone="+421903942831" street="Horná 34" zip="03861" />
          <ATHLETES>
            <ATHLETE birthdate="1967-12-18" firstname="Branislav" gender="M" lastname="Turanský" nation="SVK" license="SVK13190" athleteid="15922">
              <RESULTS>
                <RESULT eventid="1079" points="416" reactiontime="+76" swimtime="00:00:27.12" resultid="15923" heatid="19298" lane="8" entrytime="00:00:27.63" />
                <RESULT eventid="1113" points="321" reactiontime="+91" swimtime="00:02:40.06" resultid="15924" heatid="19313" lane="1" entrytime="00:02:49.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.07" />
                    <SPLIT distance="100" swimtime="00:01:14.89" />
                    <SPLIT distance="150" swimtime="00:02:03.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="395" reactiontime="+85" swimtime="00:01:01.22" resultid="15925" heatid="19384" lane="5" entrytime="00:01:00.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="332" reactiontime="+74" swimtime="00:01:10.63" resultid="15926" heatid="19476" lane="2" entrytime="00:01:11.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="289" reactiontime="+89" swimtime="00:05:56.19" resultid="15927" heatid="19510" lane="5" entrytime="00:05:57.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.04" />
                    <SPLIT distance="100" swimtime="00:01:19.49" />
                    <SPLIT distance="150" swimtime="00:02:03.35" />
                    <SPLIT distance="200" swimtime="00:02:46.98" />
                    <SPLIT distance="250" swimtime="00:03:40.72" />
                    <SPLIT distance="300" swimtime="00:04:34.44" />
                    <SPLIT distance="350" swimtime="00:05:17.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="316" reactiontime="+65" swimtime="00:02:34.92" resultid="15928" heatid="19536" lane="2" entrytime="00:02:36.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                    <SPLIT distance="100" swimtime="00:01:14.49" />
                    <SPLIT distance="150" swimtime="00:01:54.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-02-18" firstname="Lívia" gender="F" lastname="Velitsová" nation="SVK" license="SVK18938" athleteid="15959">
              <RESULTS>
                <RESULT eventid="1222" points="166" reactiontime="+134" swimtime="00:04:04.50" resultid="15960" heatid="19355" lane="3" entrytime="00:04:19.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.38" />
                    <SPLIT distance="100" swimtime="00:01:57.39" />
                    <SPLIT distance="150" swimtime="00:03:00.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="176" reactiontime="+129" swimtime="00:01:51.13" resultid="15961" heatid="19428" lane="7" entrytime="00:01:57.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="193" reactiontime="+132" swimtime="00:00:49.48" resultid="15962" heatid="19540" lane="3" entrytime="00:00:50.51" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-06-16" firstname="Katarína" gender="F" lastname="Turanská" nation="SVK" license="SVK17844" athleteid="15929">
              <RESULTS>
                <RESULT eventid="1062" points="114" reactiontime="+103" swimtime="00:00:47.87" resultid="15930" heatid="19276" lane="1" entrytime="00:00:50.54" />
                <RESULT eventid="1222" points="181" reactiontime="+115" swimtime="00:03:57.67" resultid="15931" heatid="19355" lane="4" entrytime="00:04:10.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.77" />
                    <SPLIT distance="100" swimtime="00:01:55.75" />
                    <SPLIT distance="150" swimtime="00:02:57.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="81" reactiontime="+88" swimtime="00:00:56.16" resultid="15932" heatid="19445" lane="8" entrytime="00:00:56.24" />
                <RESULT eventid="1664" points="191" reactiontime="+100" swimtime="00:00:49.65" resultid="15933" heatid="19540" lane="7" entrytime="00:00:51.45" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-11-26" firstname="Darina" gender="F" lastname="Krausová" nation="SVK" license="SVK20932" athleteid="15963">
              <RESULTS>
                <RESULT eventid="1595" points="240" reactiontime="+72" swimtime="00:01:27.86" resultid="15964" heatid="19515" lane="0" entrytime="00:01:23.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-05-10" firstname="Miroslav" gender="M" lastname="Kočalka" nation="SVK" license="SVK17837" athleteid="15918">
              <RESULTS>
                <RESULT eventid="1273" points="131" reactiontime="+88" swimtime="00:01:28.34" resultid="15919" heatid="19376" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="168" reactiontime="+85" swimtime="00:00:39.46" resultid="15920" heatid="19453" lane="1" entrytime="00:00:37.31" />
                <RESULT comment="O4 - Start wykonany przed sygnłem (przedwczesny start) (Time: 9:20)" eventid="1613" reactiontime="+61" status="DSQ" swimtime="00:01:29.98" resultid="15921" heatid="19519" lane="7" entrytime="00:01:29.24" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-02-16" firstname="Ladislav" gender="M" lastname="Zvarík" nation="SVK" license="SVK17846" athleteid="15915">
              <RESULTS>
                <RESULT eventid="1406" points="119" reactiontime="+115" swimtime="00:01:52.87" resultid="15916" heatid="19435" lane="1" entrytime="00:01:53.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="142" reactiontime="+105" swimtime="00:00:48.38" resultid="15917" heatid="19549" lane="7" entrytime="00:00:47.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-06-08" firstname="Ján" gender="M" lastname="Vanko" nation="SVK" license="SVK17842" athleteid="15934">
              <RESULTS>
                <RESULT eventid="1079" points="202" reactiontime="+106" swimtime="00:00:34.51" resultid="15935" heatid="19288" lane="4" entrytime="00:00:34.60" />
                <RESULT eventid="1113" points="136" reactiontime="+102" swimtime="00:03:32.93" resultid="15936" heatid="19311" lane="7" entrytime="00:03:35.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.06" />
                    <SPLIT distance="100" swimtime="00:01:40.84" />
                    <SPLIT distance="150" swimtime="00:02:44.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="120" reactiontime="+94" swimtime="00:00:45.03" resultid="15937" heatid="19345" lane="1" entrytime="00:00:44.58" />
                <RESULT eventid="14243" points="153" reactiontime="+103" swimtime="00:01:33.92" resultid="15938" heatid="19399" lane="1" entrytime="00:01:40.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="180" reactiontime="+90" swimtime="00:00:38.58" resultid="15939" heatid="19452" lane="3" entrytime="00:00:40.93" />
                <RESULT eventid="1647" points="84" reactiontime="+89" swimtime="00:04:00.70" resultid="15940" heatid="19532" lane="6" entrytime="00:04:09.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.02" />
                    <SPLIT distance="100" swimtime="00:01:51.80" />
                    <SPLIT distance="150" swimtime="00:02:55.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-02-03" firstname="Adriana" gender="F" lastname="Salaiová" nation="SVK" license="SVK17833" athleteid="15944">
              <RESULTS>
                <RESULT eventid="1062" points="56" swimtime="00:01:00.43" resultid="15945" heatid="19276" lane="9" entrytime="00:01:00.89" />
                <RESULT eventid="1256" points="53" reactiontime="+117" swimtime="00:02:15.05" resultid="15946" heatid="19367" lane="6" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="96" reactiontime="+138" swimtime="00:01:02.50" resultid="15947" heatid="19539" lane="2" entrytime="00:01:06.21" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-12-26" firstname="Michaela" gender="F" lastname="Janovská" nation="SVK" license="SVK21011" athleteid="15954">
              <RESULTS>
                <RESULT eventid="14225" points="234" reactiontime="+84" swimtime="00:01:31.94" resultid="15955" heatid="19391" lane="3" entrytime="00:01:34.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="188" reactiontime="+83" swimtime="00:00:42.52" resultid="15956" heatid="19446" lane="0" entrytime="00:00:43.27" />
                <RESULT eventid="1491" points="229" reactiontime="+115" swimtime="00:03:01.01" resultid="15957" heatid="19481" lane="5" entrytime="00:03:05.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.69" />
                    <SPLIT distance="100" swimtime="00:01:23.65" />
                    <SPLIT distance="150" swimtime="00:02:12.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="232" reactiontime="+91" swimtime="00:06:21.22" resultid="15958" heatid="19696" lane="6" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.78" />
                    <SPLIT distance="100" swimtime="00:01:27.08" />
                    <SPLIT distance="150" swimtime="00:02:14.54" />
                    <SPLIT distance="200" swimtime="00:03:03.16" />
                    <SPLIT distance="250" swimtime="00:03:52.27" />
                    <SPLIT distance="300" swimtime="00:04:42.01" />
                    <SPLIT distance="350" swimtime="00:05:32.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-18" firstname="Linda" gender="F" lastname="Spišáková" nation="SVK" license="SVK18707" athleteid="15948">
              <RESULTS>
                <RESULT eventid="1096" points="208" reactiontime="+90" swimtime="00:03:25.58" resultid="15949" heatid="19306" lane="8" entrytime="00:03:39.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.33" />
                    <SPLIT distance="100" swimtime="00:01:43.25" />
                    <SPLIT distance="150" swimtime="00:02:38.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="206" reactiontime="+105" swimtime="00:01:35.91" resultid="15950" heatid="19391" lane="1" entrytime="00:01:37.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="270" reactiontime="+97" swimtime="00:01:36.41" resultid="15951" heatid="19429" lane="4" entrytime="00:01:37.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="130" reactiontime="+85" swimtime="00:00:48.12" resultid="15952" heatid="19446" lane="9" entrytime="00:00:43.70" />
                <RESULT eventid="1664" points="291" reactiontime="+87" swimtime="00:00:43.19" resultid="15953" heatid="19542" lane="8" entrytime="00:00:43.42" />
                <RESULT eventid="1222" points="263" reactiontime="+83" swimtime="00:03:29.83" resultid="17754" heatid="19357" lane="9" entrytime="00:03:32.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.02" />
                    <SPLIT distance="100" swimtime="00:01:41.79" />
                    <SPLIT distance="150" swimtime="00:02:37.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-12-14" firstname="Roman" gender="M" lastname="Kubera" nation="SVK" license="SVK21009" athleteid="15941">
              <RESULTS>
                <RESULT eventid="1079" points="196" reactiontime="+85" swimtime="00:00:34.85" resultid="15942" heatid="19287" lane="4" entrytime="00:00:35.28" />
                <RESULT eventid="1273" points="157" reactiontime="+105" swimtime="00:01:23.19" resultid="15943" heatid="19376" lane="6" entrytime="00:01:25.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="196" reactiontime="+75" swimtime="00:02:35.66" resultid="15969" heatid="19422" lane="0" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                    <SPLIT distance="100" swimtime="00:01:20.97" />
                    <SPLIT distance="150" swimtime="00:02:00.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15922" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="15915" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="15918" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="15934" number="4" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" points="229" reactiontime="+84" swimtime="00:02:14.93" resultid="15970" heatid="19500" lane="9" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                    <SPLIT distance="100" swimtime="00:01:12.93" />
                    <SPLIT distance="150" swimtime="00:01:47.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15918" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="15934" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="15941" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="15922" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1358" points="168" swimtime="00:03:07.10" resultid="15967" heatid="19420" lane="8" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.14" />
                    <SPLIT distance="150" swimtime="00:02:26.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15954" number="1" />
                    <RELAYPOSITION athleteid="15959" number="2" />
                    <RELAYPOSITION athleteid="15929" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="15948" number="4" reactiontime="+7" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1525" points="122" reactiontime="+92" swimtime="00:03:09.99" resultid="15968" heatid="19497" lane="5" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.15" />
                    <SPLIT distance="100" swimtime="00:01:31.98" />
                    <SPLIT distance="150" swimtime="00:02:07.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15948" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="15959" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="15954" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="15944" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="217" reactiontime="+95" swimtime="00:02:27.28" resultid="15965" heatid="19320" lane="2" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                    <SPLIT distance="100" swimtime="00:01:11.61" />
                    <SPLIT distance="150" swimtime="00:01:59.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15941" number="1" reactiontime="+95" />
                    <RELAYPOSITION athleteid="15948" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="15929" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="15922" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="181" reactiontime="+97" swimtime="00:02:51.51" resultid="15966" heatid="19562" lane="1" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.84" />
                    <SPLIT distance="100" swimtime="00:01:34.76" />
                    <SPLIT distance="150" swimtime="00:02:16.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15918" number="1" reactiontime="+97" />
                    <RELAYPOSITION athleteid="15948" number="2" reactiontime="+27" />
                    <RELAYPOSITION athleteid="15954" number="3" reactiontime="+23" />
                    <RELAYPOSITION athleteid="15941" number="4" reactiontime="+5" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1698" points="237" reactiontime="+73" swimtime="00:02:37.01" resultid="15971" heatid="19562" lane="5" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                    <SPLIT distance="100" swimtime="00:01:24.73" />
                    <SPLIT distance="150" swimtime="00:02:02.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15922" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="15929" number="2" reactiontime="+85" />
                    <RELAYPOSITION athleteid="15963" number="3" reactiontime="+30" />
                    <RELAYPOSITION athleteid="15934" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SLPL" nation="CZE" clubid="18412" name="Plavecký klub Slávia VŠ Plzeň">
          <CONTACT email="Vlastimil.Havlicek@seznam.cz" name="Vlastimil Havlicek" phone="+421602892172" />
          <ATHLETES>
            <ATHLETE birthdate="1977-04-29" firstname="Petr" gender="M" lastname="Hejnic" nation="CZE" athleteid="18416">
              <RESULTS>
                <RESULT eventid="1113" points="376" reactiontime="+81" swimtime="00:02:31.82" resultid="18417" heatid="19317" lane="9" entrytime="00:02:28.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.06" />
                    <SPLIT distance="100" swimtime="00:01:12.55" />
                    <SPLIT distance="150" swimtime="00:01:55.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="382" reactiontime="+84" swimtime="00:02:45.94" resultid="18418" heatid="19364" lane="6" entrytime="00:02:44.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.62" />
                    <SPLIT distance="100" swimtime="00:01:20.56" />
                    <SPLIT distance="150" swimtime="00:02:02.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="379" reactiontime="+86" swimtime="00:01:09.48" resultid="18419" heatid="19407" lane="7" entrytime="00:01:08.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="389" reactiontime="+86" swimtime="00:01:16.14" resultid="18420" heatid="19441" lane="7" entrytime="00:01:14.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-08-20" firstname="Vlastimil" gender="M" lastname="Havlíček" nation="CZE" athleteid="18413">
              <RESULTS>
                <RESULT eventid="1079" points="574" reactiontime="+75" swimtime="00:00:24.37" resultid="18414" heatid="19303" lane="4" entrytime="00:00:24.32" />
                <RESULT eventid="1440" points="580" reactiontime="+71" swimtime="00:00:26.14" resultid="18415" heatid="19464" lane="9" entrytime="00:00:26.28" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="CZE" clubid="18525" name="Plavecký klub Zábřeh">
          <CONTACT city="Zábřeh na Moravě" email="sipjir73@seznam.cz" name="Jiří Šíp" state="CZE" />
          <ATHLETES>
            <ATHLETE birthdate="1973-09-19" firstname="Jiří" gender="M" lastname="Šíp" nation="CZE" athleteid="18526">
              <RESULTS>
                <RESULT eventid="1113" points="371" reactiontime="+86" swimtime="00:02:32.46" resultid="18527" heatid="19315" lane="8" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                    <SPLIT distance="100" swimtime="00:01:11.95" />
                    <SPLIT distance="150" swimtime="00:01:58.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="328" reactiontime="+83" swimtime="00:00:32.21" resultid="18528" heatid="19350" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="14243" points="416" reactiontime="+89" swimtime="00:01:07.37" resultid="18529" heatid="19406" lane="4" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="359" reactiontime="+82" swimtime="00:01:08.77" resultid="18530" heatid="19476" lane="5" entrytime="00:01:10.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O4 - Start wykonany przed sygnłem (przedwczesny start) (Time: 10:32)" eventid="1647" reactiontime="+61" status="DSQ" swimtime="00:02:37.33" resultid="18531" heatid="19536" lane="9" entrytime="00:02:41.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                    <SPLIT distance="100" swimtime="00:01:15.10" />
                    <SPLIT distance="150" swimtime="00:01:56.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="RUS" clubid="16122" name="Pregel">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1965-01-01" firstname="Vadim" gender="M" lastname="Ezhkov" nation="RUS" athleteid="16123">
              <RESULTS>
                <RESULT eventid="1079" points="291" reactiontime="+67" swimtime="00:00:30.54" resultid="16124" heatid="19292" lane="8" entrytime="00:00:30.50" />
                <RESULT eventid="1113" points="260" reactiontime="+68" swimtime="00:02:51.68" resultid="16125" heatid="19313" lane="9" entrytime="00:02:53.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.97" />
                    <SPLIT distance="100" swimtime="00:01:21.89" />
                    <SPLIT distance="150" swimtime="00:02:09.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="302" reactiontime="+75" swimtime="00:01:06.95" resultid="16126" heatid="19380" lane="1" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="293" reactiontime="+76" swimtime="00:01:15.70" resultid="16127" heatid="19403" lane="1" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="319" reactiontime="+73" swimtime="00:01:21.35" resultid="16128" heatid="19438" lane="5" entrytime="00:01:24.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="196" reactiontime="+78" swimtime="00:01:24.11" resultid="16129" heatid="19473" lane="5" entrytime="00:01:27.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="338" reactiontime="+72" swimtime="00:00:36.24" resultid="16130" heatid="19553" lane="6" entrytime="00:00:37.50" />
                <RESULT eventid="1744" points="280" reactiontime="+74" swimtime="00:05:24.25" resultid="16131" heatid="19704" lane="1" entrytime="00:05:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                    <SPLIT distance="100" swimtime="00:01:15.79" />
                    <SPLIT distance="150" swimtime="00:01:56.67" />
                    <SPLIT distance="200" swimtime="00:02:38.24" />
                    <SPLIT distance="250" swimtime="00:03:19.58" />
                    <SPLIT distance="300" swimtime="00:04:01.93" />
                    <SPLIT distance="350" swimtime="00:04:43.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Aleksandr" gender="M" lastname="Smirnov" nation="RUS" athleteid="16132">
              <RESULTS>
                <RESULT eventid="14207" points="389" reactiontime="+96" swimtime="00:19:21.01" resultid="16133" heatid="19623" lane="7" entrytime="00:19:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                    <SPLIT distance="200" swimtime="00:02:27.72" />
                    <SPLIT distance="250" swimtime="00:03:05.47" />
                    <SPLIT distance="300" swimtime="00:03:43.42" />
                    <SPLIT distance="350" swimtime="00:04:21.74" />
                    <SPLIT distance="400" swimtime="00:05:00.17" />
                    <SPLIT distance="450" swimtime="00:05:38.54" />
                    <SPLIT distance="500" swimtime="00:06:17.02" />
                    <SPLIT distance="550" swimtime="00:06:55.68" />
                    <SPLIT distance="600" swimtime="00:07:34.71" />
                    <SPLIT distance="650" swimtime="00:08:13.55" />
                    <SPLIT distance="700" swimtime="00:08:53.10" />
                    <SPLIT distance="750" swimtime="00:09:32.20" />
                    <SPLIT distance="800" swimtime="00:10:11.47" />
                    <SPLIT distance="850" swimtime="00:10:50.53" />
                    <SPLIT distance="900" swimtime="00:11:29.79" />
                    <SPLIT distance="950" swimtime="00:12:09.35" />
                    <SPLIT distance="1000" swimtime="00:12:48.63" />
                    <SPLIT distance="1050" swimtime="00:13:28.28" />
                    <SPLIT distance="1100" swimtime="00:14:07.95" />
                    <SPLIT distance="1150" swimtime="00:14:47.57" />
                    <SPLIT distance="1200" swimtime="00:15:27.12" />
                    <SPLIT distance="1250" swimtime="00:16:06.65" />
                    <SPLIT distance="1300" swimtime="00:16:46.53" />
                    <SPLIT distance="1350" swimtime="00:17:25.95" />
                    <SPLIT distance="1400" swimtime="00:18:05.16" />
                    <SPLIT distance="1450" swimtime="00:18:44.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="16134" heatid="19493" lane="1" entrytime="00:02:19.50" />
                <RESULT eventid="1744" points="398" reactiontime="+98" swimtime="00:04:48.51" resultid="16135" heatid="19706" lane="6" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                    <SPLIT distance="100" swimtime="00:01:08.87" />
                    <SPLIT distance="150" swimtime="00:01:45.89" />
                    <SPLIT distance="200" swimtime="00:02:22.67" />
                    <SPLIT distance="250" swimtime="00:02:59.91" />
                    <SPLIT distance="300" swimtime="00:03:36.96" />
                    <SPLIT distance="350" swimtime="00:04:13.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="617" nation="CZE" clubid="14539" name="PVK Brno">
          <CONTACT name="Mr. Smerda" street="Velkopavlovicka" zip="60200" />
          <ATHLETES>
            <ATHLETE birthdate="1979-02-05" firstname="Michal" gender="M" lastname="Fiala" nation="CZE" athleteid="14552">
              <RESULTS>
                <RESULT eventid="1239" points="239" reactiontime="+96" swimtime="00:03:14.05" resultid="14553" heatid="19362" lane="7" entrytime="00:03:11.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.31" />
                    <SPLIT distance="100" swimtime="00:01:33.74" />
                    <SPLIT distance="150" swimtime="00:02:25.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="219" reactiontime="+90" swimtime="00:01:23.34" resultid="14554" heatid="19402" lane="9" entrytime="00:01:20.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="233" reactiontime="+88" swimtime="00:01:30.28" resultid="14555" heatid="19438" lane="0" entrytime="00:01:27.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="257" reactiontime="+93" swimtime="00:02:36.20" resultid="14556" heatid="19490" lane="5" entrytime="00:02:38.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                    <SPLIT distance="100" swimtime="00:01:15.48" />
                    <SPLIT distance="150" swimtime="00:01:57.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="188" reactiontime="+89" swimtime="00:01:23.81" resultid="14557" heatid="19520" lane="8" entrytime="00:01:19.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O4 - Start wykonany przed sygnłem (przedwczesny start) (Time: 11:13)" eventid="1681" status="DSQ" swimtime="00:00:00.00" resultid="14558" heatid="19553" lane="9" entrytime="00:00:38.88" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1941-12-06" firstname="Frantisek" gender="M" lastname="Pokorny" nation="CZE" athleteid="14559">
              <RESULTS>
                <RESULT eventid="14243" points="182" reactiontime="+97" swimtime="00:01:28.62" resultid="14560" heatid="19400" lane="3" entrytime="00:01:28.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="232" reactiontime="+99" swimtime="00:00:35.46" resultid="14561" heatid="19454" lane="1" entrytime="00:00:35.58" />
                <RESULT eventid="1681" points="214" reactiontime="+96" swimtime="00:00:42.19" resultid="14562" heatid="19550" lane="5" entrytime="00:00:42.49" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-03-05" firstname="Michaela" gender="F" lastname="Konecna" nation="CZE" athleteid="14570">
              <RESULTS>
                <RESULT eventid="1256" points="297" reactiontime="+94" swimtime="00:01:16.27" resultid="14571" heatid="19370" lane="2" entrytime="00:01:15.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="278" reactiontime="+90" swimtime="00:01:26.83" resultid="14572" heatid="19392" lane="4" entrytime="00:01:26.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="220" reactiontime="+141" swimtime="00:00:40.36" resultid="14573" heatid="19447" lane="9" entrytime="00:00:38.05" />
                <RESULT eventid="1491" points="267" reactiontime="+81" swimtime="00:02:51.86" resultid="14574" heatid="19482" lane="9" entrytime="00:03:01.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.65" />
                    <SPLIT distance="100" swimtime="00:01:21.97" />
                    <SPLIT distance="150" swimtime="00:02:07.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="235" reactiontime="+83" swimtime="00:01:28.46" resultid="14575" heatid="19514" lane="8" entrytime="00:01:28.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-12" firstname="Jaroslava" gender="F" lastname="Stritezska" nation="CZE" athleteid="14576">
              <RESULTS>
                <RESULT eventid="1187" points="101" reactiontime="+78" swimtime="00:00:55.07" resultid="14577" heatid="19337" lane="0" entrytime="00:00:54.23" />
                <RESULT eventid="14225" points="108" reactiontime="+96" swimtime="00:01:58.70" resultid="14578" heatid="19390" lane="8" entrytime="00:02:03.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="140" reactiontime="+117" swimtime="00:01:59.94" resultid="14579" heatid="19428" lane="0" entrytime="00:02:04.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="156" reactiontime="+130" swimtime="00:00:53.12" resultid="14580" heatid="19540" lane="1" entrytime="00:00:53.11" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-02-15" firstname="Rudolf" gender="M" lastname="Smerda" nation="CZE" athleteid="14563">
              <RESULTS>
                <RESULT eventid="1273" points="259" reactiontime="+88" swimtime="00:01:10.46" resultid="14564" heatid="19379" lane="8" entrytime="00:01:12.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="188" reactiontime="+96" swimtime="00:03:09.45" resultid="14565" heatid="19415" lane="2" entrytime="00:03:18.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="266" reactiontime="+84" swimtime="00:00:33.87" resultid="14566" heatid="19455" lane="7" entrytime="00:00:34.11" />
                <RESULT eventid="1508" points="252" reactiontime="+94" swimtime="00:02:37.21" resultid="14567" heatid="19489" lane="4" entrytime="00:02:47.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.83" />
                    <SPLIT distance="100" swimtime="00:01:18.18" />
                    <SPLIT distance="150" swimtime="00:02:00.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="193" reactiontime="+82" swimtime="00:01:23.12" resultid="14568" heatid="19520" lane="9" entrytime="00:01:23.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="14569" heatid="19703" lane="1" entrytime="00:05:57.33" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="RMKS" nation="POL" region="SLA" clubid="14581" name="RMKS Rybnik">
          <CONTACT city="Rybnik" email="aniaduda0511@tlen.pl" name="DUDA ANNA" phone="792666159" state="SLA" street="orzepowicka 22a/37" zip="44-217" />
          <ATHLETES>
            <ATHLETE birthdate="1981-04-15" firstname="Anna" gender="F" lastname="Duda" nation="POL" athleteid="14587">
              <RESULTS>
                <RESULT eventid="1062" points="603" reactiontime="+83" swimtime="00:00:27.50" resultid="14588" heatid="19283" lane="6" entrytime="00:00:27.80" />
                <RESULT eventid="1096" points="447" reactiontime="+90" swimtime="00:02:39.29" resultid="14589" heatid="19309" lane="1" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                    <SPLIT distance="100" swimtime="00:01:16.52" />
                    <SPLIT distance="150" swimtime="00:02:02.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="542" reactiontime="+85" swimtime="00:01:02.43" resultid="14590" heatid="19372" lane="1" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="477" reactiontime="+86" swimtime="00:01:12.48" resultid="14591" heatid="19396" lane="0" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1423" points="585" reactiontime="+78" swimtime="00:00:29.14" resultid="14592" heatid="19449" lane="5" entrytime="00:00:29.90" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1555" points="414" reactiontime="+100" swimtime="00:05:48.01" resultid="14593" heatid="19505" lane="1" entrytime="00:05:50.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.31" />
                    <SPLIT distance="150" swimtime="00:02:05.83" />
                    <SPLIT distance="200" swimtime="00:02:51.91" />
                    <SPLIT distance="250" swimtime="00:03:43.22" />
                    <SPLIT distance="300" swimtime="00:04:33.74" />
                    <SPLIT distance="350" swimtime="00:05:12.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="512" reactiontime="+83" swimtime="00:01:08.22" resultid="14594" heatid="19515" lane="5" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="452" reactiontime="+82" swimtime="00:00:37.31" resultid="14595" heatid="19544" lane="6" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-03" firstname="Agnieszka" gender="F" lastname="Bieniak" nation="POL" athleteid="14582">
              <RESULTS>
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="14583" heatid="19341" lane="9" entrytime="00:00:34.00" />
                <RESULT eventid="1388" status="DNS" swimtime="00:00:00.00" resultid="14584" heatid="19432" lane="8" entrytime="00:01:23.00" />
                <RESULT eventid="1457" status="DNS" swimtime="00:00:00.00" resultid="14585" heatid="19469" lane="8" entrytime="00:01:12.00" />
                <RESULT eventid="1630" points="416" reactiontime="+71" swimtime="00:02:39.66" resultid="14586" heatid="19529" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                    <SPLIT distance="100" swimtime="00:01:14.23" />
                    <SPLIT distance="150" swimtime="00:01:55.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="14303" name="Rydułtoeska Akademia Aktywnego Seniora" shortname="Rydułtoeska Akademia Aktywnego">
          <CONTACT email="otelom.090866@interia.pl" name="Otlik Marian" />
          <ATHLETES>
            <ATHLETE birthdate="1946-02-02" firstname="Lippa" gender="F" lastname="Maria" nation="POL" athleteid="14402">
              <RESULTS>
                <RESULT eventid="1147" reactiontime="+152" status="OTL" swimtime="00:23:04.35" resultid="14403" heatid="19594" lane="3" entrytime="00:23:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.60" />
                    <SPLIT distance="100" swimtime="00:02:36.39" />
                    <SPLIT distance="150" swimtime="00:04:04.43" />
                    <SPLIT distance="200" swimtime="00:05:33.72" />
                    <SPLIT distance="250" swimtime="00:07:01.45" />
                    <SPLIT distance="300" swimtime="00:08:30.29" />
                    <SPLIT distance="350" swimtime="00:09:58.11" />
                    <SPLIT distance="400" swimtime="00:11:25.51" />
                    <SPLIT distance="450" swimtime="00:12:51.99" />
                    <SPLIT distance="500" swimtime="00:14:20.37" />
                    <SPLIT distance="550" swimtime="00:15:47.34" />
                    <SPLIT distance="600" swimtime="00:17:15.12" />
                    <SPLIT distance="650" swimtime="00:18:42.46" />
                    <SPLIT distance="750" swimtime="00:21:37.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="29" reactiontime="+190" swimtime="00:01:22.89" resultid="14404" heatid="19336" lane="1" />
                <RESULT eventid="1256" points="28" reactiontime="+122" swimtime="00:02:47.12" resultid="14405" heatid="19367" lane="7" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="29" reactiontime="+97" swimtime="00:02:57.46" resultid="14406" heatid="19465" lane="3" entrytime="00:03:06.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:25.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="37" reactiontime="+133" swimtime="00:05:29.95" resultid="14407" heatid="19479" lane="4" entrytime="00:05:21.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.64" />
                    <SPLIT distance="100" swimtime="00:02:36.75" />
                    <SPLIT distance="150" swimtime="00:04:04.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="34" reactiontime="+138" swimtime="00:06:07.74" resultid="14408" heatid="19526" lane="1" entrytime="00:06:32.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.77" />
                    <SPLIT distance="100" swimtime="00:02:57.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="44" reactiontime="+133" swimtime="00:11:01.83" resultid="14409" heatid="19695" lane="0" entrytime="00:10:45.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.52" />
                    <SPLIT distance="100" swimtime="00:02:35.04" />
                    <SPLIT distance="150" swimtime="00:03:57.64" />
                    <SPLIT distance="200" swimtime="00:05:22.59" />
                    <SPLIT distance="250" swimtime="00:06:47.86" />
                    <SPLIT distance="300" swimtime="00:08:12.93" />
                    <SPLIT distance="350" swimtime="00:09:37.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1945-12-07" firstname="Miron" gender="M" lastname="Starosta" nation="POL" athleteid="14410">
              <RESULTS>
                <RESULT eventid="1079" points="74" reactiontime="+147" swimtime="00:00:48.05" resultid="14411" heatid="19284" lane="0" />
                <RESULT eventid="1113" points="58" reactiontime="+153" swimtime="00:04:42.53" resultid="14412" heatid="19310" lane="0" entrytime="00:04:46.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.41" />
                    <SPLIT distance="100" swimtime="00:02:17.98" />
                    <SPLIT distance="150" swimtime="00:03:40.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="66" reactiontime="+106" swimtime="00:04:57.67" resultid="14413" heatid="19359" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.01" />
                    <SPLIT distance="100" swimtime="00:02:24.26" />
                    <SPLIT distance="150" swimtime="00:03:42.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="60" reactiontime="+87" swimtime="00:02:08.48" resultid="14414" heatid="19397" lane="4" entrytime="00:02:12.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="65" swimtime="00:02:18.00" resultid="14415" heatid="19434" lane="0" entrytime="00:02:24.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" reactiontime="+99" status="DNF" swimtime="00:09:18.14" resultid="14416" heatid="19507" lane="8" entrytime="00:10:47.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.81" />
                    <SPLIT distance="100" swimtime="00:02:44.94" />
                    <SPLIT distance="150" swimtime="00:04:08.87" />
                    <SPLIT distance="200" swimtime="00:05:31.19" />
                    <SPLIT distance="250" swimtime="00:06:58.60" />
                    <SPLIT distance="350" swimtime="00:08:07.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="44" reactiontime="+103" swimtime="00:04:57.00" resultid="14417" heatid="19530" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.63" />
                    <SPLIT distance="100" swimtime="00:02:15.06" />
                    <SPLIT distance="150" swimtime="00:03:38.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="71" reactiontime="+92" swimtime="00:01:00.73" resultid="14418" heatid="19546" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-11-24" firstname="Jerzy" gender="M" lastname="Ciecior" nation="POL" athleteid="14393">
              <RESULTS>
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="14394" heatid="19318" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="14207" points="191" reactiontime="+90" swimtime="00:24:30.60" resultid="14395" heatid="19620" lane="4" entrytime="00:25:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.50" />
                    <SPLIT distance="100" swimtime="00:01:29.42" />
                    <SPLIT distance="150" swimtime="00:02:17.54" />
                    <SPLIT distance="200" swimtime="00:03:05.88" />
                    <SPLIT distance="250" swimtime="00:03:54.74" />
                    <SPLIT distance="300" swimtime="00:04:43.80" />
                    <SPLIT distance="350" swimtime="00:05:33.20" />
                    <SPLIT distance="400" swimtime="00:06:22.54" />
                    <SPLIT distance="450" swimtime="00:07:11.83" />
                    <SPLIT distance="500" swimtime="00:08:01.26" />
                    <SPLIT distance="550" swimtime="00:08:50.53" />
                    <SPLIT distance="600" swimtime="00:09:40.19" />
                    <SPLIT distance="650" swimtime="00:10:30.01" />
                    <SPLIT distance="700" swimtime="00:11:19.93" />
                    <SPLIT distance="750" swimtime="00:12:10.14" />
                    <SPLIT distance="800" swimtime="00:13:00.09" />
                    <SPLIT distance="850" swimtime="00:13:50.04" />
                    <SPLIT distance="900" swimtime="00:14:39.38" />
                    <SPLIT distance="950" swimtime="00:15:28.85" />
                    <SPLIT distance="1000" swimtime="00:16:18.40" />
                    <SPLIT distance="1050" swimtime="00:17:08.00" />
                    <SPLIT distance="1100" swimtime="00:17:57.66" />
                    <SPLIT distance="1150" swimtime="00:18:47.09" />
                    <SPLIT distance="1200" swimtime="00:19:36.88" />
                    <SPLIT distance="1250" swimtime="00:20:26.30" />
                    <SPLIT distance="1300" swimtime="00:21:16.18" />
                    <SPLIT distance="1350" swimtime="00:22:05.47" />
                    <SPLIT distance="1400" swimtime="00:22:55.14" />
                    <SPLIT distance="1450" swimtime="00:23:43.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="170" swimtime="00:00:40.08" resultid="14396" heatid="19346" lane="8" entrytime="00:00:42.00" />
                <RESULT eventid="1341" points="99" reactiontime="+94" swimtime="00:03:54.04" resultid="14397" heatid="19415" lane="0" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.84" />
                    <SPLIT distance="100" swimtime="00:01:47.93" />
                    <SPLIT distance="150" swimtime="00:02:52.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="157" reactiontime="+82" swimtime="00:01:30.61" resultid="14398" heatid="19473" lane="1" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="14399" heatid="19508" lane="1" entrytime="00:07:15.00" />
                <RESULT eventid="1613" points="140" reactiontime="+73" swimtime="00:01:32.53" resultid="14400" heatid="19519" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="146" reactiontime="+91" swimtime="00:03:20.17" resultid="14401" heatid="19533" lane="5" entrytime="00:03:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.99" />
                    <SPLIT distance="100" swimtime="00:01:37.15" />
                    <SPLIT distance="150" swimtime="00:02:30.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-05-26" firstname="Władysław" gender="M" lastname="Szurek" nation="POL" athleteid="14386">
              <RESULTS>
                <RESULT eventid="1205" points="14" reactiontime="+120" swimtime="00:01:30.83" resultid="14387" heatid="19342" lane="3" entrytime="00:01:29.00" />
                <RESULT eventid="1273" points="23" reactiontime="+119" swimtime="00:02:37.60" resultid="14388" heatid="19374" lane="8" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="13" reactiontime="+99" swimtime="00:03:25.99" resultid="14389" heatid="19470" lane="6" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:35.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="22" reactiontime="+118" swimtime="00:05:50.84" resultid="14390" heatid="19486" lane="1" entrytime="00:05:30.00" />
                <RESULT eventid="1647" points="14" reactiontime="+98" swimtime="00:07:12.70" resultid="14391" heatid="19531" lane="1" entrytime="00:07:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:35.43" />
                    <SPLIT distance="100" swimtime="00:03:26.23" />
                    <SPLIT distance="150" swimtime="00:05:20.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="25" reactiontime="+116" swimtime="00:12:03.01" resultid="14392" heatid="19699" lane="6" entrytime="00:11:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.02" />
                    <SPLIT distance="100" swimtime="00:02:39.37" />
                    <SPLIT distance="200" swimtime="00:05:43.24" />
                    <SPLIT distance="250" swimtime="00:07:17.69" />
                    <SPLIT distance="300" swimtime="00:08:52.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-05-16" firstname="Rudolf" gender="M" lastname="Bugla" nation="POL" athleteid="14377">
              <RESULTS>
                <RESULT eventid="1079" points="67" reactiontime="+110" swimtime="00:00:49.86" resultid="14378" heatid="19285" lane="8" entrytime="00:00:45.00" />
                <RESULT eventid="1113" points="60" reactiontime="+114" swimtime="00:04:39.04" resultid="14379" heatid="19310" lane="1" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.03" />
                    <SPLIT distance="100" swimtime="00:02:17.23" />
                    <SPLIT distance="150" swimtime="00:03:36.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="46" reactiontime="+87" swimtime="00:01:01.59" resultid="14380" heatid="19343" lane="4" entrytime="00:00:55.30" />
                <RESULT eventid="1341" points="32" reactiontime="+102" swimtime="00:05:38.94" resultid="14381" heatid="19414" lane="8" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.46" />
                    <SPLIT distance="100" swimtime="00:02:38.17" />
                    <SPLIT distance="150" swimtime="00:04:07.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="42" reactiontime="+112" swimtime="00:01:02.40" resultid="14382" heatid="19451" lane="8" entrytime="00:00:59.50" />
                <RESULT eventid="1578" points="51" reactiontime="+108" swimtime="00:10:34.56" resultid="14383" heatid="19507" lane="1" entrytime="00:09:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.97" />
                    <SPLIT distance="100" swimtime="00:02:44.17" />
                    <SPLIT distance="150" swimtime="00:05:29.09" />
                    <SPLIT distance="200" swimtime="00:06:52.00" />
                    <SPLIT distance="250" swimtime="00:08:14.09" />
                    <SPLIT distance="350" swimtime="00:09:25.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="36" reactiontime="+102" swimtime="00:02:24.78" resultid="14384" heatid="19517" lane="1" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="45" reactiontime="+89" swimtime="00:04:56.43" resultid="14385" heatid="19532" lane="0" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.43" />
                    <SPLIT distance="100" swimtime="00:02:24.72" />
                    <SPLIT distance="150" swimtime="00:03:42.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-08-21" firstname="Michał" gender="M" lastname="Kądzioła" nation="POL" athleteid="14419">
              <RESULTS>
                <RESULT eventid="1079" points="370" reactiontime="+84" swimtime="00:00:28.22" resultid="14420" heatid="19294" lane="1" entrytime="00:00:29.50" />
                <RESULT eventid="1113" points="252" reactiontime="+95" swimtime="00:02:53.50" resultid="14421" heatid="19313" lane="0" entrytime="00:02:52.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                    <SPLIT distance="100" swimtime="00:01:15.58" />
                    <SPLIT distance="150" swimtime="00:02:09.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="307" reactiontime="+77" swimtime="00:00:32.93" resultid="14422" heatid="19349" lane="3" entrytime="00:00:33.11" />
                <RESULT eventid="14243" points="310" reactiontime="+87" swimtime="00:01:14.31" resultid="14423" heatid="19404" lane="3" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="342" reactiontime="+77" swimtime="00:00:31.16" resultid="14424" heatid="19459" lane="9" entrytime="00:00:30.88" />
                <RESULT eventid="1474" points="282" reactiontime="+84" swimtime="00:01:14.58" resultid="14425" heatid="19475" lane="4" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="14426" heatid="19509" lane="2" entrytime="00:06:15.00" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="14427" heatid="19521" lane="8" entrytime="00:01:14.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="17523" name="SBC">
          <CONTACT email="blochmaciek8@gmail.com" name="Bloch" phone="668800005" />
          <ATHLETES>
            <ATHLETE birthdate="1972-03-11" firstname="Dorota" gender="F" lastname="Batóg" nation="POL" athleteid="17555">
              <RESULTS>
                <RESULT eventid="1062" points="340" reactiontime="+91" swimtime="00:00:33.29" resultid="17556" heatid="19279" lane="4" entrytime="00:00:34.34" />
                <RESULT eventid="1187" points="240" reactiontime="+112" swimtime="00:00:41.26" resultid="17557" heatid="19338" lane="3" entrytime="00:00:41.73" />
                <RESULT eventid="1256" points="305" reactiontime="+85" swimtime="00:01:15.57" resultid="17558" heatid="19370" lane="9" entrytime="00:01:19.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="292" reactiontime="+82" swimtime="00:01:25.35" resultid="17559" heatid="19392" lane="8" entrytime="00:01:29.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="237" reactiontime="+87" swimtime="00:00:39.37" resultid="17560" heatid="19446" lane="6" entrytime="00:00:39.35" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-05-11" firstname="Joanna" gender="F" lastname="Krowicka" nation="POL" athleteid="17547">
              <RESULTS>
                <RESULT eventid="1062" points="232" reactiontime="+81" swimtime="00:00:37.82" resultid="17548" heatid="19278" lane="7" entrytime="00:00:38.90" />
                <RESULT eventid="1096" points="169" reactiontime="+72" swimtime="00:03:40.13" resultid="17549" heatid="19306" lane="9" entrytime="00:03:50.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.35" />
                    <SPLIT distance="100" swimtime="00:01:53.22" />
                    <SPLIT distance="150" swimtime="00:02:51.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="219" reactiontime="+87" swimtime="00:03:43.19" resultid="17550" heatid="19356" lane="3" entrytime="00:03:41.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.50" />
                    <SPLIT distance="100" swimtime="00:01:47.69" />
                    <SPLIT distance="150" swimtime="00:02:46.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="200" reactiontime="+82" swimtime="00:01:36.81" resultid="17551" heatid="19391" lane="8" entrytime="00:01:39.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="221" reactiontime="+83" swimtime="00:01:43.14" resultid="17552" heatid="19429" lane="7" entrytime="00:01:41.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="117" reactiontime="+87" swimtime="00:00:49.81" resultid="17553" heatid="19445" lane="6" entrytime="00:00:49.19" />
                <RESULT eventid="1664" points="248" reactiontime="+71" swimtime="00:00:45.56" resultid="17554" heatid="19541" lane="6" entrytime="00:00:45.72" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-07" firstname="Radosław" gender="M" lastname="Stefurak" nation="POL" athleteid="17542">
              <RESULTS>
                <RESULT eventid="1239" points="266" reactiontime="+84" swimtime="00:03:07.13" resultid="17543" heatid="19363" lane="9" entrytime="00:03:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                    <SPLIT distance="100" swimtime="00:01:26.45" />
                    <SPLIT distance="150" swimtime="00:02:16.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="267" reactiontime="+106" swimtime="00:01:26.36" resultid="17544" heatid="19438" lane="4" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="223" reactiontime="+87" swimtime="00:02:43.63" resultid="17545" heatid="19490" lane="6" entrytime="00:02:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.10" />
                    <SPLIT distance="100" swimtime="00:01:16.80" />
                    <SPLIT distance="150" swimtime="00:02:00.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="17546" heatid="19554" lane="9" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DIA" nation="AUT" region="WLSV" clubid="14753" name="SC Diana" shortname="Diana">
          <ATHLETES>
            <ATHLETE birthdate="1985-07-16" firstname="Agata" gender="F" lastname="Wycisk" nation="POL" license="44612" athleteid="14754">
              <RESULTS>
                <RESULT eventid="1062" points="101" reactiontime="+89" swimtime="00:00:49.78" resultid="14755" heatid="19276" lane="6" entrytime="00:00:49.66" />
                <RESULT eventid="1222" points="191" reactiontime="+100" swimtime="00:03:53.61" resultid="14756" heatid="19354" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.43" />
                    <SPLIT distance="100" swimtime="00:01:54.30" />
                    <SPLIT distance="150" swimtime="00:02:54.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="103" swimtime="00:01:48.59" resultid="14757" heatid="19368" lane="0" entrytime="00:01:46.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="172" reactiontime="+95" swimtime="00:01:52.07" resultid="14758" heatid="19428" lane="3" entrytime="00:01:52.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="106" reactiontime="+89" swimtime="00:03:53.45" resultid="14759" heatid="19480" lane="7" entrytime="00:03:52.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.96" />
                    <SPLIT distance="100" swimtime="00:01:52.95" />
                    <SPLIT distance="150" swimtime="00:02:54.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" status="DNS" swimtime="00:00:00.00" resultid="14760" heatid="19540" lane="8" entrytime="00:00:53.43" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="14295" name="SG Erkelenz - Hückelhoven">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1967-01-29" firstname="Dariusz" gender="M" lastname="Andrzejczak" nation="GER" athleteid="14296">
              <RESULTS>
                <RESULT eventid="1079" points="489" swimtime="00:00:25.70" resultid="14297" heatid="19301" lane="0" entrytime="00:00:26.00" />
                <RESULT eventid="1205" points="342" reactiontime="+60" swimtime="00:00:31.77" resultid="14298" heatid="19351" lane="9" entrytime="00:00:31.00" />
                <RESULT eventid="14243" points="388" reactiontime="+76" swimtime="00:01:08.91" resultid="14299" heatid="19408" lane="8" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="436" reactiontime="+80" swimtime="00:00:28.74" resultid="14300" heatid="19461" lane="4" entrytime="00:00:28.00" />
                <RESULT eventid="1613" points="363" reactiontime="+85" swimtime="00:01:07.37" resultid="14301" heatid="19524" lane="4" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="414" reactiontime="+86" swimtime="00:00:33.86" resultid="14302" heatid="19557" lane="5" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="16145" name="SiKReT Gliwice">
          <CONTACT city="GLIWICE" email="joannaeco@tlen.pl" name="JOANNA ZAGAŁA" phone="601427257" state="ŚLĄSK" street="JAGIELOŃSKA 21" zip="44-100" />
          <ATHLETES>
            <ATHLETE birthdate="1959-06-24" firstname="Joanna" gender="F" lastname="Zagała" nation="POL" athleteid="16146">
              <RESULTS>
                <RESULT eventid="1062" points="240" reactiontime="+78" swimtime="00:00:37.35" resultid="16147" heatid="19278" lane="8" entrytime="00:00:39.00" />
                <RESULT eventid="1165" points="193" reactiontime="+98" swimtime="00:26:28.79" resultid="16148" heatid="19624" lane="1" entrytime="00:30:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.07" />
                    <SPLIT distance="100" swimtime="00:02:32.73" />
                    <SPLIT distance="150" swimtime="00:04:20.24" />
                    <SPLIT distance="200" swimtime="00:05:14.29" />
                    <SPLIT distance="250" swimtime="00:06:07.74" />
                    <SPLIT distance="300" swimtime="00:07:55.98" />
                    <SPLIT distance="350" swimtime="00:16:50.92" />
                    <SPLIT distance="400" swimtime="00:19:31.60" />
                    <SPLIT distance="450" swimtime="00:21:18.56" />
                    <SPLIT distance="500" swimtime="00:23:04.74" />
                    <SPLIT distance="850" swimtime="00:23:57.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="156" reactiontime="+78" swimtime="00:00:47.66" resultid="16149" heatid="19337" lane="6" entrytime="00:00:50.00" />
                <RESULT eventid="14225" points="183" reactiontime="+81" swimtime="00:01:39.69" resultid="16150" heatid="19390" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" status="DNS" swimtime="00:00:00.00" resultid="16151" heatid="19466" lane="9" entrytime="00:02:00.00" />
                <RESULT eventid="1491" points="208" reactiontime="+84" swimtime="00:03:06.89" resultid="16152" heatid="19481" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.89" />
                    <SPLIT distance="100" swimtime="00:01:31.36" />
                    <SPLIT distance="150" swimtime="00:02:18.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="146" reactiontime="+91" swimtime="00:03:46.12" resultid="16153" heatid="19527" lane="0" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.49" />
                    <SPLIT distance="100" swimtime="00:01:52.84" />
                    <SPLIT distance="150" swimtime="00:02:51.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="195" reactiontime="+84" swimtime="00:00:49.38" resultid="16154" heatid="19539" lane="3" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-04-20" firstname="Wojciech" gender="M" lastname="Kosiak" nation="POL" athleteid="16176">
              <RESULTS>
                <RESULT eventid="1079" points="117" reactiontime="+116" swimtime="00:00:41.38" resultid="16177" heatid="19285" lane="2" entrytime="00:00:43.00" />
                <RESULT eventid="1273" points="95" reactiontime="+106" swimtime="00:01:38.46" resultid="16178" heatid="19375" lane="7" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="77" reactiontime="+120" swimtime="00:00:51.22" resultid="16179" heatid="19451" lane="9" entrytime="00:01:00.00" />
                <RESULT eventid="1508" points="82" reactiontime="+116" swimtime="00:03:48.04" resultid="16180" heatid="19486" lane="4" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.33" />
                    <SPLIT distance="100" swimtime="00:01:50.12" />
                    <SPLIT distance="150" swimtime="00:02:49.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-03-28" firstname="Łukasz" gender="M" lastname="Stolarczyk" nation="POL" athleteid="16202">
              <RESULTS>
                <RESULT eventid="1273" points="511" reactiontime="+77" swimtime="00:00:56.18" resultid="16203" heatid="19388" lane="9" entrytime="00:00:55.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="491" reactiontime="+84" swimtime="00:00:27.63" resultid="16204" heatid="19462" lane="4" entrytime="00:00:27.15" />
                <RESULT eventid="1613" points="481" reactiontime="+85" swimtime="00:01:01.34" resultid="16205" heatid="19525" lane="1" entrytime="00:01:00.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-02-14" firstname="Dawid" gender="M" lastname="Zimkowski" nation="POL" athleteid="16189">
              <RESULTS>
                <RESULT eventid="1079" points="233" reactiontime="+86" swimtime="00:00:32.90" resultid="16190" heatid="19293" lane="8" entrytime="00:00:30.00" />
                <RESULT eventid="1205" points="247" reactiontime="+68" swimtime="00:00:35.37" resultid="16191" heatid="19348" lane="8" entrytime="00:00:36.00" />
                <RESULT eventid="14243" points="290" reactiontime="+82" swimtime="00:01:15.98" resultid="16192" heatid="19402" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="354" reactiontime="+83" swimtime="00:00:30.80" resultid="16193" heatid="19457" lane="2" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-16" firstname="Stanisław" gender="M" lastname="Twardysko" nation="POL" athleteid="16181">
              <RESULTS>
                <RESULT eventid="1079" points="199" reactiontime="+81" swimtime="00:00:34.68" resultid="16182" heatid="19288" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1205" points="142" reactiontime="+87" swimtime="00:00:42.55" resultid="16183" heatid="19345" lane="2" entrytime="00:00:44.00" />
                <RESULT eventid="1273" points="195" reactiontime="+97" swimtime="00:01:17.45" resultid="16184" heatid="19377" lane="4" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="131" reactiontime="+67" swimtime="00:01:36.24" resultid="16185" heatid="19472" lane="4" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.93" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O4 - Start wykonany przed sygnłem (przedwczesny start) (Time: 18:56)" eventid="1508" reactiontime="+77" status="DSQ" swimtime="00:02:54.64" resultid="16186" heatid="19488" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.33" />
                    <SPLIT distance="100" swimtime="00:01:21.21" />
                    <SPLIT distance="150" swimtime="00:02:08.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="16187" heatid="19533" lane="8" entrytime="00:03:40.00" />
                <RESULT eventid="1744" points="171" reactiontime="+92" swimtime="00:06:22.21" resultid="16188" heatid="19702" lane="8" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.02" />
                    <SPLIT distance="100" swimtime="00:01:23.70" />
                    <SPLIT distance="150" swimtime="00:02:11.12" />
                    <SPLIT distance="200" swimtime="00:03:50.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-08-11" firstname="Agnieszka" gender="F" lastname="Drejka" nation="POL" athleteid="16164">
              <RESULTS>
                <RESULT eventid="1062" status="DNS" swimtime="00:00:00.00" resultid="16165" heatid="19278" lane="1" entrytime="00:00:39.00" />
                <RESULT eventid="1222" points="193" reactiontime="+97" swimtime="00:03:52.53" resultid="16166" heatid="19356" lane="2" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.81" />
                    <SPLIT distance="100" swimtime="00:01:50.88" />
                    <SPLIT distance="150" swimtime="00:02:52.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="183" swimtime="00:01:29.51" resultid="16167" heatid="19369" lane="0" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="176" reactiontime="+85" swimtime="00:01:51.24" resultid="16168" heatid="19429" lane="9" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="157" reactiontime="+100" swimtime="00:03:25.27" resultid="16169" heatid="19481" lane="1" entrytime="00:03:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.20" />
                    <SPLIT distance="100" swimtime="00:01:33.52" />
                    <SPLIT distance="150" swimtime="00:02:29.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="178" reactiontime="+90" swimtime="00:00:50.90" resultid="16170" heatid="19540" lane="4" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-13" firstname="Błażej" gender="M" lastname="Dyga" nation="POL" athleteid="16171">
              <RESULTS>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="16172" heatid="19374" lane="9" entrytime="00:03:00.00" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="16173" heatid="19472" lane="6" entrytime="00:01:40.00" />
                <RESULT eventid="1647" points="126" reactiontime="+102" swimtime="00:03:30.39" resultid="16174" heatid="19533" lane="7" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.70" />
                    <SPLIT distance="100" swimtime="00:01:42.64" />
                    <SPLIT distance="150" swimtime="00:02:35.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="161" reactiontime="+113" swimtime="00:06:29.41" resultid="16175" heatid="19702" lane="9" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.28" />
                    <SPLIT distance="100" swimtime="00:01:28.21" />
                    <SPLIT distance="150" swimtime="00:02:18.39" />
                    <SPLIT distance="200" swimtime="00:03:09.22" />
                    <SPLIT distance="250" swimtime="00:04:00.20" />
                    <SPLIT distance="300" swimtime="00:04:51.04" />
                    <SPLIT distance="350" swimtime="00:05:41.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-02-05" firstname="Zofia" gender="F" lastname="Dąbrowska" nation="POL" athleteid="16155">
              <RESULTS>
                <RESULT eventid="1062" points="167" reactiontime="+88" swimtime="00:00:42.18" resultid="16156" heatid="19277" lane="5" entrytime="00:00:41.00" />
                <RESULT eventid="1147" reactiontime="+86" status="OTL" swimtime="00:15:38.12" resultid="16157" heatid="19595" lane="8" entrytime="00:15:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.13" />
                    <SPLIT distance="100" swimtime="00:01:48.62" />
                    <SPLIT distance="150" swimtime="00:02:50.09" />
                    <SPLIT distance="200" swimtime="00:05:49.99" />
                    <SPLIT distance="300" swimtime="00:06:49.53" />
                    <SPLIT distance="350" swimtime="00:07:49.20" />
                    <SPLIT distance="400" swimtime="00:08:48.17" />
                    <SPLIT distance="450" swimtime="00:09:46.56" />
                    <SPLIT distance="600" swimtime="00:13:42.46" />
                    <SPLIT distance="650" swimtime="00:14:41.44" />
                    <SPLIT distance="700" swimtime="00:15:36.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="118" reactiontime="+88" swimtime="00:04:34.25" resultid="16158" heatid="19356" lane="8" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.11" />
                    <SPLIT distance="100" swimtime="00:02:03.64" />
                    <SPLIT distance="150" swimtime="00:03:15.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" status="DNS" swimtime="00:00:00.00" resultid="16159" heatid="19411" lane="5" entrytime="00:04:30.00" />
                <RESULT eventid="1388" points="143" reactiontime="+86" swimtime="00:01:59.10" resultid="16160" heatid="19428" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="103" reactiontime="+91" swimtime="00:09:13.28" resultid="16161" heatid="19503" lane="6" entrytime="00:08:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.94" />
                    <SPLIT distance="150" swimtime="00:03:42.78" />
                    <SPLIT distance="200" swimtime="00:04:57.48" />
                    <SPLIT distance="250" swimtime="00:06:09.55" />
                    <SPLIT distance="300" swimtime="00:07:19.73" />
                    <SPLIT distance="350" swimtime="00:08:18.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="84" reactiontime="+83" swimtime="00:02:04.51" resultid="16162" heatid="19513" lane="7" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="180" reactiontime="+78" swimtime="00:00:50.68" resultid="16163" heatid="19540" lane="6" entrytime="00:00:51.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" status="DNS" swimtime="00:00:00.00" resultid="16209" heatid="19500" lane="0" entrytime="00:02:12.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16202" number="1" />
                    <RELAYPOSITION athleteid="16176" number="2" />
                    <RELAYPOSITION athleteid="16181" number="3" />
                    <RELAYPOSITION athleteid="16189" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" status="DNS" swimtime="00:00:00.00" resultid="16210" heatid="19422" lane="9" entrytime="00:02:38.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16181" number="1" />
                    <RELAYPOSITION athleteid="16189" number="2" />
                    <RELAYPOSITION athleteid="16202" number="3" />
                    <RELAYPOSITION athleteid="16176" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" points="216" reactiontime="+78" swimtime="00:02:30.62" resultid="16211" heatid="19421" lane="4" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.35" />
                    <SPLIT distance="100" swimtime="00:01:20.95" />
                    <SPLIT distance="150" swimtime="00:01:48.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16181" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="16189" number="2" reactiontime="+43" />
                    <RELAYPOSITION athleteid="16202" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="16176" number="4" reactiontime="+71" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="236" reactiontime="+95" swimtime="00:02:23.13" resultid="16206" heatid="19320" lane="1" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.14" />
                    <SPLIT distance="100" swimtime="00:01:16.38" />
                    <SPLIT distance="150" swimtime="00:01:54.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16155" number="1" reactiontime="+95" />
                    <RELAYPOSITION athleteid="16181" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="16146" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="16189" number="4" reactiontime="-3" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="214" reactiontime="+82" swimtime="00:02:42.28" resultid="16207" heatid="19562" lane="8" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.67" />
                    <SPLIT distance="100" swimtime="00:01:39.63" />
                    <SPLIT distance="150" swimtime="00:02:07.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16146" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="16155" number="2" />
                    <RELAYPOSITION athleteid="16202" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="16181" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="CZE" clubid="14367" name="SK Spolchemie Usti nad Labem">
          <CONTACT email="benova.dana@seznam.cz" name="Spolchemie Usti nad Labem" phone="+420728212656" />
          <ATHLETES>
            <ATHLETE birthdate="1956-01-26" firstname="Dana" gender="F" lastname="Benova" nation="CZE" license="565126" athleteid="14368">
              <RESULTS>
                <RESULT eventid="1096" points="82" reactiontime="+87" swimtime="00:04:39.43" resultid="14369" heatid="19305" lane="2" entrytime="00:04:56.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.92" />
                    <SPLIT distance="100" swimtime="00:02:18.44" />
                    <SPLIT distance="150" swimtime="00:03:32.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="85" reactiontime="+98" swimtime="00:34:50.42" resultid="14370" heatid="19624" lane="0" entrytime="00:34:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.53" />
                    <SPLIT distance="100" swimtime="00:02:05.22" />
                    <SPLIT distance="150" swimtime="00:03:13.24" />
                    <SPLIT distance="200" swimtime="00:04:21.19" />
                    <SPLIT distance="250" swimtime="00:05:31.25" />
                    <SPLIT distance="300" swimtime="00:06:40.75" />
                    <SPLIT distance="350" swimtime="00:07:49.76" />
                    <SPLIT distance="400" swimtime="00:08:59.40" />
                    <SPLIT distance="450" swimtime="00:10:09.31" />
                    <SPLIT distance="500" swimtime="00:11:19.08" />
                    <SPLIT distance="550" swimtime="00:12:28.96" />
                    <SPLIT distance="600" swimtime="00:13:39.33" />
                    <SPLIT distance="650" swimtime="00:14:49.10" />
                    <SPLIT distance="700" swimtime="00:15:59.08" />
                    <SPLIT distance="750" swimtime="00:17:10.06" />
                    <SPLIT distance="800" swimtime="00:18:20.06" />
                    <SPLIT distance="850" swimtime="00:19:29.82" />
                    <SPLIT distance="900" swimtime="00:20:40.22" />
                    <SPLIT distance="950" swimtime="00:21:50.87" />
                    <SPLIT distance="1000" swimtime="00:23:02.04" />
                    <SPLIT distance="1050" swimtime="00:24:12.93" />
                    <SPLIT distance="1100" swimtime="00:25:23.90" />
                    <SPLIT distance="1150" swimtime="00:26:35.72" />
                    <SPLIT distance="1200" swimtime="00:27:46.85" />
                    <SPLIT distance="1250" swimtime="00:28:57.62" />
                    <SPLIT distance="1300" swimtime="00:30:09.42" />
                    <SPLIT distance="1350" swimtime="00:31:20.94" />
                    <SPLIT distance="1400" swimtime="00:32:32.42" />
                    <SPLIT distance="1450" swimtime="00:33:43.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="93" reactiontime="+93" swimtime="00:04:56.70" resultid="14371" heatid="19355" lane="6" entrytime="00:04:52.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.87" />
                    <SPLIT distance="100" swimtime="00:02:25.66" />
                    <SPLIT distance="150" swimtime="00:03:45.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="37" reactiontime="+92" swimtime="00:05:57.86" resultid="14372" heatid="19411" lane="2" entrytime="00:06:37.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.52" />
                    <SPLIT distance="100" swimtime="00:02:51.41" />
                    <SPLIT distance="150" swimtime="00:04:30.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="79" reactiontime="+89" swimtime="00:04:18.07" resultid="14373" heatid="19480" lane="9" entrytime="00:04:14.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.95" />
                    <SPLIT distance="100" swimtime="00:02:04.84" />
                    <SPLIT distance="150" swimtime="00:03:13.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="75" reactiontime="+98" swimtime="00:10:13.37" resultid="14374" heatid="19503" lane="2" entrytime="00:10:21.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.23" />
                    <SPLIT distance="150" swimtime="00:02:53.60" />
                    <SPLIT distance="200" swimtime="00:04:12.61" />
                    <SPLIT distance="250" swimtime="00:05:24.84" />
                    <SPLIT distance="300" swimtime="00:06:41.10" />
                    <SPLIT distance="350" swimtime="00:07:56.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="78" reactiontime="+83" swimtime="00:04:38.52" resultid="14375" heatid="19526" lane="5" entrytime="00:04:27.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.39" />
                    <SPLIT distance="100" swimtime="00:02:19.75" />
                    <SPLIT distance="150" swimtime="00:03:30.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="79" reactiontime="+89" swimtime="00:09:04.99" resultid="14376" heatid="19695" lane="7" entrytime="00:08:48.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.49" />
                    <SPLIT distance="100" swimtime="00:02:05.18" />
                    <SPLIT distance="150" swimtime="00:03:16.24" />
                    <SPLIT distance="200" swimtime="00:04:26.14" />
                    <SPLIT distance="250" swimtime="00:05:37.21" />
                    <SPLIT distance="300" swimtime="00:06:48.17" />
                    <SPLIT distance="350" swimtime="00:07:58.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="MAL" clubid="16274" name="Solne Miasto Wieliczka">
          <CONTACT email="zychkubaa@gmail.com" name="Zych Jakub" phone="784177829" />
          <ATHLETES>
            <ATHLETE birthdate="1960-03-20" firstname="Elżbieta" gender="F" lastname="Hamowska" nation="POL" athleteid="16295">
              <RESULTS>
                <RESULT eventid="1062" points="63" swimtime="00:00:58.27" resultid="16296" heatid="19276" lane="0" entrytime="00:00:55.00" />
                <RESULT comment="K11 - Nierównoczesne lub naprzemienne ruchy nóg (Time: 9:52)" eventid="1222" reactiontime="+88" status="DSQ" swimtime="00:04:51.74" resultid="16297" heatid="19356" lane="9" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.59" />
                    <SPLIT distance="100" swimtime="00:02:17.59" />
                    <SPLIT distance="150" swimtime="00:03:37.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="102" reactiontime="+97" swimtime="00:02:13.18" resultid="16298" heatid="19428" lane="8" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-03-23" firstname="Agnieszka" gender="F" lastname="Kuna" nation="POL" athleteid="16283">
              <RESULTS>
                <RESULT eventid="1096" points="102" reactiontime="+105" swimtime="00:04:20.53" resultid="16284" heatid="19306" lane="0" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.21" />
                    <SPLIT distance="100" swimtime="00:02:03.64" />
                    <SPLIT distance="150" swimtime="00:03:14.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="134" reactiontime="+114" swimtime="00:04:22.61" resultid="16285" heatid="19355" lane="5" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.60" />
                    <SPLIT distance="100" swimtime="00:02:00.63" />
                    <SPLIT distance="150" swimtime="00:03:11.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="173" reactiontime="+110" swimtime="00:01:51.80" resultid="16286" heatid="19428" lane="6" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-12-28" firstname="Darek" gender="M" lastname="Jania" nation="POL" athleteid="16275">
              <RESULTS>
                <RESULT eventid="1113" points="136" reactiontime="+90" swimtime="00:03:32.84" resultid="16276" heatid="19312" lane="5" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.32" />
                    <SPLIT distance="100" swimtime="00:01:43.00" />
                    <SPLIT distance="150" swimtime="00:02:39.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="151" reactiontime="+82" swimtime="00:01:34.40" resultid="16277" heatid="19400" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="152" reactiontime="+87" swimtime="00:00:40.79" resultid="16278" heatid="19452" lane="6" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-12-08" firstname="Jakub" gender="M" lastname="Jakubiński" nation="POL" athleteid="16299">
              <RESULTS>
                <RESULT eventid="1079" points="215" reactiontime="+86" swimtime="00:00:33.78" resultid="16300" heatid="19287" lane="5" entrytime="00:00:35.50" />
                <RESULT eventid="1273" points="160" reactiontime="+82" swimtime="00:01:22.63" resultid="16301" heatid="19376" lane="0" entrytime="00:01:29.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="135" reactiontime="+81" swimtime="00:03:13.70" resultid="16302" heatid="19487" lane="3" entrytime="00:03:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                    <SPLIT distance="100" swimtime="00:01:26.20" />
                    <SPLIT distance="150" swimtime="00:02:19.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-08-02" firstname="Edyta" gender="F" lastname="Żmijewska" nation="POL" athleteid="16291">
              <RESULTS>
                <RESULT eventid="1062" points="157" reactiontime="+98" swimtime="00:00:43.00" resultid="16292" heatid="19277" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="1187" points="123" reactiontime="+85" swimtime="00:00:51.50" resultid="16293" heatid="19337" lane="3" entrytime="00:00:50.00" />
                <RESULT eventid="1457" points="112" reactiontime="+81" swimtime="00:01:53.99" resultid="16294" heatid="19466" lane="1" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-02-07" firstname="Szymon" gender="M" lastname="Markiewicz" nation="POL" athleteid="16279">
              <RESULTS>
                <RESULT eventid="1079" points="168" reactiontime="+101" swimtime="00:00:36.70" resultid="16280" heatid="19288" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1273" points="171" reactiontime="+100" swimtime="00:01:20.85" resultid="16281" heatid="19376" lane="8" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="146" reactiontime="+100" swimtime="00:03:08.48" resultid="16282" heatid="19487" lane="4" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.19" />
                    <SPLIT distance="100" swimtime="00:01:25.40" />
                    <SPLIT distance="150" swimtime="00:02:16.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-03-27" firstname="Agnieszka" gender="F" lastname="DanekWiśniak" nation="POL" athleteid="16287">
              <RESULTS>
                <RESULT eventid="1062" points="137" reactiontime="+97" swimtime="00:00:45.03" resultid="16288" heatid="19277" lane="1" entrytime="00:00:43.00" />
                <RESULT eventid="1256" points="125" reactiontime="+97" swimtime="00:01:41.74" resultid="16289" heatid="19368" lane="8" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="129" reactiontime="+118" swimtime="00:03:38.99" resultid="16290" heatid="19480" lane="6" entrytime="00:03:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.12" />
                    <SPLIT distance="100" swimtime="00:01:45.71" />
                    <SPLIT distance="150" swimtime="00:02:44.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1358" points="124" reactiontime="+87" swimtime="00:03:26.60" resultid="16303" heatid="19419" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.94" />
                    <SPLIT distance="100" swimtime="00:01:51.14" />
                    <SPLIT distance="150" swimtime="00:02:40.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16291" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="16295" number="2" reactiontime="+100" />
                    <RELAYPOSITION athleteid="16283" number="3" reactiontime="+79" />
                    <RELAYPOSITION athleteid="16287" number="4" reactiontime="+74" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="174" reactiontime="+96" swimtime="00:02:38.41" resultid="16304" heatid="19319" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.13" />
                    <SPLIT distance="100" swimtime="00:01:28.64" />
                    <SPLIT distance="150" swimtime="00:02:04.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16283" number="1" reactiontime="+96" />
                    <RELAYPOSITION athleteid="16291" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="16279" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="16299" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="18444" name="Start Poznań">
          <CONTACT city="Poznań" email="robert.beym@gmail.com" name="Beym Robert" phone="512111513" street="os. Batorego 8/67" zip="60-687" />
          <ATHLETES>
            <ATHLETE birthdate="1982-07-01" firstname="Michał" gender="M" lastname="Kaczmarek" nation="POL" athleteid="18462">
              <RESULTS>
                <RESULT eventid="1273" points="273" reactiontime="+95" swimtime="00:01:09.25" resultid="18463" heatid="19379" lane="3" entrytime="00:01:10.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="242" reactiontime="+101" swimtime="00:01:20.71" resultid="18464" heatid="19401" lane="5" entrytime="00:01:22.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="262" reactiontime="+85" swimtime="00:01:26.82" resultid="18465" heatid="19437" lane="7" entrytime="00:01:29.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="176" reactiontime="+95" swimtime="00:00:38.83" resultid="18466" heatid="19453" lane="6" entrytime="00:00:36.97" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-07-01" firstname="Wojciech" gender="M" lastname="Dmytrów" nation="POL" athleteid="18467">
              <RESULTS>
                <RESULT eventid="1239" points="284" reactiontime="+95" swimtime="00:03:03.16" resultid="18468" heatid="19363" lane="0" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.10" />
                    <SPLIT distance="100" swimtime="00:01:23.62" />
                    <SPLIT distance="150" swimtime="00:02:12.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="357" reactiontime="+82" swimtime="00:01:18.36" resultid="18469" heatid="19439" lane="0" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="18470" heatid="19554" lane="8" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-07-01" firstname="Piotr" gender="M" lastname="Monczak" nation="POL" athleteid="18454">
              <RESULTS>
                <RESULT eventid="1079" points="419" reactiontime="+82" swimtime="00:00:27.07" resultid="18455" heatid="19300" lane="1" entrytime="00:00:26.40" />
                <RESULT eventid="1113" points="379" reactiontime="+86" swimtime="00:02:31.45" resultid="18456" heatid="19317" lane="1" entrytime="00:02:27.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                    <SPLIT distance="100" swimtime="00:01:10.81" />
                    <SPLIT distance="150" swimtime="00:01:56.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="457" reactiontime="+83" swimtime="00:00:58.33" resultid="18457" heatid="19386" lane="2" entrytime="00:00:57.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="380" swimtime="00:01:09.42" resultid="18458" heatid="19408" lane="0" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="434" swimtime="00:02:11.19" resultid="18459" heatid="19495" lane="0" entrytime="00:02:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                    <SPLIT distance="100" swimtime="00:01:04.54" />
                    <SPLIT distance="150" swimtime="00:01:37.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="18460" heatid="19511" lane="4" entrytime="00:05:25.00" />
                <RESULT eventid="1744" points="412" reactiontime="+84" swimtime="00:04:45.04" resultid="18461" heatid="19707" lane="4" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                    <SPLIT distance="100" swimtime="00:01:09.01" />
                    <SPLIT distance="150" swimtime="00:01:45.59" />
                    <SPLIT distance="200" swimtime="00:02:23.06" />
                    <SPLIT distance="250" swimtime="00:03:00.13" />
                    <SPLIT distance="300" swimtime="00:03:35.38" />
                    <SPLIT distance="350" swimtime="00:04:10.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-01-07" firstname="Robert" gender="M" lastname="Beym" nation="POL" athleteid="18445">
              <RESULTS>
                <RESULT eventid="1079" points="469" reactiontime="+83" swimtime="00:00:26.06" resultid="18446" heatid="19301" lane="5" entrytime="00:00:26.00" />
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="18447" heatid="19315" lane="6" entrytime="00:02:35.00" />
                <RESULT eventid="1205" points="371" reactiontime="+79" swimtime="00:00:30.91" resultid="18448" heatid="19351" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="14243" points="455" reactiontime="+83" swimtime="00:01:05.36" resultid="18449" heatid="19408" lane="5" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="453" reactiontime="+80" swimtime="00:00:28.38" resultid="18450" heatid="19460" lane="2" entrytime="00:00:29.00" />
                <RESULT eventid="1474" points="385" reactiontime="+81" swimtime="00:01:07.24" resultid="18451" heatid="19477" lane="4" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="420" reactiontime="+94" swimtime="00:01:04.18" resultid="18452" heatid="19523" lane="4" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="18453" heatid="19537" lane="8" entrytime="00:02:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="STEEF" nation="POL" region="DOL" clubid="18619" name="steef">
          <CONTACT city="Wrocław" email="ste1@wp.pl" name="Skrzypek Stefan" street="Edyty Stein" zip="50-322" />
          <ATHLETES>
            <ATHLETE birthdate="1956-09-02" firstname="Stefan" gender="M" lastname="Skrzypek" nation="POL" athleteid="18628">
              <RESULTS>
                <RESULT eventid="14207" points="167" reactiontime="+111" swimtime="00:25:38.48" resultid="18629" heatid="19620" lane="6" entrytime="00:26:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.17" />
                    <SPLIT distance="100" swimtime="00:01:30.13" />
                    <SPLIT distance="150" swimtime="00:02:17.84" />
                    <SPLIT distance="200" swimtime="00:03:06.43" />
                    <SPLIT distance="250" swimtime="00:03:55.61" />
                    <SPLIT distance="300" swimtime="00:04:47.06" />
                    <SPLIT distance="350" swimtime="00:05:38.15" />
                    <SPLIT distance="400" swimtime="00:06:29.62" />
                    <SPLIT distance="450" swimtime="00:07:21.48" />
                    <SPLIT distance="500" swimtime="00:08:13.82" />
                    <SPLIT distance="550" swimtime="00:09:05.02" />
                    <SPLIT distance="600" swimtime="00:09:56.83" />
                    <SPLIT distance="650" swimtime="00:10:48.79" />
                    <SPLIT distance="700" swimtime="00:11:39.96" />
                    <SPLIT distance="750" swimtime="00:12:32.09" />
                    <SPLIT distance="800" swimtime="00:13:23.89" />
                    <SPLIT distance="850" swimtime="00:14:15.50" />
                    <SPLIT distance="900" swimtime="00:15:09.15" />
                    <SPLIT distance="950" swimtime="00:16:02.53" />
                    <SPLIT distance="1000" swimtime="00:16:56.50" />
                    <SPLIT distance="1050" swimtime="00:17:49.05" />
                    <SPLIT distance="1100" swimtime="00:18:42.02" />
                    <SPLIT distance="1150" swimtime="00:19:35.28" />
                    <SPLIT distance="1200" swimtime="00:20:28.33" />
                    <SPLIT distance="1250" swimtime="00:21:21.80" />
                    <SPLIT distance="1300" swimtime="00:22:14.35" />
                    <SPLIT distance="1350" swimtime="00:23:07.05" />
                    <SPLIT distance="1400" swimtime="00:24:00.19" />
                    <SPLIT distance="1450" swimtime="00:24:51.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="198" reactiontime="+106" swimtime="00:02:50.26" resultid="18630" heatid="19489" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.58" />
                    <SPLIT distance="100" swimtime="00:01:21.59" />
                    <SPLIT distance="150" swimtime="00:02:05.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="183" reactiontime="+99" swimtime="00:06:13.55" resultid="18631" heatid="19703" lane="8" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.90" />
                    <SPLIT distance="100" swimtime="00:01:29.71" />
                    <SPLIT distance="150" swimtime="00:02:17.66" />
                    <SPLIT distance="200" swimtime="00:03:06.32" />
                    <SPLIT distance="250" swimtime="00:03:54.40" />
                    <SPLIT distance="300" swimtime="00:04:42.18" />
                    <SPLIT distance="350" swimtime="00:05:29.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-03-19" firstname="Ewa" gender="F" lastname="Szała" nation="POL" athleteid="18620">
              <RESULTS>
                <RESULT eventid="1096" points="283" reactiontime="+93" swimtime="00:03:05.58" resultid="18621" heatid="19307" lane="2" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.71" />
                    <SPLIT distance="100" swimtime="00:01:27.71" />
                    <SPLIT distance="150" swimtime="00:02:19.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="269" reactiontime="+93" swimtime="00:00:39.76" resultid="18622" heatid="19338" lane="4" entrytime="00:00:41.00" />
                <RESULT eventid="14225" points="261" reactiontime="+82" swimtime="00:01:28.60" resultid="18623" heatid="19393" lane="9" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="259" swimtime="00:01:26.27" resultid="18624" heatid="19467" lane="2" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="281" reactiontime="+97" swimtime="00:06:35.69" resultid="18625" heatid="19504" lane="6" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.52" />
                    <SPLIT distance="100" swimtime="00:01:37.59" />
                    <SPLIT distance="150" swimtime="00:02:26.03" />
                    <SPLIT distance="200" swimtime="00:03:16.17" />
                    <SPLIT distance="250" swimtime="00:04:10.19" />
                    <SPLIT distance="300" swimtime="00:05:06.10" />
                    <SPLIT distance="350" swimtime="00:05:51.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="261" swimtime="00:03:06.45" resultid="18626" heatid="19528" lane="1" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.69" />
                    <SPLIT distance="100" swimtime="00:01:31.65" />
                    <SPLIT distance="150" swimtime="00:02:20.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="248" reactiontime="+99" swimtime="00:06:12.87" resultid="18627" heatid="19697" lane="8" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                    <SPLIT distance="100" swimtime="00:02:16.46" />
                    <SPLIT distance="150" swimtime="00:03:03.93" />
                    <SPLIT distance="200" swimtime="00:03:50.50" />
                    <SPLIT distance="250" swimtime="00:04:37.35" />
                    <SPLIT distance="300" swimtime="00:05:25.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MASTERS LU" nation="POL" region="LBL" clubid="14934" name="Stowarzyszenie Pływackie MASTERS Lublin" shortname="Stowarzyszenie Pływackie MASTE">
          <CONTACT city="Lublin" email="masters_lublin@wp.pl" name="Rafał Wójcicki" phone="+48501794954" state="LUBEL" street="Stanisława Lema 18" zip="20-445" />
          <ATHLETES>
            <ATHLETE birthdate="1975-04-28" firstname="Rafał" gender="M" lastname="Wójcicki" nation="POL" license="103503700001" athleteid="14935">
              <RESULTS>
                <RESULT eventid="1205" points="242" reactiontime="+72" swimtime="00:00:35.64" resultid="14936" heatid="19348" lane="3" entrytime="00:00:35.53" entrycourse="SCM" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="14937" heatid="19475" lane="1" entrytime="00:01:17.64" entrycourse="SCM" />
                <RESULT eventid="1681" points="282" reactiontime="+82" swimtime="00:00:38.46" resultid="14938" heatid="19553" lane="8" entrytime="00:00:38.42" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-11-07" firstname="Konrad" gender="M" lastname="Ćwikła" nation="POL" license="103503700005" athleteid="14948">
              <RESULTS>
                <RESULT eventid="14243" points="358" reactiontime="+101" swimtime="00:01:10.80" resultid="14949" heatid="19405" lane="1" entrytime="00:01:12.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="324" reactiontime="+95" swimtime="00:00:31.74" resultid="14950" heatid="19459" lane="8" entrytime="00:00:30.59" entrycourse="SCM" />
                <RESULT eventid="1744" points="283" reactiontime="+90" swimtime="00:05:22.91" resultid="14951" heatid="19704" lane="8" entrytime="00:05:30.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.17" />
                    <SPLIT distance="100" swimtime="00:01:13.56" />
                    <SPLIT distance="150" swimtime="00:01:54.34" />
                    <SPLIT distance="200" swimtime="00:02:35.49" />
                    <SPLIT distance="250" swimtime="00:04:00.14" />
                    <SPLIT distance="300" swimtime="00:04:42.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-06-05" firstname="Marek" gender="M" lastname="Żuber" nation="POL" license="103503700009" athleteid="14952">
              <RESULTS>
                <RESULT eventid="1079" points="352" reactiontime="+90" swimtime="00:00:28.69" resultid="14953" heatid="19300" lane="6" entrytime="00:00:26.11" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-05-28" firstname="Anna" gender="F" lastname="Michalska" nation="POL" license="103503600002" athleteid="14939">
              <RESULTS>
                <RESULT eventid="1062" points="331" swimtime="00:00:33.57" resultid="14940" heatid="19281" lane="0" entrytime="00:00:32.88" entrycourse="SCM" />
                <RESULT eventid="1187" points="357" reactiontime="+88" swimtime="00:00:36.16" resultid="14941" heatid="19340" lane="2" entrytime="00:00:35.54" entrycourse="SCM" />
                <RESULT eventid="1457" points="329" reactiontime="+89" swimtime="00:01:19.66" resultid="14942" heatid="19468" lane="7" entrytime="00:01:19.76" entrycourse="SCM" />
                <RESULT eventid="1630" points="329" reactiontime="+95" swimtime="00:02:52.66" resultid="14943" heatid="19528" lane="3" entrytime="00:02:58.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.30" />
                    <SPLIT distance="100" swimtime="00:01:22.62" />
                    <SPLIT distance="150" swimtime="00:02:08.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-26" firstname="Rafał" gender="M" lastname="Zielonka" nation="POL" license="103503700008" athleteid="14944">
              <RESULTS>
                <RESULT eventid="14189" points="459" reactiontime="+80" swimtime="00:09:34.53" resultid="14945" heatid="19618" lane="7" entrytime="00:09:30.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.39" />
                    <SPLIT distance="100" swimtime="00:01:05.92" />
                    <SPLIT distance="150" swimtime="00:01:41.13" />
                    <SPLIT distance="200" swimtime="00:02:17.23" />
                    <SPLIT distance="250" swimtime="00:02:52.72" />
                    <SPLIT distance="300" swimtime="00:03:28.82" />
                    <SPLIT distance="350" swimtime="00:04:05.13" />
                    <SPLIT distance="400" swimtime="00:04:41.56" />
                    <SPLIT distance="450" swimtime="00:05:17.63" />
                    <SPLIT distance="500" swimtime="00:05:53.88" />
                    <SPLIT distance="550" swimtime="00:06:30.56" />
                    <SPLIT distance="600" swimtime="00:07:07.71" />
                    <SPLIT distance="650" swimtime="00:07:44.68" />
                    <SPLIT distance="700" swimtime="00:08:21.66" />
                    <SPLIT distance="750" swimtime="00:08:58.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="511" reactiontime="+91" swimtime="00:02:04.29" resultid="14946" heatid="19495" lane="2" entrytime="00:02:07.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.01" />
                    <SPLIT distance="100" swimtime="00:01:00.83" />
                    <SPLIT distance="150" swimtime="00:01:33.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="497" reactiontime="+87" swimtime="00:04:27.81" resultid="14947" heatid="19708" lane="2" entrytime="00:04:29.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                    <SPLIT distance="100" swimtime="00:01:03.23" />
                    <SPLIT distance="150" swimtime="00:01:36.62" />
                    <SPLIT distance="200" swimtime="00:02:10.68" />
                    <SPLIT distance="250" swimtime="00:02:44.74" />
                    <SPLIT distance="300" swimtime="00:03:19.74" />
                    <SPLIT distance="350" swimtime="00:03:54.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="MASTERS Lublin" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="360" reactiontime="+74" swimtime="00:02:07.12" resultid="14954" heatid="19423" lane="0" entrytime="00:02:10.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                    <SPLIT distance="100" swimtime="00:01:08.30" />
                    <SPLIT distance="150" swimtime="00:01:39.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14935" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="14944" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="14952" number="3" reactiontime="+75" />
                    <RELAYPOSITION athleteid="14948" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="404" reactiontime="+102" swimtime="00:01:51.69" resultid="14955" heatid="19501" lane="1" entrytime="00:01:55.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.11" />
                    <SPLIT distance="100" swimtime="00:00:57.98" />
                    <SPLIT distance="150" swimtime="00:01:26.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14948" number="1" reactiontime="+102" />
                    <RELAYPOSITION athleteid="14935" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="14952" number="3" reactiontime="+143" />
                    <RELAYPOSITION athleteid="14944" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="17684" name="Swim2tri">
          <CONTACT name="Hanczewska Marta" />
          <ATHLETES>
            <ATHLETE birthdate="1984-10-05" firstname="Marta" gender="F" lastname="Hanczewska" nation="POL" athleteid="17685">
              <RESULTS>
                <RESULT eventid="1062" points="362" reactiontime="+98" swimtime="00:00:32.59" resultid="17686" heatid="19280" lane="2" entrytime="00:00:33.50" />
                <RESULT eventid="14225" points="293" reactiontime="+95" swimtime="00:01:25.32" resultid="17687" heatid="19392" lane="6" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="299" reactiontime="+98" swimtime="00:01:33.19" resultid="17688" heatid="19430" lane="3" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="308" reactiontime="+90" swimtime="00:00:42.37" resultid="17689" heatid="19543" lane="9" entrytime="00:00:41.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="079/14" nation="POL" region="WA" clubid="17269" name="Swimmers St. Pływackie">
          <CONTACT city="WARSZAWA" email="REMOG@SWIMMERSTEAM.PL" name="GOŁĘBIOWSKI REMIGIUSZ" phone="601333782" state="MAZ" street="GŁADKA 18" zip="02-172" />
          <ATHLETES>
            <ATHLETE birthdate="1993-03-07" firstname="Michał" gender="M" lastname="Hudyka" nation="POL" athleteid="17278">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="17279" heatid="19299" lane="2" entrytime="00:00:27.00" />
                <RESULT eventid="14243" status="DNS" swimtime="00:00:00.00" resultid="17280" heatid="19406" lane="5" entrytime="00:01:09.00" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="17281" heatid="19558" lane="9" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-28" firstname="Marek" gender="M" lastname="Brożyna" nation="POL" athleteid="17270">
              <RESULTS>
                <RESULT eventid="1079" points="323" reactiontime="+88" swimtime="00:00:29.50" resultid="17271" heatid="19296" lane="4" entrytime="00:00:28.39" />
                <RESULT eventid="1113" points="324" reactiontime="+78" swimtime="00:02:39.47" resultid="17272" heatid="19314" lane="9" entrytime="00:02:44.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                    <SPLIT distance="100" swimtime="00:01:14.88" />
                    <SPLIT distance="150" swimtime="00:02:04.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="303" reactiontime="+73" swimtime="00:00:33.05" resultid="17273" heatid="19349" lane="6" entrytime="00:00:33.24" />
                <RESULT eventid="14243" points="332" reactiontime="+88" swimtime="00:01:12.57" resultid="17274" heatid="19404" lane="4" entrytime="00:01:13.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="317" swimtime="00:01:11.73" resultid="17275" heatid="19476" lane="7" entrytime="00:01:12.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="319" reactiontime="+90" swimtime="00:05:44.50" resultid="17276" heatid="19509" lane="4" entrytime="00:06:06.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.67" />
                    <SPLIT distance="100" swimtime="00:01:19.17" />
                    <SPLIT distance="150" swimtime="00:02:01.59" />
                    <SPLIT distance="200" swimtime="00:02:42.46" />
                    <SPLIT distance="250" swimtime="00:03:33.91" />
                    <SPLIT distance="300" swimtime="00:04:25.29" />
                    <SPLIT distance="350" swimtime="00:05:06.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="329" swimtime="00:02:32.87" resultid="17277" heatid="19536" lane="1" entrytime="00:02:38.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.46" />
                    <SPLIT distance="100" swimtime="00:01:13.49" />
                    <SPLIT distance="150" swimtime="00:01:53.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="17879" name="Swimminmg Masters Team Szczecin" shortname="Swimminmg Masters Team Szczeci">
          <CONTACT city="Szczecin" email="aga.krzyzostaniak@gmail.com" name="Krzyżostaniak Agnieszka" phone="603772862" street="Żupańskiego 12/8" zip="71-440" />
          <ATHLETES>
            <ATHLETE birthdate="1996-02-15" firstname="Filip" gender="M" lastname="Przybyłowski" nation="POL" athleteid="17988">
              <RESULTS>
                <RESULT eventid="14189" reactiontime="+66" status="OTL" swimtime="00:10:13.07" resultid="17989" heatid="19617" lane="4" entrytime="00:10:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                    <SPLIT distance="100" swimtime="00:01:09.70" />
                    <SPLIT distance="150" swimtime="00:01:47.43" />
                    <SPLIT distance="200" swimtime="00:02:26.22" />
                    <SPLIT distance="250" swimtime="00:03:05.04" />
                    <SPLIT distance="300" swimtime="00:03:44.18" />
                    <SPLIT distance="350" swimtime="00:04:23.48" />
                    <SPLIT distance="400" swimtime="00:05:02.26" />
                    <SPLIT distance="450" swimtime="00:05:41.92" />
                    <SPLIT distance="500" swimtime="00:06:21.56" />
                    <SPLIT distance="550" swimtime="00:07:01.89" />
                    <SPLIT distance="600" swimtime="00:07:41.43" />
                    <SPLIT distance="650" swimtime="00:08:20.88" />
                    <SPLIT distance="700" swimtime="00:08:59.84" />
                    <SPLIT distance="750" swimtime="00:09:38.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="393" reactiontime="+68" swimtime="00:00:29.74" resultid="17990" heatid="19456" lane="3" entrytime="00:00:32.13" entrycourse="SCM" />
                <RESULT comment="K16 - Niejednoczesne dotknięcie ściany dłońmi przy nawrocie lub na zakończenie wyścigu (Time: 21:05)" eventid="1578" reactiontime="+69" status="DSQ" swimtime="00:05:27.00" resultid="17991" heatid="19510" lane="3" entrytime="00:05:57.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                    <SPLIT distance="100" swimtime="00:01:11.79" />
                    <SPLIT distance="150" swimtime="00:01:55.96" />
                    <SPLIT distance="200" swimtime="00:02:40.29" />
                    <SPLIT distance="250" swimtime="00:03:27.22" />
                    <SPLIT distance="300" swimtime="00:04:14.40" />
                    <SPLIT distance="350" swimtime="00:04:52.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="372" reactiontime="+70" swimtime="00:01:06.80" resultid="17992" heatid="19521" lane="1" entrytime="00:01:13.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-11-04" firstname="Kamil" gender="M" lastname="Zieliński" nation="POL" athleteid="17934">
              <RESULTS>
                <RESULT eventid="14189" reactiontime="+98" status="OTL" swimtime="00:12:06.36" resultid="17935" heatid="19616" lane="8" entrytime="00:12:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.28" />
                    <SPLIT distance="100" swimtime="00:02:48.55" />
                    <SPLIT distance="600" swimtime="00:08:17.63" />
                    <SPLIT distance="650" swimtime="00:09:04.88" />
                    <SPLIT distance="700" swimtime="00:10:37.17" />
                    <SPLIT distance="750" swimtime="00:11:24.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="198" reactiontime="+74" swimtime="00:00:38.09" resultid="17936" heatid="19346" lane="5" entrytime="00:00:40.00" entrycourse="SCM" />
                <RESULT eventid="1273" points="253" reactiontime="+96" swimtime="00:01:10.99" resultid="17937" heatid="19379" lane="2" entrytime="00:01:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="184" reactiontime="+72" swimtime="00:01:25.93" resultid="17938" heatid="19473" lane="2" entrytime="00:01:30.00" entrycourse="SCM" />
                <RESULT eventid="1647" points="171" reactiontime="+80" swimtime="00:03:10.25" resultid="17939" heatid="19533" lane="3" entrytime="00:03:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.17" />
                    <SPLIT distance="100" swimtime="00:01:29.96" />
                    <SPLIT distance="150" swimtime="00:02:21.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-17" firstname="Grzegorz" gender="M" lastname="Juszkiewicz" nation="POL" athleteid="17993">
              <RESULTS>
                <RESULT eventid="1273" points="88" reactiontime="+185" swimtime="00:01:40.86" resultid="17994" heatid="19374" lane="4" entrytime="00:01:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="65" reactiontime="+127" swimtime="00:02:05.05" resultid="17995" heatid="19398" lane="9" entrytime="00:02:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-06-09" firstname="Marcin" gender="M" lastname="Kaczmarek" nation="POL" athleteid="17996">
              <RESULTS>
                <RESULT eventid="1273" points="198" reactiontime="+84" swimtime="00:01:17.01" resultid="17997" heatid="19376" lane="4" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="170" reactiontime="+82" swimtime="00:02:59.32" resultid="17998" heatid="19487" lane="6" entrytime="00:03:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.58" />
                    <SPLIT distance="100" swimtime="00:01:26.96" />
                    <SPLIT distance="150" swimtime="00:02:14.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="17999" heatid="19700" lane="2" entrytime="00:07:20.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-03-20" firstname="Marcin" gender="M" lastname="Łogin" nation="POL" athleteid="18000">
              <RESULTS>
                <RESULT eventid="1079" points="298" reactiontime="+109" swimtime="00:00:30.33" resultid="18001" heatid="19293" lane="0" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="1239" points="234" reactiontime="+103" swimtime="00:03:15.26" resultid="18002" heatid="19362" lane="1" entrytime="00:03:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.85" />
                    <SPLIT distance="100" swimtime="00:01:34.71" />
                    <SPLIT distance="150" swimtime="00:02:25.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="264" reactiontime="+105" swimtime="00:01:26.68" resultid="18003" heatid="19438" lane="3" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="18004" heatid="19554" lane="0" entrytime="00:00:37.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-09" firstname="Helena" gender="F" lastname="Szulc" nation="POL" athleteid="17960">
              <RESULTS>
                <RESULT eventid="1096" points="314" reactiontime="+92" swimtime="00:02:59.17" resultid="17961" heatid="19308" lane="0" entrytime="00:03:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.51" />
                    <SPLIT distance="100" swimtime="00:01:23.39" />
                    <SPLIT distance="150" swimtime="00:02:15.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="347" reactiontime="+85" swimtime="00:01:20.63" resultid="17962" heatid="19394" lane="8" entrytime="00:01:21.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="227" reactiontime="+97" swimtime="00:03:16.02" resultid="17963" heatid="19412" lane="1" entrytime="00:03:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.21" />
                    <SPLIT distance="100" swimtime="00:01:34.34" />
                    <SPLIT distance="150" swimtime="00:02:26.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="305" swimtime="00:00:36.21" resultid="17964" heatid="19447" lane="0" entrytime="00:00:37.00" entrycourse="SCM" />
                <RESULT eventid="1555" points="299" reactiontime="+100" swimtime="00:06:27.81" resultid="17965" heatid="19504" lane="4" entrytime="00:06:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.70" />
                    <SPLIT distance="100" swimtime="00:01:33.61" />
                    <SPLIT distance="150" swimtime="00:02:22.96" />
                    <SPLIT distance="200" swimtime="00:03:11.30" />
                    <SPLIT distance="250" swimtime="00:04:05.21" />
                    <SPLIT distance="300" swimtime="00:04:59.98" />
                    <SPLIT distance="350" swimtime="00:05:44.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="267" reactiontime="+86" swimtime="00:01:24.77" resultid="17966" heatid="19515" lane="8" entrytime="00:01:23.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-05-09" firstname="Łukasz" gender="M" lastname="Rożek" nation="POL" athleteid="17982">
              <RESULTS>
                <RESULT eventid="1079" points="200" reactiontime="+113" swimtime="00:00:34.59" resultid="17983" heatid="19289" lane="7" entrytime="00:00:33.14" entrycourse="SCM" />
                <RESULT eventid="14189" reactiontime="+101" status="OTL" swimtime="00:14:04.01" resultid="17984" heatid="19615" lane="6" entrytime="00:14:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.82" />
                    <SPLIT distance="100" swimtime="00:01:33.47" />
                    <SPLIT distance="150" swimtime="00:02:23.19" />
                    <SPLIT distance="200" swimtime="00:03:15.19" />
                    <SPLIT distance="250" swimtime="00:04:08.56" />
                    <SPLIT distance="300" swimtime="00:05:03.38" />
                    <SPLIT distance="350" swimtime="00:05:57.61" />
                    <SPLIT distance="400" swimtime="00:06:53.01" />
                    <SPLIT distance="450" swimtime="00:07:48.16" />
                    <SPLIT distance="500" swimtime="00:08:42.77" />
                    <SPLIT distance="550" swimtime="00:09:37.17" />
                    <SPLIT distance="600" swimtime="00:10:31.45" />
                    <SPLIT distance="650" swimtime="00:11:25.55" />
                    <SPLIT distance="700" swimtime="00:12:20.81" />
                    <SPLIT distance="750" swimtime="00:13:14.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="217" reactiontime="+83" swimtime="00:01:14.74" resultid="17985" heatid="19377" lane="7" entrytime="00:01:20.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="181" reactiontime="+92" swimtime="00:02:55.64" resultid="17986" heatid="19487" lane="5" entrytime="00:03:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.08" />
                    <SPLIT distance="100" swimtime="00:01:22.47" />
                    <SPLIT distance="150" swimtime="00:02:09.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="154" reactiontime="+86" swimtime="00:06:35.27" resultid="17987" heatid="19700" lane="4" entrytime="00:07:05.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.13" />
                    <SPLIT distance="100" swimtime="00:01:27.73" />
                    <SPLIT distance="150" swimtime="00:02:16.42" />
                    <SPLIT distance="200" swimtime="00:03:06.32" />
                    <SPLIT distance="250" swimtime="00:03:56.86" />
                    <SPLIT distance="300" swimtime="00:04:49.46" />
                    <SPLIT distance="350" swimtime="00:05:42.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-03-13" firstname="Boguś" gender="M" lastname="Michalak" nation="POL" athleteid="18005">
              <RESULTS>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="18006" heatid="19344" lane="5" entrytime="00:00:50.00" entrycourse="SCM" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="18007" heatid="19374" lane="1" entrytime="00:02:15.00" entrycourse="SCM" />
                <RESULT comment="K14 - Praca nóg w płaszczyźnie pionowej w dół (z wyjątkiem jednego ruchu po starcie i nawrocie) (Time: 16:39)" eventid="1406" reactiontime="+119" status="DSQ" swimtime="00:02:27.10" resultid="18008" heatid="19434" lane="9" entrytime="00:02:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="40" reactiontime="+104" swimtime="00:02:22.36" resultid="18009" heatid="19470" lane="3" entrytime="00:02:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-12-12" firstname="Dominika" gender="F" lastname="Zielińska" nation="POL" athleteid="17926">
              <RESULTS>
                <RESULT eventid="1096" points="424" reactiontime="+89" swimtime="00:02:42.13" resultid="17927" heatid="19308" lane="4" entrytime="00:02:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                    <SPLIT distance="100" swimtime="00:01:15.10" />
                    <SPLIT distance="150" swimtime="00:02:02.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="371" reactiontime="+90" swimtime="00:11:06.56" resultid="17928" heatid="19596" lane="7" entrytime="00:10:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                    <SPLIT distance="100" swimtime="00:01:16.18" />
                    <SPLIT distance="150" swimtime="00:01:57.55" />
                    <SPLIT distance="200" swimtime="00:02:39.46" />
                    <SPLIT distance="250" swimtime="00:03:21.92" />
                    <SPLIT distance="300" swimtime="00:04:04.45" />
                    <SPLIT distance="350" swimtime="00:04:47.04" />
                    <SPLIT distance="400" swimtime="00:05:29.86" />
                    <SPLIT distance="450" swimtime="00:06:12.75" />
                    <SPLIT distance="500" swimtime="00:06:55.13" />
                    <SPLIT distance="550" swimtime="00:07:37.25" />
                    <SPLIT distance="600" swimtime="00:08:20.35" />
                    <SPLIT distance="650" swimtime="00:09:02.43" />
                    <SPLIT distance="700" swimtime="00:09:44.51" />
                    <SPLIT distance="750" swimtime="00:10:25.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="373" reactiontime="+57" swimtime="00:00:35.64" resultid="17929" heatid="19340" lane="7" entrytime="00:00:36.00" entrycourse="SCM" />
                <RESULT eventid="14225" points="422" reactiontime="+87" swimtime="00:01:15.51" resultid="17930" heatid="19394" lane="3" entrytime="00:01:16.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="385" reactiontime="+74" swimtime="00:01:15.58" resultid="17931" heatid="19468" lane="3" entrytime="00:01:16.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="405" reactiontime="+70" swimtime="00:02:29.62" resultid="17932" heatid="19484" lane="0" entrytime="00:02:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.62" />
                    <SPLIT distance="100" swimtime="00:01:11.19" />
                    <SPLIT distance="150" swimtime="00:01:50.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="383" swimtime="00:02:44.07" resultid="17933" heatid="19529" lane="8" entrytime="00:02:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:02:02.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-05-26" firstname="Grzegorz" gender="M" lastname="Król" nation="POL" athleteid="17969">
              <RESULTS>
                <RESULT eventid="1205" reactiontime="+123" status="DNS" swimtime="00:00:00.00" resultid="17970" heatid="19346" lane="3" entrytime="00:00:40.00" entrycourse="SCM" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="17971" heatid="19373" lane="4" entrytime="00:01:47.00" entrycourse="SCM" />
                <RESULT eventid="1508" points="151" reactiontime="+113" swimtime="00:03:06.25" resultid="17972" heatid="19489" lane="6" entrytime="00:02:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.24" />
                    <SPLIT distance="100" swimtime="00:01:24.68" />
                    <SPLIT distance="150" swimtime="00:02:16.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-06-19" firstname="Tomasz" gender="M" lastname="Mazur" nation="POL" athleteid="17967">
              <RESULTS>
                <RESULT eventid="1273" points="127" reactiontime="+89" swimtime="00:01:29.23" resultid="17968" heatid="19375" lane="3" entrytime="00:01:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-29" firstname="Robert" gender="M" lastname="Szota" nation="POL" athleteid="17973">
              <RESULTS>
                <RESULT eventid="1079" points="366" reactiontime="+77" swimtime="00:00:28.31" resultid="17974" heatid="19292" lane="5" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="14189" reactiontime="+79" status="OTL" swimtime="00:10:37.40" resultid="17975" heatid="19617" lane="5" entrytime="00:10:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.00" />
                    <SPLIT distance="100" swimtime="00:01:11.90" />
                    <SPLIT distance="150" swimtime="00:01:50.92" />
                    <SPLIT distance="200" swimtime="00:02:30.12" />
                    <SPLIT distance="250" swimtime="00:03:09.76" />
                    <SPLIT distance="300" swimtime="00:03:49.82" />
                    <SPLIT distance="350" swimtime="00:04:30.78" />
                    <SPLIT distance="400" swimtime="00:05:11.40" />
                    <SPLIT distance="450" swimtime="00:05:52.16" />
                    <SPLIT distance="500" swimtime="00:06:33.73" />
                    <SPLIT distance="550" swimtime="00:07:15.01" />
                    <SPLIT distance="600" swimtime="00:07:56.66" />
                    <SPLIT distance="700" swimtime="00:09:19.14" />
                    <SPLIT distance="750" swimtime="00:09:59.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="356" reactiontime="+73" swimtime="00:01:03.35" resultid="17976" heatid="19382" lane="8" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="319" swimtime="00:01:13.56" resultid="17977" heatid="19403" lane="0" entrytime="00:01:17.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="285" reactiontime="+66" swimtime="00:00:33.09" resultid="17978" heatid="19455" lane="8" entrytime="00:00:34.50" entrycourse="SCM" />
                <RESULT eventid="1508" points="349" reactiontime="+70" swimtime="00:02:21.09" resultid="17979" heatid="19492" lane="3" entrytime="00:02:23.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                    <SPLIT distance="100" swimtime="00:01:09.41" />
                    <SPLIT distance="150" swimtime="00:01:46.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="280" reactiontime="+77" swimtime="00:00:38.59" resultid="17980" heatid="19553" lane="7" entrytime="00:00:38.00" entrycourse="SCM" />
                <RESULT eventid="1744" points="332" reactiontime="+71" swimtime="00:05:06.49" resultid="17981" heatid="19706" lane="9" entrytime="00:05:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                    <SPLIT distance="100" swimtime="00:01:12.79" />
                    <SPLIT distance="150" swimtime="00:01:52.12" />
                    <SPLIT distance="200" swimtime="00:02:31.93" />
                    <SPLIT distance="300" swimtime="00:03:52.14" />
                    <SPLIT distance="350" swimtime="00:04:31.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-06-12" firstname="Kamila" gender="F" lastname="Gębka" nation="POL" athleteid="17947">
              <RESULTS>
                <RESULT eventid="1222" points="317" reactiontime="+98" swimtime="00:03:17.23" resultid="17948" heatid="19356" lane="7" entrytime="00:03:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.14" />
                    <SPLIT distance="100" swimtime="00:01:36.41" />
                    <SPLIT distance="150" swimtime="00:02:25.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" status="DNS" swimtime="00:00:00.00" resultid="17949" heatid="19429" lane="6" entrytime="00:01:40.00" entrycourse="SCM" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="17950" heatid="19483" lane="9" entrytime="00:02:50.00" entrycourse="SCM" />
                <RESULT eventid="1664" status="DNS" swimtime="00:00:00.00" resultid="17951" heatid="19541" lane="5" entrytime="00:00:45.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-02-24" firstname="Maciej" gender="M" lastname="Brodacki" nation="POL" athleteid="17914">
              <RESULTS>
                <RESULT eventid="1079" points="514" reactiontime="+88" swimtime="00:00:25.28" resultid="17915" heatid="19301" lane="1" entrytime="00:00:26.00" entrycourse="SCM" />
                <RESULT eventid="1273" points="521" reactiontime="+79" swimtime="00:00:55.84" resultid="17916" heatid="19387" lane="8" entrytime="00:00:56.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="458" reactiontime="+83" swimtime="00:01:05.23" resultid="17917" heatid="19408" lane="4" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="448" reactiontime="+82" swimtime="00:00:28.47" resultid="17918" heatid="19460" lane="6" entrytime="00:00:29.00" entrycourse="SCM" />
                <RESULT eventid="1474" points="377" reactiontime="+87" swimtime="00:01:07.71" resultid="17919" heatid="19475" lane="0" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="436" reactiontime="+85" swimtime="00:01:03.40" resultid="17920" heatid="19523" lane="5" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="400" reactiontime="+85" swimtime="00:00:34.26" resultid="17921" heatid="19554" lane="2" entrytime="00:00:37.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-08-12" firstname="Marek" gender="M" lastname="Zienkiewicz" nation="POL" athleteid="17952">
              <RESULTS>
                <RESULT eventid="1079" points="334" reactiontime="+82" swimtime="00:00:29.20" resultid="17953" heatid="19293" lane="5" entrytime="00:00:29.59" entrycourse="SCM" />
                <RESULT eventid="1273" points="288" reactiontime="+74" swimtime="00:01:07.98" resultid="17954" heatid="19380" lane="7" entrytime="00:01:08.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="245" reactiontime="+82" swimtime="00:01:20.28" resultid="17955" heatid="19402" lane="2" entrytime="00:01:19.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="298" reactiontime="+76" swimtime="00:00:32.61" resultid="17956" heatid="19456" lane="0" entrytime="00:00:32.97" entrycourse="SCM" />
                <RESULT eventid="1508" points="242" reactiontime="+73" swimtime="00:02:39.36" resultid="17957" heatid="19490" lane="2" entrytime="00:02:41.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.78" />
                    <SPLIT distance="100" swimtime="00:01:16.15" />
                    <SPLIT distance="150" swimtime="00:01:57.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="294" reactiontime="+74" swimtime="00:00:37.95" resultid="17958" heatid="19553" lane="5" entrytime="00:00:37.09" entrycourse="SCM" />
                <RESULT eventid="1744" points="217" reactiontime="+58" swimtime="00:05:53.17" resultid="17959" heatid="19702" lane="6" entrytime="00:06:07.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                    <SPLIT distance="100" swimtime="00:01:18.99" />
                    <SPLIT distance="150" swimtime="00:02:03.21" />
                    <SPLIT distance="200" swimtime="00:02:48.32" />
                    <SPLIT distance="250" swimtime="00:03:34.15" />
                    <SPLIT distance="300" swimtime="00:04:21.50" />
                    <SPLIT distance="350" swimtime="00:05:08.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-06-14" firstname="Kinga" gender="F" lastname="Maciupa" nation="POL" athleteid="17940">
              <RESULTS>
                <RESULT eventid="1096" points="484" reactiontime="+67" swimtime="00:02:35.11" resultid="17941" heatid="19309" lane="8" entrytime="00:02:40.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                    <SPLIT distance="100" swimtime="00:01:12.47" />
                    <SPLIT distance="150" swimtime="00:01:57.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="477" reactiontime="+78" swimtime="00:00:32.85" resultid="17942" heatid="19341" lane="0" entrytime="00:00:33.12" entrycourse="SCM" />
                <RESULT eventid="14225" points="497" reactiontime="+72" swimtime="00:01:11.50" resultid="17943" heatid="19395" lane="5" entrytime="00:01:13.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="434" reactiontime="+76" swimtime="00:00:32.20" resultid="17944" heatid="19449" lane="0" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1555" points="466" reactiontime="+78" swimtime="00:05:34.43" resultid="17945" heatid="19505" lane="2" entrytime="00:05:40.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.96" />
                    <SPLIT distance="100" swimtime="00:01:13.96" />
                    <SPLIT distance="150" swimtime="00:01:56.89" />
                    <SPLIT distance="200" swimtime="00:02:38.74" />
                    <SPLIT distance="250" swimtime="00:03:25.46" />
                    <SPLIT distance="300" swimtime="00:04:13.75" />
                    <SPLIT distance="350" swimtime="00:04:55.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="424" reactiontime="+82" swimtime="00:01:12.67" resultid="17946" heatid="19515" lane="3" entrytime="00:01:11.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-20" firstname="Agnieszka" gender="F" lastname="Krzyżostaniak" nation="POL" athleteid="17901">
              <RESULTS>
                <RESULT eventid="1062" points="543" reactiontime="+85" swimtime="00:00:28.48" resultid="17902" heatid="19283" lane="7" entrytime="00:00:28.00" entrycourse="SCM" />
                <RESULT eventid="1187" points="553" reactiontime="+76" swimtime="00:00:31.27" resultid="17903" heatid="19341" lane="5" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="14225" points="482" reactiontime="+82" swimtime="00:01:12.25" resultid="17904" heatid="19396" lane="9" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" status="DNS" swimtime="00:00:00.00" resultid="17905" heatid="19448" lane="0" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1457" points="484" reactiontime="+70" swimtime="00:01:10.06" resultid="17906" heatid="19469" lane="6" entrytime="00:01:09.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="391" reactiontime="+86" swimtime="00:00:39.16" resultid="17907" heatid="19543" lane="4" entrytime="00:00:40.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-18" firstname="Jan" gender="M" lastname="Roenig" nation="POL" athleteid="17908">
              <RESULTS>
                <RESULT eventid="1079" points="426" reactiontime="+90" swimtime="00:00:26.92" resultid="17909" heatid="19295" lane="5" entrytime="00:00:29.00" entrycourse="SCM" />
                <RESULT eventid="1273" points="387" reactiontime="+80" swimtime="00:01:01.65" resultid="17910" heatid="19383" lane="9" entrytime="00:01:03.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="389" reactiontime="+94" swimtime="00:01:16.12" resultid="17911" heatid="19439" lane="1" entrytime="00:01:22.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="369" reactiontime="+85" swimtime="00:00:30.39" resultid="17912" heatid="19454" lane="4" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1681" points="430" reactiontime="+76" swimtime="00:00:33.45" resultid="17913" heatid="19557" lane="9" entrytime="00:00:34.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-28" firstname="Tomasz" gender="M" lastname="Panasiuk" nation="POL" athleteid="17922">
              <RESULTS>
                <RESULT eventid="1273" points="125" reactiontime="+92" swimtime="00:01:29.78" resultid="17923" heatid="19374" lane="2" entrytime="00:01:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="95" reactiontime="+93" swimtime="00:01:49.98" resultid="17924" heatid="19398" lane="2" entrytime="00:01:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="17925" heatid="19451" lane="1" entrytime="00:00:55.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="SMT SZCZECIN 1" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="332" reactiontime="+74" swimtime="00:02:10.66" resultid="18016" heatid="19422" lane="4" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                    <SPLIT distance="100" swimtime="00:01:14.54" />
                    <SPLIT distance="150" swimtime="00:01:42.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17934" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="18000" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="17914" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="17973" number="4" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="422" reactiontime="+82" swimtime="00:01:50.07" resultid="18017" heatid="19501" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.84" />
                    <SPLIT distance="100" swimtime="00:00:55.07" />
                    <SPLIT distance="150" swimtime="00:01:25.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17908" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="17973" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="18000" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="17914" number="4" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="SMT SZCZECIN 2" number="2">
              <RESULTS>
                <RESULT eventid="1381" points="100" reactiontime="+105" swimtime="00:03:14.79" resultid="18018" heatid="19421" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.89" />
                    <SPLIT distance="100" swimtime="00:01:57.01" />
                    <SPLIT distance="150" swimtime="00:02:42.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18005" number="1" reactiontime="+105" />
                    <RELAYPOSITION athleteid="17993" number="2" reactiontime="+90" />
                    <RELAYPOSITION athleteid="17922" number="3" reactiontime="+81" />
                    <RELAYPOSITION athleteid="17982" number="4" reactiontime="+63" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="159" reactiontime="+74" swimtime="00:02:32.36" resultid="18019" heatid="19499" lane="3" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.35" />
                    <SPLIT distance="100" swimtime="00:01:07.57" />
                    <SPLIT distance="150" swimtime="00:01:42.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17952" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="17993" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="17969" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="18005" number="4" reactiontime="+78" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" name="SMT SZCZECIN 3" number="3">
              <RESULTS>
                <RESULT eventid="1548" points="245" reactiontime="+78" swimtime="00:02:11.97" resultid="18020" heatid="19499" lane="4" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.18" />
                    <SPLIT distance="100" swimtime="00:01:11.21" />
                    <SPLIT distance="150" swimtime="00:01:39.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17996" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="17967" number="2" reactiontime="+63" />
                    <RELAYPOSITION athleteid="17988" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="17934" number="4" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" name="SMT SZCZECIN 1" number="1">
              <RESULTS>
                <RESULT eventid="1358" points="453" reactiontime="+76" swimtime="00:02:14.42" resultid="18014" heatid="19420" lane="2" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                    <SPLIT distance="100" swimtime="00:01:11.83" />
                    <SPLIT distance="150" swimtime="00:01:44.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17901" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="17947" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="17940" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="17926" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1525" status="DNS" swimtime="00:00:00.00" resultid="18015" heatid="19498" lane="2" entrytime="00:02:06.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17926" number="1" />
                    <RELAYPOSITION athleteid="17940" number="2" />
                    <RELAYPOSITION athleteid="17960" number="3" />
                    <RELAYPOSITION athleteid="17901" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="SMT SZCZECIN 1" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="444" reactiontime="+87" swimtime="00:01:56.03" resultid="18010" heatid="19321" lane="5" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.08" />
                    <SPLIT distance="100" swimtime="00:00:59.90" />
                    <SPLIT distance="150" swimtime="00:01:31.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17908" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="17960" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="17926" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="17914" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="493" reactiontime="+74" swimtime="00:02:02.97" resultid="18011" heatid="19563" lane="4" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                    <SPLIT distance="100" swimtime="00:01:04.68" />
                    <SPLIT distance="150" swimtime="00:01:37.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17901" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="17908" number="2" reactiontime="+69" />
                    <RELAYPOSITION athleteid="17926" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="17914" number="4" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="SMT SZCZECIN 2" number="2">
              <RESULTS>
                <RESULT eventid="1130" points="432" reactiontime="+73" swimtime="00:01:57.15" resultid="18012" heatid="19321" lane="4" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.80" />
                    <SPLIT distance="100" swimtime="00:00:59.23" />
                    <SPLIT distance="150" swimtime="00:01:29.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17952" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="17940" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="18000" number="3" reactiontime="+72" />
                    <RELAYPOSITION athleteid="17901" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" name="SMT SZCZECIN 2" number="2">
              <RESULTS>
                <RESULT eventid="1698" status="DNS" swimtime="00:00:00.00" resultid="18013" heatid="19563" lane="2" entrytime="00:02:20.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17934" number="1" />
                    <RELAYPOSITION athleteid="17901" number="2" />
                    <RELAYPOSITION athleteid="17988" number="3" />
                    <RELAYPOSITION athleteid="17940" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="15734" name="T.P.Masters Opole">
          <CONTACT city="OPOLE" name="KRASNODĘBSKI" />
          <ATHLETES>
            <ATHLETE birthdate="1988-01-01" firstname="Tomasz" gender="M" lastname="Samsel" nation="POL" athleteid="15747">
              <RESULTS>
                <RESULT eventid="1079" points="496" reactiontime="+74" swimtime="00:00:25.58" resultid="15748" heatid="19301" lane="4" entrytime="00:00:25.98" />
                <RESULT eventid="1113" points="409" reactiontime="+78" swimtime="00:02:27.69" resultid="15749" heatid="19314" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                    <SPLIT distance="100" swimtime="00:01:09.62" />
                    <SPLIT distance="150" swimtime="00:01:53.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="516" reactiontime="+72" swimtime="00:00:56.00" resultid="15750" heatid="19386" lane="7" entrytime="00:00:57.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="426" reactiontime="+73" swimtime="00:01:06.83" resultid="15751" heatid="19407" lane="8" entrytime="00:01:08.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="475" reactiontime="+84" swimtime="00:02:07.31" resultid="15752" heatid="19495" lane="1" entrytime="00:02:08.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.01" />
                    <SPLIT distance="100" swimtime="00:01:01.57" />
                    <SPLIT distance="150" swimtime="00:01:34.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="333" reactiontime="+80" swimtime="00:01:09.31" resultid="15753" heatid="19522" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="373" reactiontime="+82" swimtime="00:00:35.07" resultid="15754" heatid="19552" lane="0" entrytime="00:00:39.49" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-01" firstname="Grzegorz" gender="M" lastname="Radomski" nation="POL" athleteid="15755">
              <RESULTS>
                <RESULT eventid="1113" points="529" reactiontime="+79" swimtime="00:02:15.54" resultid="15756" heatid="19317" lane="2" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.52" />
                    <SPLIT distance="100" swimtime="00:01:02.67" />
                    <SPLIT distance="150" swimtime="00:01:41.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14189" points="468" reactiontime="+76" swimtime="00:09:30.79" resultid="15757" heatid="19617" lane="7" entrytime="00:10:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                    <SPLIT distance="100" swimtime="00:01:04.31" />
                    <SPLIT distance="150" swimtime="00:01:39.78" />
                    <SPLIT distance="200" swimtime="00:02:15.35" />
                    <SPLIT distance="250" swimtime="00:02:51.12" />
                    <SPLIT distance="300" swimtime="00:03:26.86" />
                    <SPLIT distance="350" swimtime="00:04:03.26" />
                    <SPLIT distance="400" swimtime="00:04:39.74" />
                    <SPLIT distance="450" swimtime="00:05:16.08" />
                    <SPLIT distance="500" swimtime="00:05:52.57" />
                    <SPLIT distance="550" swimtime="00:06:29.58" />
                    <SPLIT distance="600" swimtime="00:07:05.97" />
                    <SPLIT distance="650" swimtime="00:07:42.31" />
                    <SPLIT distance="700" swimtime="00:08:19.27" />
                    <SPLIT distance="750" swimtime="00:08:56.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-01" firstname="Agnieszka" gender="F" lastname="Bartnikowska" nation="POL" athleteid="15735">
              <RESULTS>
                <RESULT eventid="1423" points="487" reactiontime="+82" swimtime="00:00:30.98" resultid="15736" heatid="19444" lane="6" />
                <RESULT eventid="1457" points="481" reactiontime="+76" swimtime="00:01:10.23" resultid="15737" heatid="19469" lane="9" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="465" reactiontime="+89" swimtime="00:02:33.83" resultid="15738" heatid="19529" lane="6" entrytime="00:02:36.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                    <SPLIT distance="100" swimtime="00:01:15.90" />
                    <SPLIT distance="150" swimtime="00:01:55.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-01-01" firstname="Tadeusz" gender="M" lastname="Witkowski" nation="POL" athleteid="15761">
              <RESULTS>
                <RESULT eventid="1079" points="89" reactiontime="+126" swimtime="00:00:45.31" resultid="15762" heatid="19285" lane="3" entrytime="00:00:42.00" />
                <RESULT eventid="1205" points="48" reactiontime="+95" swimtime="00:01:00.83" resultid="15763" heatid="19343" lane="2" entrytime="00:00:59.00" />
                <RESULT eventid="1273" points="66" reactiontime="+129" swimtime="00:01:50.86" resultid="15764" heatid="19374" lane="3" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="39" reactiontime="+90" swimtime="00:02:23.38" resultid="15765" heatid="19471" lane="9" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="15766" heatid="19486" lane="5" entrytime="00:04:00.00" />
                <RESULT eventid="1647" points="34" reactiontime="+98" swimtime="00:05:23.69" resultid="15767" heatid="19532" lane="1" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.37" />
                    <SPLIT distance="100" swimtime="00:02:37.13" />
                    <SPLIT distance="150" swimtime="00:04:01.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="73" reactiontime="+121" swimtime="00:01:00.39" resultid="15768" heatid="19547" lane="5" entrytime="00:00:59.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-01" firstname="Oskar" gender="M" lastname="Orski" nation="POL" athleteid="15758">
              <RESULTS>
                <RESULT eventid="1273" points="285" reactiontime="+98" swimtime="00:01:08.26" resultid="15759" heatid="19380" lane="4" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="251" reactiontime="+107" swimtime="00:01:28.14" resultid="15760" heatid="19437" lane="3" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-01" firstname="Zbigniew" gender="M" lastname="Januszkiewicz" nation="POL" athleteid="15739">
              <RESULTS>
                <RESULT eventid="1079" points="423" reactiontime="+75" swimtime="00:00:26.97" resultid="15740" heatid="19298" lane="9" entrytime="00:00:27.80" />
                <RESULT eventid="1113" points="402" reactiontime="+77" swimtime="00:02:28.47" resultid="15741" heatid="19316" lane="9" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.03" />
                    <SPLIT distance="100" swimtime="00:01:08.45" />
                    <SPLIT distance="150" swimtime="00:01:54.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="368" reactiontime="+71" swimtime="00:00:30.99" resultid="15742" heatid="19351" lane="2" entrytime="00:00:30.90" />
                <RESULT eventid="1341" points="338" reactiontime="+88" swimtime="00:02:35.72" resultid="15743" heatid="19417" lane="0" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.71" />
                    <SPLIT distance="100" swimtime="00:01:13.58" />
                    <SPLIT distance="150" swimtime="00:01:53.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="426" reactiontime="+84" swimtime="00:00:28.95" resultid="15744" heatid="19450" lane="3" />
                <RESULT eventid="1474" points="419" reactiontime="+75" swimtime="00:01:05.36" resultid="15745" heatid="19477" lane="3" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.91" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Europy Masters" eventid="1647" points="417" reactiontime="+62" swimtime="00:02:21.37" resultid="15746" heatid="19537" lane="7" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.18" />
                    <SPLIT distance="100" swimtime="00:01:09.32" />
                    <SPLIT distance="150" swimtime="00:01:45.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="SVK" clubid="14747" name="THREE POOLS Bernolákovo">
          <ATHLETES>
            <ATHLETE birthdate="1957-07-19" firstname="Jozef" gender="M" lastname="Krčík" nation="SVK" athleteid="14748">
              <RESULTS>
                <RESULT eventid="14207" points="303" reactiontime="+118" swimtime="00:21:01.85" resultid="14749" heatid="19621" lane="4" entrytime="00:23:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.22" />
                    <SPLIT distance="100" swimtime="00:01:19.14" />
                    <SPLIT distance="150" swimtime="00:02:01.58" />
                    <SPLIT distance="200" swimtime="00:02:44.21" />
                    <SPLIT distance="250" swimtime="00:03:26.57" />
                    <SPLIT distance="300" swimtime="00:04:08.75" />
                    <SPLIT distance="350" swimtime="00:04:50.66" />
                    <SPLIT distance="400" swimtime="00:05:32.71" />
                    <SPLIT distance="450" swimtime="00:06:14.55" />
                    <SPLIT distance="500" swimtime="00:07:38.57" />
                    <SPLIT distance="550" swimtime="00:08:20.54" />
                    <SPLIT distance="600" swimtime="00:09:02.73" />
                    <SPLIT distance="650" swimtime="00:09:44.74" />
                    <SPLIT distance="700" swimtime="00:10:26.36" />
                    <SPLIT distance="750" swimtime="00:11:08.44" />
                    <SPLIT distance="800" swimtime="00:11:50.84" />
                    <SPLIT distance="850" swimtime="00:12:32.85" />
                    <SPLIT distance="950" swimtime="00:13:15.39" />
                    <SPLIT distance="1000" swimtime="00:13:57.63" />
                    <SPLIT distance="1050" swimtime="00:14:40.02" />
                    <SPLIT distance="1100" swimtime="00:15:22.15" />
                    <SPLIT distance="1150" swimtime="00:16:04.61" />
                    <SPLIT distance="1200" swimtime="00:16:46.79" />
                    <SPLIT distance="1250" swimtime="00:17:29.46" />
                    <SPLIT distance="1300" swimtime="00:18:12.36" />
                    <SPLIT distance="1350" swimtime="00:18:55.07" />
                    <SPLIT distance="1400" swimtime="00:19:37.49" />
                    <SPLIT distance="1450" swimtime="00:20:19.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="224" reactiontime="+112" swimtime="00:01:22.82" resultid="14750" heatid="19400" lane="5" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="262" reactiontime="+102" swimtime="00:02:35.21" resultid="14751" heatid="19490" lane="0" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.73" />
                    <SPLIT distance="100" swimtime="00:01:15.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="279" reactiontime="+109" swimtime="00:05:24.76" resultid="14752" heatid="19703" lane="3" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                    <SPLIT distance="100" swimtime="00:01:18.21" />
                    <SPLIT distance="150" swimtime="00:01:58.53" />
                    <SPLIT distance="200" swimtime="00:02:40.05" />
                    <SPLIT distance="250" swimtime="00:03:21.52" />
                    <SPLIT distance="300" swimtime="00:04:02.92" />
                    <SPLIT distance="350" swimtime="00:04:44.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="CZE" clubid="18532" name="TJ Alcedo Vsetín">
          <CONTACT city="Vsetín" email="pavel.obr@czechswimming.cz" name="Pavel Obr" state="CZE" street="Dolní Jasenka 770" zip="75501" />
          <ATHLETES>
            <ATHLETE birthdate="1967-05-03" firstname="Pavel" gender="M" lastname="Obr" nation="CZE" athleteid="18533">
              <RESULTS>
                <RESULT eventid="1079" points="361" reactiontime="+81" swimtime="00:00:28.45" resultid="18534" heatid="19298" lane="6" entrytime="00:00:27.50" />
                <RESULT eventid="1113" points="343" reactiontime="+81" swimtime="00:02:36.50" resultid="18535" heatid="19315" lane="9" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                    <SPLIT distance="100" swimtime="00:01:13.58" />
                    <SPLIT distance="150" swimtime="00:01:58.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="423" reactiontime="+82" swimtime="00:00:59.84" resultid="18536" heatid="19383" lane="5" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.67" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K16 - Niejednoczesne dotknięcie ściany dłońmi przy nawrocie lub na zakończenie wyścigu (Time: 12:03)" eventid="14243" reactiontime="+84" status="DSQ" swimtime="00:01:09.75" resultid="18537" heatid="19405" lane="3" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="387" reactiontime="+91" swimtime="00:00:29.91" resultid="18538" heatid="19459" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1578" points="262" reactiontime="+93" swimtime="00:06:07.90" resultid="18539" heatid="19510" lane="1" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                    <SPLIT distance="100" swimtime="00:01:12.01" />
                    <SPLIT distance="150" swimtime="00:01:59.91" />
                    <SPLIT distance="200" swimtime="00:02:48.56" />
                    <SPLIT distance="250" swimtime="00:03:40.98" />
                    <SPLIT distance="300" swimtime="00:04:36.74" />
                    <SPLIT distance="350" swimtime="00:05:21.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="372" reactiontime="+91" swimtime="00:00:35.10" resultid="18540" heatid="19556" lane="1" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="020/16" nation="POL" region="ZAC" clubid="17755" name="TKKF Koszalin Masters">
          <CONTACT city="Koszalin" email="jakubkielar3@gmail.com" internet="www.masterskoszalin.pl" name="Kielar" phone="693193137" />
          <ATHLETES>
            <ATHLETE birthdate="1995-01-01" firstname="Kamil" gender="M" lastname="Mika" nation="POL" athleteid="17842">
              <RESULTS>
                <RESULT eventid="14243" points="381" reactiontime="+90" swimtime="00:01:09.35" resultid="17843" heatid="19404" lane="6" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="444" reactiontime="+79" swimtime="00:01:12.85" resultid="17844" heatid="19442" lane="9" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="446" reactiontime="+82" swimtime="00:00:33.04" resultid="17845" heatid="19558" lane="5" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-03-14" firstname="Sylwia" gender="F" lastname="Kuśpiet" nation="POL" athleteid="17853">
              <RESULTS>
                <RESULT eventid="1062" points="480" swimtime="00:00:29.67" resultid="17854" heatid="19283" lane="9" entrytime="00:00:29.00" />
                <RESULT eventid="14225" points="507" reactiontime="+94" swimtime="00:01:11.05" resultid="17855" heatid="19396" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="453" reactiontime="+84" swimtime="00:00:31.74" resultid="17856" heatid="19449" lane="8" entrytime="00:00:32.00" />
                <RESULT eventid="1664" points="423" reactiontime="+89" swimtime="00:00:38.14" resultid="17857" heatid="19543" lane="3" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-02-20" firstname="Artur" gender="M" lastname="Rutkowski" nation="POL" athleteid="17791">
              <RESULTS>
                <RESULT eventid="1113" points="309" reactiontime="+91" swimtime="00:02:42.15" resultid="17792" heatid="19314" lane="0" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.22" />
                    <SPLIT distance="100" swimtime="00:01:16.98" />
                    <SPLIT distance="150" swimtime="00:02:04.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="234" reactiontime="+75" swimtime="00:00:36.01" resultid="17793" heatid="19348" lane="1" entrytime="00:00:36.00" />
                <RESULT eventid="1341" points="255" reactiontime="+91" swimtime="00:02:51.00" resultid="17794" heatid="19416" lane="6" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                    <SPLIT distance="100" swimtime="00:01:17.61" />
                    <SPLIT distance="150" swimtime="00:02:02.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="333" reactiontime="+87" swimtime="00:00:31.44" resultid="17795" heatid="19456" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1578" points="278" reactiontime="+94" swimtime="00:06:00.44" resultid="17796" heatid="19509" lane="3" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.04" />
                    <SPLIT distance="100" swimtime="00:01:22.54" />
                    <SPLIT distance="150" swimtime="00:02:09.44" />
                    <SPLIT distance="200" swimtime="00:02:56.68" />
                    <SPLIT distance="250" swimtime="00:03:46.99" />
                    <SPLIT distance="300" swimtime="00:04:39.22" />
                    <SPLIT distance="350" swimtime="00:05:21.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="292" reactiontime="+89" swimtime="00:01:12.44" resultid="17797" heatid="19521" lane="7" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="315" reactiontime="+94" swimtime="00:00:37.11" resultid="17798" heatid="19554" lane="1" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-08-26" firstname="Dorota" gender="F" lastname="Gudaniec" nation="POL" athleteid="17812">
              <RESULTS>
                <RESULT eventid="1165" points="235" reactiontime="+106" swimtime="00:24:50.25" resultid="17813" heatid="19624" lane="3" entrytime="00:24:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.64" />
                    <SPLIT distance="100" swimtime="00:01:30.40" />
                    <SPLIT distance="150" swimtime="00:02:19.83" />
                    <SPLIT distance="200" swimtime="00:03:09.32" />
                    <SPLIT distance="250" swimtime="00:03:59.22" />
                    <SPLIT distance="300" swimtime="00:04:49.11" />
                    <SPLIT distance="350" swimtime="00:05:39.43" />
                    <SPLIT distance="400" swimtime="00:06:29.21" />
                    <SPLIT distance="450" swimtime="00:07:19.30" />
                    <SPLIT distance="500" swimtime="00:08:09.44" />
                    <SPLIT distance="550" swimtime="00:08:59.28" />
                    <SPLIT distance="600" swimtime="00:09:49.64" />
                    <SPLIT distance="650" swimtime="00:10:40.03" />
                    <SPLIT distance="700" swimtime="00:11:29.82" />
                    <SPLIT distance="750" swimtime="00:12:19.98" />
                    <SPLIT distance="800" swimtime="00:13:10.12" />
                    <SPLIT distance="850" swimtime="00:14:00.28" />
                    <SPLIT distance="900" swimtime="00:14:50.23" />
                    <SPLIT distance="950" swimtime="00:15:40.50" />
                    <SPLIT distance="1000" swimtime="00:16:30.50" />
                    <SPLIT distance="1050" swimtime="00:17:20.70" />
                    <SPLIT distance="1100" swimtime="00:18:10.86" />
                    <SPLIT distance="1150" swimtime="00:19:01.08" />
                    <SPLIT distance="1200" swimtime="00:19:51.35" />
                    <SPLIT distance="1250" swimtime="00:20:41.53" />
                    <SPLIT distance="1300" swimtime="00:21:31.94" />
                    <SPLIT distance="1350" swimtime="00:22:22.65" />
                    <SPLIT distance="1400" swimtime="00:23:12.76" />
                    <SPLIT distance="1450" swimtime="00:24:02.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="182" reactiontime="+107" swimtime="00:03:57.25" resultid="17814" heatid="19356" lane="6" entrytime="00:03:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.48" />
                    <SPLIT distance="100" swimtime="00:01:52.44" />
                    <SPLIT distance="150" swimtime="00:02:55.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="194" reactiontime="+107" swimtime="00:01:37.78" resultid="17815" heatid="19391" lane="2" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="178" reactiontime="+113" swimtime="00:01:50.76" resultid="17816" heatid="19429" lane="1" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="198" reactiontime="+109" swimtime="00:07:25.01" resultid="17817" heatid="19504" lane="0" entrytime="00:07:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.77" />
                    <SPLIT distance="100" swimtime="00:01:48.69" />
                    <SPLIT distance="150" swimtime="00:02:46.09" />
                    <SPLIT distance="200" swimtime="00:03:41.46" />
                    <SPLIT distance="250" swimtime="00:04:42.79" />
                    <SPLIT distance="300" swimtime="00:05:45.39" />
                    <SPLIT distance="350" swimtime="00:06:35.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="175" reactiontime="+83" swimtime="00:03:32.83" resultid="17818" heatid="19527" lane="2" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.67" />
                    <SPLIT distance="100" swimtime="00:01:45.20" />
                    <SPLIT distance="150" swimtime="00:02:40.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="218" reactiontime="+99" swimtime="00:06:29.22" resultid="17819" heatid="19696" lane="5" entrytime="00:06:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.69" />
                    <SPLIT distance="100" swimtime="00:01:30.34" />
                    <SPLIT distance="150" swimtime="00:02:19.81" />
                    <SPLIT distance="200" swimtime="00:03:09.28" />
                    <SPLIT distance="250" swimtime="00:03:59.50" />
                    <SPLIT distance="300" swimtime="00:04:49.83" />
                    <SPLIT distance="350" swimtime="00:05:40.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-03-29" firstname="Marcin" gender="M" lastname="Jaworski" nation="POL" athleteid="17833">
              <RESULTS>
                <RESULT eventid="1079" points="270" reactiontime="+95" swimtime="00:00:31.31" resultid="17834" heatid="19295" lane="7" entrytime="00:00:29.00" />
                <RESULT eventid="1205" points="230" reactiontime="+95" swimtime="00:00:36.23" resultid="17835" heatid="19347" lane="3" entrytime="00:00:37.00" />
                <RESULT eventid="1474" points="247" reactiontime="+81" swimtime="00:01:17.88" resultid="17836" heatid="19474" lane="7" entrytime="00:01:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-03-24" firstname="Radosław" gender="M" lastname="Bor" nation="POL" athleteid="17828">
              <RESULTS>
                <RESULT eventid="1079" points="539" reactiontime="+76" swimtime="00:00:24.88" resultid="17829" heatid="19304" lane="0" entrytime="00:00:24.00" />
                <RESULT eventid="1205" points="420" reactiontime="+74" swimtime="00:00:29.65" resultid="17830" heatid="19353" lane="8" entrytime="00:00:28.00" />
                <RESULT eventid="1273" points="589" reactiontime="+76" swimtime="00:00:53.60" resultid="17831" heatid="19388" lane="2" entrytime="00:00:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="445" reactiontime="+78" swimtime="00:01:04.03" resultid="17832" heatid="19477" lane="0" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-11-19" firstname="Małgorzata" gender="F" lastname="Milczarek" nation="POL" athleteid="17850">
              <RESULTS>
                <RESULT eventid="1062" points="133" reactiontime="+94" swimtime="00:00:45.44" resultid="17851" heatid="19276" lane="7" entrytime="00:00:50.00" />
                <RESULT eventid="1664" points="191" reactiontime="+75" swimtime="00:00:49.67" resultid="17852" heatid="19541" lane="9" entrytime="00:00:49.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-08-22" firstname="Grzegorz" gender="M" lastname="Ćwikła" nation="POL" athleteid="17756">
              <RESULTS>
                <RESULT eventid="1113" points="293" reactiontime="+86" swimtime="00:02:44.92" resultid="17757" heatid="19313" lane="2" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                    <SPLIT distance="100" swimtime="00:01:20.55" />
                    <SPLIT distance="150" swimtime="00:02:09.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14207" points="280" reactiontime="+86" swimtime="00:21:35.11" resultid="17758" heatid="19622" lane="1" entrytime="00:22:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.07" />
                    <SPLIT distance="100" swimtime="00:01:16.76" />
                    <SPLIT distance="150" swimtime="00:01:59.20" />
                    <SPLIT distance="200" swimtime="00:02:42.24" />
                    <SPLIT distance="250" swimtime="00:03:25.51" />
                    <SPLIT distance="300" swimtime="00:04:08.51" />
                    <SPLIT distance="350" swimtime="00:04:52.13" />
                    <SPLIT distance="400" swimtime="00:05:35.26" />
                    <SPLIT distance="450" swimtime="00:06:19.06" />
                    <SPLIT distance="500" swimtime="00:07:02.61" />
                    <SPLIT distance="550" swimtime="00:07:46.26" />
                    <SPLIT distance="600" swimtime="00:08:30.02" />
                    <SPLIT distance="650" swimtime="00:09:13.48" />
                    <SPLIT distance="700" swimtime="00:09:57.18" />
                    <SPLIT distance="750" swimtime="00:10:41.09" />
                    <SPLIT distance="800" swimtime="00:11:24.84" />
                    <SPLIT distance="850" swimtime="00:12:08.40" />
                    <SPLIT distance="900" swimtime="00:12:52.46" />
                    <SPLIT distance="950" swimtime="00:13:37.09" />
                    <SPLIT distance="1000" swimtime="00:14:21.33" />
                    <SPLIT distance="1050" swimtime="00:15:05.53" />
                    <SPLIT distance="1100" swimtime="00:15:49.93" />
                    <SPLIT distance="1150" swimtime="00:16:34.19" />
                    <SPLIT distance="1200" swimtime="00:17:18.67" />
                    <SPLIT distance="1250" swimtime="00:18:03.31" />
                    <SPLIT distance="1300" swimtime="00:18:47.03" />
                    <SPLIT distance="1350" swimtime="00:19:30.60" />
                    <SPLIT distance="1400" swimtime="00:20:13.35" />
                    <SPLIT distance="1450" swimtime="00:20:56.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="279" reactiontime="+74" swimtime="00:00:33.99" resultid="17759" heatid="19348" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="14243" points="294" reactiontime="+77" swimtime="00:01:15.59" resultid="17760" heatid="19404" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="281" reactiontime="+70" swimtime="00:01:14.63" resultid="17761" heatid="19475" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="271" reactiontime="+88" swimtime="00:06:03.63" resultid="17762" heatid="19509" lane="6" entrytime="00:06:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.52" />
                    <SPLIT distance="100" swimtime="00:01:24.43" />
                    <SPLIT distance="150" swimtime="00:02:13.46" />
                    <SPLIT distance="200" swimtime="00:03:01.03" />
                    <SPLIT distance="250" swimtime="00:03:53.81" />
                    <SPLIT distance="300" swimtime="00:04:46.12" />
                    <SPLIT distance="350" swimtime="00:05:25.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="233" reactiontime="+71" swimtime="00:02:51.65" resultid="17763" heatid="19535" lane="7" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.07" />
                    <SPLIT distance="100" swimtime="00:01:22.98" />
                    <SPLIT distance="150" swimtime="00:02:08.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="296" reactiontime="+89" swimtime="00:05:18.44" resultid="17764" heatid="19705" lane="2" entrytime="00:05:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                    <SPLIT distance="100" swimtime="00:01:14.94" />
                    <SPLIT distance="150" swimtime="00:01:56.10" />
                    <SPLIT distance="200" swimtime="00:02:37.71" />
                    <SPLIT distance="250" swimtime="00:03:19.39" />
                    <SPLIT distance="300" swimtime="00:04:00.86" />
                    <SPLIT distance="350" swimtime="00:04:41.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-02-24" firstname="Wioletta" gender="F" lastname="Pawliczek" nation="POL" athleteid="17799">
              <RESULTS>
                <RESULT eventid="1062" points="293" reactiontime="+85" swimtime="00:00:34.99" resultid="17800" heatid="19279" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1187" points="261" reactiontime="+76" swimtime="00:00:40.16" resultid="17801" heatid="19339" lane="7" entrytime="00:00:39.00" />
                <RESULT eventid="1256" points="277" swimtime="00:01:18.08" resultid="17802" heatid="19370" lane="0" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="255" reactiontime="+71" swimtime="00:01:26.75" resultid="17803" heatid="19467" lane="7" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="241" reactiontime="+77" swimtime="00:03:11.56" resultid="17804" heatid="19528" lane="0" entrytime="00:03:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.85" />
                    <SPLIT distance="100" swimtime="00:01:33.70" />
                    <SPLIT distance="150" swimtime="00:02:24.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Łukasz" gender="M" lastname="Olszak" nation="POL" athleteid="17837">
              <RESULTS>
                <RESULT eventid="1079" points="541" reactiontime="+76" swimtime="00:00:24.85" resultid="17838" heatid="19304" lane="8" entrytime="00:00:24.00" />
                <RESULT eventid="1205" points="406" reactiontime="+67" swimtime="00:00:30.00" resultid="17839" heatid="19353" lane="1" entrytime="00:00:28.00" />
                <RESULT eventid="1273" points="525" reactiontime="+77" swimtime="00:00:55.68" resultid="17840" heatid="19388" lane="1" entrytime="00:00:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="406" reactiontime="+64" swimtime="00:01:06.06" resultid="17841" heatid="19477" lane="9" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Dawid" gender="M" lastname="Fremel" nation="POL" athleteid="17846">
              <RESULTS>
                <RESULT eventid="14243" points="533" reactiontime="+69" swimtime="00:01:02.00" resultid="17847" heatid="19409" lane="8" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="613" reactiontime="+70" swimtime="00:01:05.46" resultid="17848" heatid="19443" lane="8" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="608" reactiontime="+74" swimtime="00:00:29.80" resultid="17849" heatid="19560" lane="2" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-07-05" firstname="Krzysztof" gender="M" lastname="Stefański" nation="POL" athleteid="17861">
              <RESULTS>
                <RESULT eventid="1079" points="363" reactiontime="+79" swimtime="00:00:28.38" resultid="17862" heatid="19297" lane="2" entrytime="00:00:28.00" />
                <RESULT eventid="1273" points="331" reactiontime="+87" swimtime="00:01:04.92" resultid="17863" heatid="19382" lane="4" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" status="DNS" swimtime="00:00:00.00" resultid="17864" heatid="19403" lane="3" entrytime="00:01:16.00" />
                <RESULT eventid="1440" points="292" reactiontime="+88" swimtime="00:00:32.83" resultid="17865" heatid="19455" lane="2" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-06-28" firstname="Michał" gender="M" lastname="Pieślak" nation="POL" athleteid="17776">
              <RESULTS>
                <RESULT eventid="1079" points="382" reactiontime="+76" swimtime="00:00:27.92" resultid="17777" heatid="19297" lane="6" entrytime="00:00:28.00" />
                <RESULT eventid="1273" points="377" reactiontime="+88" swimtime="00:01:02.17" resultid="17778" heatid="19383" lane="2" entrytime="00:01:02.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" status="DNS" swimtime="00:00:00.00" resultid="17779" heatid="19404" lane="9" entrytime="00:01:15.00" />
                <RESULT eventid="1406" points="304" reactiontime="+78" swimtime="00:01:22.70" resultid="17780" heatid="19439" lane="7" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="17781" heatid="19492" lane="7" entrytime="00:02:25.00" />
                <RESULT eventid="1681" points="335" reactiontime="+75" swimtime="00:00:36.33" resultid="17782" heatid="19555" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="17783" heatid="19705" lane="5" entrytime="00:05:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-05" firstname="Agnieszka" gender="F" lastname="Paziewska" nation="POL" athleteid="17770">
              <RESULTS>
                <RESULT eventid="1062" points="326" reactiontime="+91" swimtime="00:00:33.74" resultid="17771" heatid="19281" lane="4" entrytime="00:00:31.90" />
                <RESULT eventid="1256" points="325" reactiontime="+90" swimtime="00:01:14.00" resultid="17772" heatid="19371" lane="7" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="218" reactiontime="+94" swimtime="00:01:43.61" resultid="17773" heatid="19429" lane="5" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="272" reactiontime="+100" swimtime="00:02:50.85" resultid="17774" heatid="19483" lane="1" entrytime="00:02:46.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.78" />
                    <SPLIT distance="100" swimtime="00:01:20.42" />
                    <SPLIT distance="150" swimtime="00:02:06.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="252" reactiontime="+94" swimtime="00:00:45.34" resultid="17775" heatid="19542" lane="5" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Krzysztof" gender="M" lastname="Wróbel" nation="POL" athleteid="17824">
              <RESULTS>
                <RESULT eventid="14243" points="483" reactiontime="+76" swimtime="00:01:04.07" resultid="17825" heatid="19408" lane="7" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="583" reactiontime="+79" swimtime="00:01:06.53" resultid="17826" heatid="19442" lane="4" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="563" reactiontime="+77" swimtime="00:00:30.57" resultid="17827" heatid="19559" lane="4" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-06-16" firstname="Marcin" gender="M" lastname="Horbacz" nation="POL" athleteid="17820">
              <RESULTS>
                <RESULT eventid="14243" points="478" reactiontime="+95" swimtime="00:01:04.30" resultid="17821" heatid="19409" lane="0" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="523" reactiontime="+75" swimtime="00:01:09.00" resultid="17822" heatid="19442" lane="7" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="520" reactiontime="+80" swimtime="00:00:31.39" resultid="17823" heatid="19559" lane="0" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-01-01" firstname="Patryk" gender="M" lastname="Marszałek" nation="POL" athleteid="17858">
              <RESULTS>
                <RESULT eventid="1079" points="389" reactiontime="+80" swimtime="00:00:27.74" resultid="17859" heatid="19297" lane="5" entrytime="00:00:28.00" />
                <RESULT eventid="1273" points="369" reactiontime="+82" swimtime="00:01:02.65" resultid="17860" heatid="19385" lane="4" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-04-29" firstname="Lidia" gender="F" lastname="Mikołajczyk" nation="POL" athleteid="17784">
              <RESULTS>
                <RESULT eventid="1096" points="398" reactiontime="+100" swimtime="00:02:45.63" resultid="17785" heatid="19308" lane="6" entrytime="00:02:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.33" />
                    <SPLIT distance="100" swimtime="00:01:17.97" />
                    <SPLIT distance="150" swimtime="00:02:05.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="371" reactiontime="+95" swimtime="00:03:07.26" resultid="17786" heatid="19358" lane="8" entrytime="00:03:09.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.11" />
                    <SPLIT distance="100" swimtime="00:01:29.65" />
                    <SPLIT distance="150" swimtime="00:02:19.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="401" reactiontime="+95" swimtime="00:01:16.82" resultid="17787" heatid="19394" lane="6" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="349" reactiontime="+99" swimtime="00:01:28.51" resultid="17788" heatid="19431" lane="5" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="342" reactiontime="+108" swimtime="00:06:10.71" resultid="17789" heatid="19504" lane="5" entrytime="00:06:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.57" />
                    <SPLIT distance="100" swimtime="00:01:27.92" />
                    <SPLIT distance="150" swimtime="00:02:15.77" />
                    <SPLIT distance="200" swimtime="00:03:02.29" />
                    <SPLIT distance="250" swimtime="00:03:53.59" />
                    <SPLIT distance="300" swimtime="00:04:45.80" />
                    <SPLIT distance="350" swimtime="00:05:30.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="392" reactiontime="+95" swimtime="00:00:39.10" resultid="17790" heatid="19543" lane="6" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-28" firstname="Roman" gender="M" lastname="Pieślak" nation="POL" athleteid="17805">
              <RESULTS>
                <RESULT eventid="1079" points="314" reactiontime="+81" swimtime="00:00:29.78" resultid="17806" heatid="19293" lane="2" entrytime="00:00:29.80" />
                <RESULT eventid="1239" points="279" reactiontime="+88" swimtime="00:03:04.24" resultid="17807" heatid="19362" lane="4" entrytime="00:03:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                    <SPLIT distance="100" swimtime="00:01:24.66" />
                    <SPLIT distance="150" swimtime="00:02:13.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="295" reactiontime="+89" swimtime="00:01:07.48" resultid="17808" heatid="19381" lane="1" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="313" reactiontime="+82" swimtime="00:01:21.87" resultid="17809" heatid="19439" lane="2" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="17810" heatid="19491" lane="0" entrytime="00:02:35.00" />
                <RESULT eventid="1681" points="312" reactiontime="+75" swimtime="00:00:37.21" resultid="17811" heatid="19554" lane="7" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="team1" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="333" reactiontime="+89" swimtime="00:02:10.56" resultid="17873" heatid="19423" lane="3" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.29" />
                    <SPLIT distance="100" swimtime="00:01:08.11" />
                    <SPLIT distance="150" swimtime="00:01:40.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17833" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="17824" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="17861" number="3" reactiontime="+29" />
                    <RELAYPOSITION athleteid="17805" number="4" reactiontime="+71" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="team1" number="1">
              <RESULTS>
                <RESULT eventid="1548" points="415" reactiontime="+78" swimtime="00:01:50.70" resultid="17876" heatid="19501" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.96" />
                    <SPLIT distance="100" swimtime="00:00:56.80" />
                    <SPLIT distance="150" swimtime="00:01:24.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17776" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="17756" number="2" reactiontime="+22" />
                    <RELAYPOSITION athleteid="17861" number="3" reactiontime="+17" />
                    <RELAYPOSITION athleteid="17820" number="4" reactiontime="+18" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="team2" number="2">
              <RESULTS>
                <RESULT eventid="1381" points="376" reactiontime="+67" swimtime="00:02:05.38" resultid="17874" heatid="19423" lane="7" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.70" />
                    <SPLIT distance="100" swimtime="00:01:06.32" />
                    <SPLIT distance="150" swimtime="00:01:37.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17756" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="17820" number="2" reactiontime="+21" />
                    <RELAYPOSITION athleteid="17791" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="17776" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="99" agetotalmin="80" gender="M" name="team2 kat 0" number="2">
              <RESULTS>
                <RESULT eventid="1548" status="DNS" swimtime="00:00:00.00" resultid="17877" heatid="19502" lane="4" entrytime="00:01:40.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17837" number="1" />
                    <RELAYPOSITION athleteid="17846" number="2" />
                    <RELAYPOSITION athleteid="17842" number="3" />
                    <RELAYPOSITION athleteid="17828" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="99" agetotalmin="80" gender="M" name="team3 kat 0" number="3">
              <RESULTS>
                <RESULT eventid="1381" points="499" reactiontime="+74" swimtime="00:01:54.04" resultid="17875" heatid="19424" lane="5" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.75" />
                    <SPLIT distance="100" swimtime="00:00:59.24" />
                    <SPLIT distance="150" swimtime="00:01:25.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17828" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="17846" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="17837" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="17842" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="team1" number="1">
              <RESULTS>
                <RESULT eventid="1358" points="391" reactiontime="+74" swimtime="00:02:21.19" resultid="17871" heatid="19420" lane="3" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                    <SPLIT distance="100" swimtime="00:01:18.05" />
                    <SPLIT distance="150" swimtime="00:01:48.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17799" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="17784" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="17853" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="17770" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1525" points="326" reactiontime="+106" swimtime="00:02:16.83" resultid="17872" heatid="19498" lane="6" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.57" />
                    <SPLIT distance="100" swimtime="00:01:12.88" />
                    <SPLIT distance="150" swimtime="00:01:43.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17853" number="1" reactiontime="+106" />
                    <RELAYPOSITION athleteid="17799" number="2" reactiontime="+3" />
                    <RELAYPOSITION athleteid="17784" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="17770" number="4" reactiontime="+10" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="team1" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="406" reactiontime="+92" swimtime="00:01:59.56" resultid="17866" heatid="19322" lane="8" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.55" />
                    <SPLIT distance="100" swimtime="00:01:03.68" />
                    <SPLIT distance="150" swimtime="00:01:31.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17784" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="17770" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="17861" number="3" reactiontime="+1" />
                    <RELAYPOSITION athleteid="17776" number="4" reactiontime="+51" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="team1" number="1">
              <RESULTS>
                <RESULT eventid="1698" points="404" reactiontime="+67" swimtime="00:02:11.35" resultid="17878" heatid="19564" lane="7" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.62" />
                    <SPLIT distance="150" swimtime="00:01:41.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17799" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="17824" number="2" />
                    <RELAYPOSITION athleteid="17853" number="3" />
                    <RELAYPOSITION athleteid="17805" number="4" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="team2" number="2">
              <RESULTS>
                <RESULT eventid="1130" status="DNS" swimtime="00:00:00.00" resultid="17867" heatid="19320" lane="5" entrytime="00:02:12.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17791" number="1" />
                    <RELAYPOSITION athleteid="17812" number="3" />
                    <RELAYPOSITION athleteid="17858" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="392" reactiontime="+77" swimtime="00:02:12.70" resultid="17868" heatid="19564" lane="0" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                    <SPLIT distance="100" swimtime="00:01:05.06" />
                    <SPLIT distance="150" swimtime="00:01:39.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17756" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="17820" number="2" reactiontime="+16" />
                    <RELAYPOSITION athleteid="17812" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="17770" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="team3" number="3">
              <RESULTS>
                <RESULT eventid="1130" points="366" reactiontime="+78" swimtime="00:02:03.77" resultid="17869" heatid="19321" lane="7" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                    <SPLIT distance="100" swimtime="00:01:04.75" />
                    <SPLIT distance="150" swimtime="00:01:34.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17756" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="17799" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="17853" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="17805" number="4" reactiontime="+51" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" status="DNS" swimtime="00:00:00.00" resultid="17870" heatid="19563" lane="0" entrytime="00:02:23.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17791" number="1" />
                    <RELAYPOSITION athleteid="17784" number="2" />
                    <RELAYPOSITION athleteid="17833" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="505815" nation="POL" region="WIE" clubid="15370" name="TMA BARRACUDA Kalisz">
          <CONTACT city="KALISZ" name="GALCZYNSKI WOJCIECH" phone="790690666" state="WLKP" zip="62-800" />
          <ATHLETES>
            <ATHLETE birthdate="1989-06-08" firstname="Mateusz" gender="M" lastname="Palczynski" nation="POL" athleteid="15386">
              <RESULTS>
                <RESULT eventid="1113" points="333" reactiontime="+89" swimtime="00:02:38.13" resultid="15387" heatid="19316" lane="0" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.67" />
                    <SPLIT distance="100" swimtime="00:01:14.52" />
                    <SPLIT distance="150" swimtime="00:01:58.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14189" reactiontime="+91" status="DNF" swimtime="00:00:00.00" resultid="15388" heatid="19617" lane="3" entrytime="00:10:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.90" />
                    <SPLIT distance="100" swimtime="00:01:16.68" />
                    <SPLIT distance="150" swimtime="00:01:58.60" />
                    <SPLIT distance="200" swimtime="00:02:42.61" />
                    <SPLIT distance="250" swimtime="00:03:28.91" />
                    <SPLIT distance="300" swimtime="00:04:15.86" />
                    <SPLIT distance="350" swimtime="00:05:03.39" />
                    <SPLIT distance="400" swimtime="00:05:51.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="321" reactiontime="+88" swimtime="00:02:55.74" resultid="15389" heatid="19364" lane="0" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                    <SPLIT distance="100" swimtime="00:01:20.76" />
                    <SPLIT distance="150" swimtime="00:02:07.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="247" reactiontime="+82" swimtime="00:02:52.87" resultid="15390" heatid="19417" lane="8" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                    <SPLIT distance="100" swimtime="00:01:16.38" />
                    <SPLIT distance="150" swimtime="00:02:04.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="405" reactiontime="+72" swimtime="00:01:15.11" resultid="15391" heatid="19442" lane="0" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="15392" heatid="19511" lane="9" entrytime="00:05:50.00" />
                <RESULT eventid="1647" points="278" reactiontime="+90" swimtime="00:02:41.77" resultid="15393" heatid="19535" lane="1" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.30" />
                    <SPLIT distance="150" swimtime="00:02:00.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="423" reactiontime="+80" swimtime="00:00:33.63" resultid="15394" heatid="19558" lane="7" entrytime="00:00:32.51" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-02-01" firstname="Andrzej" gender="M" lastname="Sypniewski" nation="POL" athleteid="15395">
              <RESULTS>
                <RESULT eventid="1079" points="259" reactiontime="+77" swimtime="00:00:31.75" resultid="15396" heatid="19289" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1113" points="231" reactiontime="+84" swimtime="00:02:58.52" resultid="15397" heatid="19312" lane="1" entrytime="00:03:06.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.84" />
                    <SPLIT distance="100" swimtime="00:01:23.76" />
                    <SPLIT distance="150" swimtime="00:02:14.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="224" reactiontime="+65" swimtime="00:03:18.03" resultid="15398" heatid="19362" lane="9" entrytime="00:03:16.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.73" />
                    <SPLIT distance="100" swimtime="00:01:32.87" />
                    <SPLIT distance="150" swimtime="00:02:25.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="247" reactiontime="+81" swimtime="00:01:20.07" resultid="15399" heatid="19402" lane="3" entrytime="00:01:18.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="244" reactiontime="+75" swimtime="00:01:28.91" resultid="15400" heatid="19437" lane="9" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="186" swimtime="00:01:25.63" resultid="15401" heatid="19474" lane="8" entrytime="00:01:25.78" />
                <RESULT eventid="1613" points="183" reactiontime="+75" swimtime="00:01:24.64" resultid="15402" heatid="19519" lane="8" entrytime="00:01:30.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="257" reactiontime="+76" swimtime="00:00:39.67" resultid="15403" heatid="19552" lane="8" entrytime="00:00:39.25" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-11" firstname="Patrycja" gender="F" lastname="Rupa" nation="POL" athleteid="15404">
              <RESULTS>
                <RESULT eventid="1096" status="DNS" swimtime="00:00:00.00" resultid="15405" heatid="19308" lane="1" entrytime="00:02:55.39" />
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="15406" heatid="19341" lane="7" entrytime="00:00:32.66" />
                <RESULT eventid="14225" status="DNS" swimtime="00:00:00.00" resultid="15407" heatid="19395" lane="0" entrytime="00:01:14.87" />
                <RESULT eventid="1457" status="DNS" swimtime="00:00:00.00" resultid="15408" heatid="19469" lane="1" entrytime="00:01:11.53" />
                <RESULT eventid="1630" status="DNS" swimtime="00:00:00.00" resultid="15409" heatid="19529" lane="7" entrytime="00:02:40.63" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-09-12" firstname="Wojciech" gender="M" lastname="Galczynski" nation="POL" athleteid="15380">
              <RESULTS>
                <RESULT eventid="1079" status="WDR" swimtime="00:00:00.00" resultid="15381" entrytime="00:00:26.20" />
                <RESULT eventid="1205" status="WDR" swimtime="00:00:00.00" resultid="15382" entrytime="00:00:32.60" />
                <RESULT eventid="14243" status="WDR" swimtime="00:00:00.00" resultid="15383" entrytime="00:01:09.50" />
                <RESULT eventid="1474" status="WDR" swimtime="00:00:00.00" resultid="15384" entrytime="00:01:14.65" />
                <RESULT eventid="1681" status="WDR" swimtime="00:00:00.00" resultid="15385" entrytime="00:00:32.73" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02602" nation="POL" region="KUJ" clubid="17025" name="Toruń Multisport Team">
          <CONTACT city="Toruń" email="szufar@o2.pl" name="Szufarski Andrzej" phone="600898866" state="KUJ-P" street="Matejki 60/7" zip="87-100" />
          <ATHLETES>
            <ATHLETE birthdate="1984-01-15" firstname="Artur" gender="M" lastname="Rybicki" nation="POL" athleteid="17078">
              <RESULTS>
                <RESULT eventid="1079" points="420" reactiontime="+90" swimtime="00:00:27.05" resultid="17079" heatid="19297" lane="3" entrytime="00:00:28.00" />
                <RESULT eventid="1273" points="406" reactiontime="+82" swimtime="00:01:00.67" resultid="17080" heatid="19383" lane="0" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="308" reactiontime="+82" swimtime="00:00:32.28" resultid="17081" heatid="19455" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1681" points="219" reactiontime="+90" swimtime="00:00:41.85" resultid="17082" heatid="19550" lane="3" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-03-03" firstname="Henryk" gender="M" lastname="Zientara" nation="POL" athleteid="17071">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="17072" heatid="19284" lane="5" entrytime="00:00:46.20" />
                <RESULT eventid="1205" points="63" reactiontime="+72" swimtime="00:00:55.76" resultid="17073" heatid="19344" lane="7" entrytime="00:00:51.02" />
                <RESULT comment="K4 - Cykl ruchowy inny niż jeden ruch ramion i jadno kopnięcie nogami (Time: 10:21)" eventid="1239" reactiontime="+95" status="DSQ" swimtime="00:04:42.93" resultid="17074" heatid="19360" lane="8" entrytime="00:04:19.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.06" />
                    <SPLIT distance="100" swimtime="00:02:11.83" />
                    <SPLIT distance="150" swimtime="00:03:29.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="86" reactiontime="+94" swimtime="00:02:05.79" resultid="17075" heatid="19434" lane="4" entrytime="00:01:59.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="48" reactiontime="+86" swimtime="00:02:13.87" resultid="17076" heatid="19471" lane="7" entrytime="00:02:11.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="17077" heatid="19548" lane="5" entrytime="00:00:51.02" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-10-25" firstname="Katarzyna" gender="F" lastname="Walenta" nation="POL" athleteid="17030">
              <RESULTS>
                <RESULT eventid="1062" points="496" reactiontime="+78" swimtime="00:00:29.34" resultid="17031" heatid="19275" lane="1" />
                <RESULT eventid="1096" points="462" reactiontime="+79" swimtime="00:02:37.55" resultid="17032" heatid="19309" lane="7" entrytime="00:02:39.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.52" />
                    <SPLIT distance="100" swimtime="00:01:14.06" />
                    <SPLIT distance="150" swimtime="00:01:59.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="424" reactiontime="+78" swimtime="00:02:59.04" resultid="17033" heatid="19358" lane="3" entrytime="00:02:55.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.72" />
                    <SPLIT distance="100" swimtime="00:01:25.87" />
                    <SPLIT distance="150" swimtime="00:02:12.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="479" reactiontime="+79" swimtime="00:01:12.38" resultid="17034" heatid="19395" lane="3" entrytime="00:01:13.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="440" reactiontime="+81" swimtime="00:01:21.97" resultid="17035" heatid="19432" lane="1" entrytime="00:01:22.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.24" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1555" points="442" reactiontime="+82" swimtime="00:05:40.51" resultid="17036" heatid="19505" lane="7" entrytime="00:05:45.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                    <SPLIT distance="100" swimtime="00:01:18.02" />
                    <SPLIT distance="150" swimtime="00:02:02.62" />
                    <SPLIT distance="200" swimtime="00:02:46.22" />
                    <SPLIT distance="250" swimtime="00:03:33.26" />
                    <SPLIT distance="300" swimtime="00:04:21.33" />
                    <SPLIT distance="350" swimtime="00:05:02.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="412" reactiontime="+82" swimtime="00:00:38.47" resultid="17037" heatid="19544" lane="1" entrytime="00:00:38.24" />
                <RESULT eventid="1721" points="422" reactiontime="+84" swimtime="00:05:12.65" resultid="17038" heatid="19697" lane="9" entrytime="00:06:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                    <SPLIT distance="100" swimtime="00:01:15.05" />
                    <SPLIT distance="150" swimtime="00:01:55.29" />
                    <SPLIT distance="200" swimtime="00:02:35.44" />
                    <SPLIT distance="250" swimtime="00:03:55.85" />
                    <SPLIT distance="300" swimtime="00:04:35.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-09-24" firstname="Anita" gender="F" lastname="Śliwa" nation="POL" athleteid="17097">
              <RESULTS>
                <RESULT eventid="1096" points="208" reactiontime="+116" swimtime="00:03:25.60" resultid="17098" heatid="19306" lane="1" entrytime="00:03:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.06" />
                    <SPLIT distance="100" swimtime="00:01:35.15" />
                    <SPLIT distance="150" swimtime="00:02:38.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="220" reactiontime="+114" swimtime="00:13:13.39" resultid="17099" heatid="19595" lane="6" entrytime="00:12:46.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.90" />
                    <SPLIT distance="100" swimtime="00:01:30.59" />
                    <SPLIT distance="150" swimtime="00:02:20.04" />
                    <SPLIT distance="200" swimtime="00:03:10.74" />
                    <SPLIT distance="250" swimtime="00:04:01.90" />
                    <SPLIT distance="300" swimtime="00:04:52.94" />
                    <SPLIT distance="350" swimtime="00:05:43.82" />
                    <SPLIT distance="400" swimtime="00:06:34.08" />
                    <SPLIT distance="450" swimtime="00:07:24.78" />
                    <SPLIT distance="500" swimtime="00:08:16.20" />
                    <SPLIT distance="550" swimtime="00:09:06.36" />
                    <SPLIT distance="600" swimtime="00:09:57.17" />
                    <SPLIT distance="650" swimtime="00:10:47.35" />
                    <SPLIT distance="700" swimtime="00:11:37.44" />
                    <SPLIT distance="750" swimtime="00:12:27.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="223" reactiontime="+97" swimtime="00:00:42.30" resultid="17100" heatid="19338" lane="8" entrytime="00:00:43.20" />
                <RESULT eventid="14225" points="207" reactiontime="+101" swimtime="00:01:35.65" resultid="17101" heatid="19391" lane="7" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="198" reactiontime="+92" swimtime="00:01:34.38" resultid="17102" heatid="19466" lane="3" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="230" reactiontime="+100" swimtime="00:03:00.61" resultid="17103" heatid="19481" lane="6" entrytime="00:03:14.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                    <SPLIT distance="100" swimtime="00:01:25.55" />
                    <SPLIT distance="150" swimtime="00:02:14.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="205" reactiontime="+100" swimtime="00:03:22.06" resultid="17104" heatid="19527" lane="3" entrytime="00:03:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.55" />
                    <SPLIT distance="100" swimtime="00:01:39.56" />
                    <SPLIT distance="150" swimtime="00:03:22.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="235" reactiontime="+103" swimtime="00:06:19.50" resultid="17105" heatid="19696" lane="3" entrytime="00:06:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.19" />
                    <SPLIT distance="100" swimtime="00:01:28.04" />
                    <SPLIT distance="150" swimtime="00:02:16.97" />
                    <SPLIT distance="200" swimtime="00:03:05.79" />
                    <SPLIT distance="250" swimtime="00:03:54.60" />
                    <SPLIT distance="300" swimtime="00:04:43.88" />
                    <SPLIT distance="350" swimtime="00:05:33.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-08-24" firstname="Jan" gender="M" lastname="Bantkowski" nation="POL" athleteid="17052">
              <RESULTS>
                <RESULT eventid="1113" points="54" reactiontime="+114" swimtime="00:04:49.98" resultid="17053" heatid="19312" lane="8" entrytime="00:05:02.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.47" />
                    <SPLIT distance="100" swimtime="00:02:26.27" />
                    <SPLIT distance="150" swimtime="00:03:52.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="28" reactiontime="+109" swimtime="00:01:12.77" resultid="17054" heatid="19343" lane="0" entrytime="00:01:05.38" />
                <RESULT eventid="1341" status="DNS" swimtime="00:00:00.00" resultid="17055" heatid="19413" lane="5" entrytime="00:05:07.78" />
                <RESULT eventid="1474" points="30" reactiontime="+88" swimtime="00:02:36.05" resultid="17056" heatid="19470" lane="5" entrytime="00:02:24.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="49" reactiontime="+127" swimtime="00:10:43.14" resultid="17057" heatid="19506" lane="4" entrytime="00:10:49.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.04" />
                    <SPLIT distance="100" swimtime="00:02:33.95" />
                    <SPLIT distance="150" swimtime="00:04:06.79" />
                    <SPLIT distance="200" swimtime="00:05:32.28" />
                    <SPLIT distance="250" swimtime="00:07:08.66" />
                    <SPLIT distance="300" swimtime="00:08:42.24" />
                    <SPLIT distance="350" swimtime="00:09:44.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="32" swimtime="00:02:31.32" resultid="17058" heatid="19517" lane="0" entrytime="00:02:20.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="28" reactiontime="+83" swimtime="00:05:46.27" resultid="17059" heatid="19531" lane="3" entrytime="00:05:04.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.83" />
                    <SPLIT distance="100" swimtime="00:02:56.58" />
                    <SPLIT distance="150" swimtime="00:04:25.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-10-13" firstname="Edward" gender="M" lastname="Korolko" nation="POL" athleteid="17060">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="17061" heatid="19285" lane="6" entrytime="00:00:42.00" />
                <RESULT eventid="1205" points="38" reactiontime="+70" swimtime="00:01:05.80" resultid="17062" heatid="19343" lane="9" entrytime="00:01:05.40" />
                <RESULT eventid="1273" points="76" reactiontime="+122" swimtime="00:01:45.64" resultid="17063" heatid="19375" lane="9" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="42" swimtime="00:02:19.91" resultid="17064" heatid="19471" lane="8" entrytime="00:02:15.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="17065" heatid="19486" lane="7" entrytime="00:04:40.50" />
                <RESULT eventid="1647" points="30" reactiontime="+88" swimtime="00:05:36.27" resultid="17066" heatid="19531" lane="4" entrytime="00:04:50.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.67" />
                    <SPLIT distance="100" swimtime="00:02:43.02" />
                    <SPLIT distance="150" swimtime="00:04:10.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-08-21" firstname="Tomasz" gender="M" lastname="Osóbka" nation="POL" athleteid="17067">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="17068" heatid="19284" lane="2" entrytime="00:01:02.45" />
                <RESULT eventid="1273" points="15" reactiontime="+137" swimtime="00:02:58.69" resultid="17069" heatid="19376" lane="3" entrytime="00:02:40.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="17070" heatid="19547" lane="8" entrytime="00:01:15.45" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-10-28" firstname="Andrzej" gender="M" lastname="Gołembiewski" nation="POL" athleteid="17083">
              <RESULTS>
                <RESULT eventid="14207" points="443" reactiontime="+86" swimtime="00:18:32.22" resultid="17084" heatid="19623" lane="5" entrytime="00:18:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                    <SPLIT distance="100" swimtime="00:01:05.42" />
                    <SPLIT distance="150" swimtime="00:01:40.53" />
                    <SPLIT distance="200" swimtime="00:02:16.44" />
                    <SPLIT distance="250" swimtime="00:02:52.78" />
                    <SPLIT distance="300" swimtime="00:03:29.65" />
                    <SPLIT distance="350" swimtime="00:04:07.08" />
                    <SPLIT distance="400" swimtime="00:04:44.48" />
                    <SPLIT distance="450" swimtime="00:05:22.01" />
                    <SPLIT distance="500" swimtime="00:05:59.49" />
                    <SPLIT distance="550" swimtime="00:06:37.26" />
                    <SPLIT distance="600" swimtime="00:07:15.12" />
                    <SPLIT distance="650" swimtime="00:07:53.02" />
                    <SPLIT distance="700" swimtime="00:08:30.95" />
                    <SPLIT distance="750" swimtime="00:09:09.11" />
                    <SPLIT distance="800" swimtime="00:09:46.69" />
                    <SPLIT distance="850" swimtime="00:10:24.15" />
                    <SPLIT distance="900" swimtime="00:11:02.25" />
                    <SPLIT distance="950" swimtime="00:11:39.90" />
                    <SPLIT distance="1000" swimtime="00:12:17.70" />
                    <SPLIT distance="1050" swimtime="00:12:55.51" />
                    <SPLIT distance="1100" swimtime="00:13:33.62" />
                    <SPLIT distance="1150" swimtime="00:14:11.45" />
                    <SPLIT distance="1200" swimtime="00:14:49.39" />
                    <SPLIT distance="1250" swimtime="00:15:26.61" />
                    <SPLIT distance="1300" swimtime="00:16:03.73" />
                    <SPLIT distance="1350" swimtime="00:16:41.68" />
                    <SPLIT distance="1400" swimtime="00:17:19.73" />
                    <SPLIT distance="1450" swimtime="00:17:57.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="471" reactiontime="+89" swimtime="00:02:34.70" resultid="17085" heatid="19364" lane="3" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                    <SPLIT distance="100" swimtime="00:01:14.70" />
                    <SPLIT distance="150" swimtime="00:01:54.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="524" reactiontime="+80" swimtime="00:01:08.95" resultid="17086" heatid="19442" lane="5" entrytime="00:01:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="478" reactiontime="+79" swimtime="00:02:07.07" resultid="17087" heatid="19496" lane="0" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.38" />
                    <SPLIT distance="100" swimtime="00:01:01.16" />
                    <SPLIT distance="150" swimtime="00:01:34.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="493" reactiontime="+75" swimtime="00:00:31.96" resultid="17088" heatid="19559" lane="7" entrytime="00:00:31.70" />
                <RESULT eventid="1744" points="479" reactiontime="+78" swimtime="00:04:31.22" resultid="17089" heatid="19708" lane="8" entrytime="00:04:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.10" />
                    <SPLIT distance="100" swimtime="00:01:03.22" />
                    <SPLIT distance="150" swimtime="00:01:36.95" />
                    <SPLIT distance="200" swimtime="00:02:11.29" />
                    <SPLIT distance="250" swimtime="00:02:46.15" />
                    <SPLIT distance="300" swimtime="00:03:21.50" />
                    <SPLIT distance="350" swimtime="00:03:57.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-03-07" firstname="Grzegorz" gender="M" lastname="Arentewicz" nation="POL" athleteid="17039">
              <RESULTS>
                <RESULT eventid="1079" points="298" reactiontime="+89" swimtime="00:00:30.30" resultid="17040" heatid="19291" lane="5" entrytime="00:00:31.20" />
                <RESULT eventid="1273" points="296" reactiontime="+92" swimtime="00:01:07.36" resultid="17041" heatid="19380" lane="2" entrytime="00:01:08.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" status="DNS" swimtime="00:00:00.00" resultid="17042" heatid="19416" lane="0" entrytime="00:03:08.15" />
                <RESULT eventid="1440" points="304" reactiontime="+83" swimtime="00:00:32.40" resultid="17043" heatid="19456" lane="8" entrytime="00:00:32.70" />
                <RESULT eventid="1508" points="248" reactiontime="+89" swimtime="00:02:38.10" resultid="17044" heatid="19490" lane="7" entrytime="00:02:42.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                    <SPLIT distance="100" swimtime="00:01:16.56" />
                    <SPLIT distance="150" swimtime="00:01:57.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="241" reactiontime="+93" swimtime="00:01:17.17" resultid="17045" heatid="19520" lane="7" entrytime="00:01:18.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="250" reactiontime="+98" swimtime="00:05:36.89" resultid="17046" heatid="19703" lane="5" entrytime="00:05:44.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.10" />
                    <SPLIT distance="100" swimtime="00:01:20.17" />
                    <SPLIT distance="150" swimtime="00:02:03.37" />
                    <SPLIT distance="200" swimtime="00:02:47.04" />
                    <SPLIT distance="250" swimtime="00:03:30.69" />
                    <SPLIT distance="300" swimtime="00:04:13.84" />
                    <SPLIT distance="350" swimtime="00:04:56.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-10-11" firstname="Kamil" gender="M" lastname="Kordowski" nation="POL" athleteid="17026">
              <RESULTS>
                <RESULT eventid="1079" points="373" reactiontime="+93" swimtime="00:00:28.14" resultid="17027" heatid="19298" lane="1" entrytime="00:00:27.53" />
                <RESULT eventid="1273" points="348" reactiontime="+89" swimtime="00:01:03.86" resultid="17028" heatid="19381" lane="5" entrytime="00:01:05.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="336" reactiontime="+80" swimtime="00:00:31.33" resultid="17029" heatid="19456" lane="6" entrytime="00:00:32.29" />
                <RESULT eventid="1744" points="219" reactiontime="+95" swimtime="00:05:51.86" resultid="18343" heatid="19701" lane="3" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.10" />
                    <SPLIT distance="100" swimtime="00:01:17.60" />
                    <SPLIT distance="150" swimtime="00:02:01.03" />
                    <SPLIT distance="200" swimtime="00:02:45.23" />
                    <SPLIT distance="250" swimtime="00:03:30.98" />
                    <SPLIT distance="300" swimtime="00:04:18.13" />
                    <SPLIT distance="350" swimtime="00:05:04.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="266" reactiontime="+91" swimtime="00:02:34.42" resultid="18472" heatid="19485" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                    <SPLIT distance="100" swimtime="00:01:12.09" />
                    <SPLIT distance="150" swimtime="00:01:55.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="238" reactiontime="+91" swimtime="00:01:17.52" resultid="18473" heatid="19516" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-02-04" firstname="Andrzej" gender="M" lastname="Marchewka" nation="POL" athleteid="17047">
              <RESULTS>
                <RESULT eventid="1205" points="341" reactiontime="+77" swimtime="00:00:31.80" resultid="17048" heatid="19349" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="14243" points="348" reactiontime="+88" swimtime="00:01:11.46" resultid="17049" heatid="19404" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="327" reactiontime="+64" swimtime="00:01:10.97" resultid="17050" heatid="19476" lane="8" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="263" reactiontime="+75" swimtime="00:02:44.74" resultid="17051" heatid="19535" lane="4" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.56" />
                    <SPLIT distance="100" swimtime="00:01:18.27" />
                    <SPLIT distance="150" swimtime="00:02:01.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-04-23" firstname="Krzysztof" gender="M" lastname="Lietz" nation="POL" athleteid="17106">
              <RESULTS>
                <RESULT eventid="1079" points="237" reactiontime="+101" swimtime="00:00:32.73" resultid="17107" heatid="19290" lane="1" entrytime="00:00:32.80" />
                <RESULT eventid="14189" points="183" reactiontime="+87" swimtime="00:13:00.73" resultid="17108" heatid="19616" lane="9" entrytime="00:13:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                    <SPLIT distance="100" swimtime="00:01:27.94" />
                    <SPLIT distance="150" swimtime="00:02:15.49" />
                    <SPLIT distance="200" swimtime="00:03:55.62" />
                    <SPLIT distance="300" swimtime="00:04:46.05" />
                    <SPLIT distance="350" swimtime="00:05:35.84" />
                    <SPLIT distance="450" swimtime="00:06:26.56" />
                    <SPLIT distance="500" swimtime="00:07:16.98" />
                    <SPLIT distance="550" swimtime="00:08:06.76" />
                    <SPLIT distance="600" swimtime="00:08:56.61" />
                    <SPLIT distance="650" swimtime="00:09:47.11" />
                    <SPLIT distance="700" swimtime="00:10:37.53" />
                    <SPLIT distance="750" swimtime="00:11:26.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="216" reactiontime="+85" swimtime="00:01:14.83" resultid="17109" heatid="19378" lane="5" entrytime="00:01:13.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="181" reactiontime="+80" swimtime="00:01:28.83" resultid="17110" heatid="19401" lane="9" entrytime="00:01:25.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="225" reactiontime="+89" swimtime="00:00:35.79" resultid="17111" heatid="19453" lane="3" entrytime="00:00:36.80" />
                <RESULT eventid="1508" points="186" reactiontime="+90" swimtime="00:02:53.80" resultid="17112" heatid="19489" lane="7" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.30" />
                    <SPLIT distance="100" swimtime="00:01:25.13" />
                    <SPLIT distance="150" swimtime="00:02:11.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="131" reactiontime="+86" swimtime="00:01:34.43" resultid="17113" heatid="19519" lane="9" entrytime="00:01:33.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="181" reactiontime="+86" swimtime="00:06:14.69" resultid="17114" heatid="19702" lane="1" entrytime="00:06:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.33" />
                    <SPLIT distance="100" swimtime="00:01:29.08" />
                    <SPLIT distance="150" swimtime="00:02:16.62" />
                    <SPLIT distance="200" swimtime="00:03:06.85" />
                    <SPLIT distance="250" swimtime="00:03:56.51" />
                    <SPLIT distance="300" swimtime="00:04:46.02" />
                    <SPLIT distance="350" swimtime="00:05:32.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-06-29" firstname="Lucyna" gender="F" lastname="Serożyńska" nation="POL" athleteid="17090">
              <RESULTS>
                <RESULT eventid="1062" points="109" reactiontime="+110" swimtime="00:00:48.60" resultid="17091" heatid="19276" lane="8" entrytime="00:00:53.56" />
                <RESULT eventid="1187" points="64" reactiontime="+93" swimtime="00:01:04.07" resultid="17092" heatid="19336" lane="3" entrytime="00:01:01.18" />
                <RESULT eventid="1256" points="72" reactiontime="+121" swimtime="00:02:02.11" resultid="17093" heatid="19367" lane="5" entrytime="00:01:55.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="114" reactiontime="+108" swimtime="00:02:08.25" resultid="17094" heatid="19428" lane="9" entrytime="00:02:07.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="67" reactiontime="+95" swimtime="00:02:15.48" resultid="17095" heatid="19465" lane="5" entrytime="00:02:19.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="67" reactiontime="+103" swimtime="00:04:52.91" resultid="17096" heatid="19526" lane="6" entrytime="00:05:02.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.43" />
                    <SPLIT distance="100" swimtime="00:02:22.25" />
                    <SPLIT distance="150" swimtime="00:03:39.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="93" swimtime="00:03:19.77" resultid="17115" heatid="19421" lane="7" entrytime="00:03:14.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.87" />
                    <SPLIT distance="100" swimtime="00:01:55.04" />
                    <SPLIT distance="150" swimtime="00:02:33.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17060" number="1" />
                    <RELAYPOSITION athleteid="17071" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="17106" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="17052" number="4" reactiontime="+108" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="108" reactiontime="+98" swimtime="00:02:53.04" resultid="17116" heatid="19499" lane="2" entrytime="00:02:53.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.98" />
                    <SPLIT distance="100" swimtime="00:01:08.29" />
                    <SPLIT distance="150" swimtime="00:02:20.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17060" number="1" reactiontime="+98" />
                    <RELAYPOSITION athleteid="17052" number="2" reactiontime="+90" />
                    <RELAYPOSITION athleteid="17071" number="3" />
                    <RELAYPOSITION athleteid="17106" number="4" reactiontime="+65" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1548" points="423" reactiontime="+91" swimtime="00:01:49.97" resultid="17119" heatid="19501" lane="2" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.44" />
                    <SPLIT distance="100" swimtime="00:00:57.33" />
                    <SPLIT distance="150" swimtime="00:01:24.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17047" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="17039" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="17078" number="3" reactiontime="+16" />
                    <RELAYPOSITION athleteid="17083" number="4" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1381" points="388" reactiontime="+86" swimtime="00:02:04.02" resultid="17120" heatid="19424" lane="0" entrytime="00:02:01.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.42" />
                    <SPLIT distance="100" swimtime="00:01:04.89" />
                    <SPLIT distance="150" swimtime="00:01:36.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17047" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="17083" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="17039" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="17078" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1130" points="410" reactiontime="+74" swimtime="00:01:59.20" resultid="17117" heatid="19322" lane="9" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.89" />
                    <SPLIT distance="100" swimtime="00:01:06.25" />
                    <SPLIT distance="150" swimtime="00:01:33.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17030" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="17097" number="2" reactiontime="+90" />
                    <RELAYPOSITION athleteid="17078" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="17083" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="384" swimtime="00:02:13.58" resultid="17118" heatid="19564" lane="8" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.02" />
                    <SPLIT distance="100" swimtime="00:01:14.14" />
                    <SPLIT distance="150" swimtime="00:01:47.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17097" number="1" />
                    <RELAYPOSITION athleteid="17083" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="17030" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="17047" number="4" reactiontime="+9" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="KUJ" clubid="18403" name="Toruński Klub Triathlonowy">
          <CONTACT email="agusianamberone@poczta.onet.pl" name="KOSTYRA AGNIESZKA" phone="722053277" state="KUJ" />
          <ATHLETES>
            <ATHLETE birthdate="1990-02-16" firstname="Agnieszka" gender="F" lastname="Kostyra" nation="POL" athleteid="18409">
              <RESULTS>
                <RESULT eventid="1096" points="303" reactiontime="+65" swimtime="00:03:01.30" resultid="18410" heatid="19307" lane="9" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                    <SPLIT distance="100" swimtime="00:01:23.80" />
                    <SPLIT distance="150" swimtime="00:02:17.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" reactiontime="+86" status="OTL" swimtime="00:11:50.74" resultid="18411" heatid="19595" lane="3" entrytime="00:12:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.45" />
                    <SPLIT distance="100" swimtime="00:01:19.81" />
                    <SPLIT distance="150" swimtime="00:02:03.69" />
                    <SPLIT distance="200" swimtime="00:02:48.13" />
                    <SPLIT distance="250" swimtime="00:03:32.91" />
                    <SPLIT distance="300" swimtime="00:04:18.21" />
                    <SPLIT distance="350" swimtime="00:05:03.86" />
                    <SPLIT distance="400" swimtime="00:05:48.73" />
                    <SPLIT distance="450" swimtime="00:06:33.93" />
                    <SPLIT distance="500" swimtime="00:07:19.55" />
                    <SPLIT distance="550" swimtime="00:08:05.37" />
                    <SPLIT distance="600" swimtime="00:08:50.96" />
                    <SPLIT distance="650" swimtime="00:09:36.30" />
                    <SPLIT distance="700" swimtime="00:10:21.64" />
                    <SPLIT distance="750" swimtime="00:11:07.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="OLPOZ" nation="POL" region="WIE" clubid="17720" name="TS Olimpia Poznań">
          <CONTACT name="Pietraszewski" phone="501 648 415" />
          <ATHLETES>
            <ATHLETE birthdate="1955-01-01" firstname="Zbigniew" gender="M" lastname="Pietraszewski" nation="POL" athleteid="17745">
              <RESULTS>
                <RESULT eventid="1113" points="200" reactiontime="+91" swimtime="00:03:07.26" resultid="17746" heatid="19312" lane="9" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.06" />
                    <SPLIT distance="100" swimtime="00:01:32.52" />
                    <SPLIT distance="150" swimtime="00:02:24.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14189" points="200" reactiontime="+103" swimtime="00:12:38.16" resultid="17747" heatid="19616" lane="0" entrytime="00:12:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.21" />
                    <SPLIT distance="100" swimtime="00:01:28.35" />
                    <SPLIT distance="150" swimtime="00:02:15.69" />
                    <SPLIT distance="200" swimtime="00:03:03.31" />
                    <SPLIT distance="250" swimtime="00:03:51.13" />
                    <SPLIT distance="300" swimtime="00:04:39.08" />
                    <SPLIT distance="350" swimtime="00:05:27.64" />
                    <SPLIT distance="400" swimtime="00:06:16.47" />
                    <SPLIT distance="450" swimtime="00:07:04.61" />
                    <SPLIT distance="500" swimtime="00:07:52.64" />
                    <SPLIT distance="550" swimtime="00:08:40.70" />
                    <SPLIT distance="600" swimtime="00:09:29.07" />
                    <SPLIT distance="650" swimtime="00:10:16.76" />
                    <SPLIT distance="700" swimtime="00:11:04.55" />
                    <SPLIT distance="750" swimtime="00:11:52.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="153" reactiontime="+74" swimtime="00:00:41.54" resultid="17748" heatid="19346" lane="9" entrytime="00:00:42.00" />
                <RESULT eventid="14243" points="213" reactiontime="+94" swimtime="00:01:24.22" resultid="17749" heatid="19401" lane="7" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="176" reactiontime="+87" swimtime="00:01:27.19" resultid="17750" heatid="19473" lane="4" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="193" reactiontime="+97" swimtime="00:06:47.33" resultid="17751" heatid="19509" lane="9" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.38" />
                    <SPLIT distance="100" swimtime="00:01:43.59" />
                    <SPLIT distance="150" swimtime="00:02:32.87" />
                    <SPLIT distance="200" swimtime="00:03:22.32" />
                    <SPLIT distance="250" swimtime="00:04:16.93" />
                    <SPLIT distance="300" swimtime="00:05:13.39" />
                    <SPLIT distance="350" swimtime="00:06:01.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="169" reactiontime="+92" swimtime="00:03:10.85" resultid="17752" heatid="19534" lane="1" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.33" />
                    <SPLIT distance="100" swimtime="00:01:32.81" />
                    <SPLIT distance="150" swimtime="00:02:21.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="17753" heatid="19702" lane="2" entrytime="00:06:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Jerzy" gender="M" lastname="Boryski" nation="POL" athleteid="17731">
              <RESULTS>
                <RESULT eventid="1079" points="146" reactiontime="+102" swimtime="00:00:38.45" resultid="17732" heatid="19287" lane="1" entrytime="00:00:37.50" />
                <RESULT eventid="14189" points="126" reactiontime="+108" swimtime="00:14:43.49" resultid="17733" heatid="19615" lane="2" entrytime="00:14:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.50" />
                    <SPLIT distance="100" swimtime="00:01:41.53" />
                    <SPLIT distance="150" swimtime="00:02:36.30" />
                    <SPLIT distance="200" swimtime="00:03:31.77" />
                    <SPLIT distance="250" swimtime="00:04:27.28" />
                    <SPLIT distance="300" swimtime="00:05:23.02" />
                    <SPLIT distance="350" swimtime="00:06:18.46" />
                    <SPLIT distance="400" swimtime="00:07:14.41" />
                    <SPLIT distance="450" swimtime="00:08:10.07" />
                    <SPLIT distance="500" swimtime="00:09:06.51" />
                    <SPLIT distance="550" swimtime="00:10:03.61" />
                    <SPLIT distance="600" swimtime="00:11:00.23" />
                    <SPLIT distance="650" swimtime="00:11:57.08" />
                    <SPLIT distance="700" swimtime="00:12:54.20" />
                    <SPLIT distance="750" swimtime="00:13:50.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="141" reactiontime="+80" swimtime="00:00:42.61" resultid="17734" heatid="19345" lane="6" entrytime="00:00:43.00" />
                <RESULT eventid="1474" points="119" reactiontime="+80" swimtime="00:01:39.23" resultid="17735" heatid="19472" lane="5" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="99" reactiontime="+109" swimtime="00:03:47.77" resultid="17736" heatid="19533" lane="0" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.60" />
                    <SPLIT distance="100" swimtime="00:01:51.13" />
                    <SPLIT distance="150" swimtime="00:02:52.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="121" reactiontime="+107" swimtime="00:07:08.87" resultid="17737" heatid="19700" lane="5" entrytime="00:07:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.68" />
                    <SPLIT distance="100" swimtime="00:01:41.65" />
                    <SPLIT distance="150" swimtime="00:02:35.67" />
                    <SPLIT distance="200" swimtime="00:03:30.87" />
                    <SPLIT distance="250" swimtime="00:04:26.31" />
                    <SPLIT distance="300" swimtime="00:05:21.28" />
                    <SPLIT distance="350" swimtime="00:06:16.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Maria" gender="F" lastname="Łutowicz" nation="POL" athleteid="17722">
              <RESULTS>
                <RESULT eventid="1062" points="190" reactiontime="+98" swimtime="00:00:40.36" resultid="17723" heatid="19277" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1096" points="141" reactiontime="+99" swimtime="00:03:53.81" resultid="17724" heatid="19305" lane="5" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.53" />
                    <SPLIT distance="100" swimtime="00:01:55.48" />
                    <SPLIT distance="150" swimtime="00:03:03.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="149" reactiontime="+44" swimtime="00:00:48.38" resultid="17725" heatid="19337" lane="1" entrytime="00:00:53.00" />
                <RESULT eventid="1256" points="161" reactiontime="+99" swimtime="00:01:33.46" resultid="17726" heatid="19368" lane="6" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="123" reactiontime="+100" swimtime="00:00:49.01" resultid="17727" heatid="19445" lane="1" entrytime="00:00:53.00" />
                <RESULT eventid="1491" points="160" reactiontime="+99" swimtime="00:03:23.73" resultid="17728" heatid="19480" lane="4" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.20" />
                    <SPLIT distance="100" swimtime="00:01:40.58" />
                    <SPLIT distance="150" swimtime="00:02:34.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="159" swimtime="00:00:52.86" resultid="17729" heatid="19540" lane="0" entrytime="00:00:54.00" />
                <RESULT eventid="1721" points="155" reactiontime="+90" swimtime="00:07:16.10" resultid="17730" heatid="19696" lane="9" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.67" />
                    <SPLIT distance="100" swimtime="00:01:44.58" />
                    <SPLIT distance="150" swimtime="00:02:41.76" />
                    <SPLIT distance="200" swimtime="00:03:38.06" />
                    <SPLIT distance="250" swimtime="00:04:34.30" />
                    <SPLIT distance="300" swimtime="00:05:30.21" />
                    <SPLIT distance="350" swimtime="00:06:24.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-01-01" firstname="Jacek" gender="M" lastname="Lesiński" nation="POL" athleteid="17738">
              <RESULTS>
                <RESULT eventid="1113" points="121" reactiontime="+103" swimtime="00:03:41.06" resultid="17739" heatid="19311" lane="0" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.25" />
                    <SPLIT distance="100" swimtime="00:01:48.53" />
                    <SPLIT distance="150" swimtime="00:02:51.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="17740" heatid="19345" lane="8" entrytime="00:00:45.00" />
                <RESULT eventid="14243" status="DNS" swimtime="00:00:00.00" resultid="17741" heatid="19399" lane="8" entrytime="00:01:45.00" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="17742" heatid="19472" lane="7" entrytime="00:01:45.00" />
                <RESULT eventid="1647" points="102" reactiontime="+84" swimtime="00:03:45.61" resultid="17743" heatid="19532" lane="4" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.17" />
                    <SPLIT distance="100" swimtime="00:01:49.33" />
                    <SPLIT distance="150" swimtime="00:02:48.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="143" reactiontime="+111" swimtime="00:00:48.21" resultid="17744" heatid="19549" lane="9" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01414" nation="POL" region="WA" clubid="14761" name="UKS Delfin Legionowo">
          <CONTACT city="LEGIONOWO" email="delfin-trener@wp.pl" internet="www.delfinlegionowo.pl" name="RAFAŁ PERL" phone="601 436 700" state="MAZ" street="KRÓLOWEJ JADWIGI 11" zip="05-120" />
          <ATHLETES>
            <ATHLETE birthdate="1997-06-23" firstname="Krzysztof" gender="M" lastname="Żbikowski" nation="POL" athleteid="14770">
              <RESULTS>
                <RESULT eventid="1079" points="513" reactiontime="+71" swimtime="00:00:25.30" resultid="14771" heatid="19301" lane="9" entrytime="00:00:26.00" />
                <RESULT comment="G1 - Głowa pływaka nie złamała powierzchni wody przed lub na lini 15m (Time: 9:31)" eventid="1205" reactiontime="+79" status="DSQ" swimtime="00:00:30.59" resultid="14772" heatid="19352" lane="0" entrytime="00:00:30.00" />
                <RESULT eventid="1406" points="585" reactiontime="+81" swimtime="00:01:06.48" resultid="14773" heatid="19443" lane="0" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="514" reactiontime="+75" swimtime="00:00:27.20" resultid="14774" heatid="19461" lane="5" entrytime="00:00:28.00" />
                <RESULT eventid="1681" points="616" reactiontime="+70" swimtime="00:00:29.67" resultid="14775" heatid="19560" lane="8" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-06-07" firstname="Michał" gender="M" lastname="Perl" nation="POL" athleteid="14762">
              <RESULTS>
                <RESULT eventid="1079" points="618" reactiontime="+75" swimtime="00:00:23.78" resultid="14763" heatid="19304" lane="3" entrytime="00:00:23.57" />
                <RESULT eventid="1273" points="574" reactiontime="+69" swimtime="00:00:54.05" resultid="14764" heatid="19388" lane="8" entrytime="00:00:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="515" reactiontime="+70" swimtime="00:01:02.74" resultid="14765" heatid="19410" lane="9" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="579" reactiontime="+72" swimtime="00:01:06.72" resultid="14766" heatid="19443" lane="5" entrytime="00:01:03.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="570" reactiontime="+72" swimtime="00:00:26.29" resultid="14767" heatid="19463" lane="4" entrytime="00:00:26.39" />
                <RESULT eventid="1681" points="632" reactiontime="+71" swimtime="00:00:29.41" resultid="14768" heatid="19560" lane="4" entrytime="00:00:28.26" />
                <RESULT eventid="1744" points="365" reactiontime="+78" swimtime="00:04:56.96" resultid="14769" heatid="19707" lane="5" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                    <SPLIT distance="100" swimtime="00:01:08.73" />
                    <SPLIT distance="150" swimtime="00:01:46.40" />
                    <SPLIT distance="200" swimtime="00:02:24.46" />
                    <SPLIT distance="250" swimtime="00:03:03.08" />
                    <SPLIT distance="300" swimtime="00:03:41.50" />
                    <SPLIT distance="350" swimtime="00:04:20.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-07-05" firstname="Karolina" gender="F" lastname="Modzelan" nation="POL" athleteid="14776">
              <RESULTS>
                <RESULT eventid="1062" points="428" reactiontime="+84" swimtime="00:00:30.83" resultid="14777" heatid="19282" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="14225" points="354" reactiontime="+92" swimtime="00:01:20.10" resultid="14778" heatid="19394" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="349" reactiontime="+72" swimtime="00:01:28.55" resultid="14779" heatid="19431" lane="0" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="360" reactiontime="+78" swimtime="00:00:40.25" resultid="14780" heatid="19543" lane="5" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00408" nation="POL" region="RZ" clubid="15998" name="UKS Delfin Masrers Tarnobrzeg">
          <CONTACT city="TARNOBRZEG" email="piotr.michalik@i-bs.pl" name="MICHALIK ANGELIKA" state="PODKA" street="SKALNA GÓRA 8/21" street2="TARNOBRZEG" zip="39-400" />
          <ATHLETES>
            <ATHLETE birthdate="1971-01-07" firstname="Albert" gender="M" lastname="Szwajkowski" nation="POL" athleteid="16082">
              <RESULTS>
                <RESULT eventid="1079" points="318" reactiontime="+97" swimtime="00:00:29.67" resultid="16083" heatid="19292" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="14207" reactiontime="+129" status="OTL" swimtime="00:00:00.00" resultid="16084" heatid="19621" lane="2" entrytime="00:24:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.17" />
                    <SPLIT distance="1450" swimtime="00:25:03.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" status="DNS" swimtime="00:00:00.00" resultid="16085" heatid="19403" lane="2" entrytime="00:01:16.00" />
                <RESULT eventid="1440" points="256" reactiontime="+93" swimtime="00:00:34.29" resultid="16086" heatid="19454" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="16097" heatid="19380" lane="0" entrytime="00:01:09.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-12" firstname="Maciej" gender="M" lastname="Płaneta" nation="POL" athleteid="16048">
              <RESULTS>
                <RESULT eventid="1079" points="325" reactiontime="+73" swimtime="00:00:29.44" resultid="16049" heatid="19293" lane="6" entrytime="00:00:29.80" />
                <RESULT eventid="14207" points="276" reactiontime="+80" swimtime="00:21:41.50" resultid="16050" heatid="19622" lane="7" entrytime="00:21:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                    <SPLIT distance="100" swimtime="00:01:17.75" />
                    <SPLIT distance="150" swimtime="00:01:59.53" />
                    <SPLIT distance="200" swimtime="00:02:40.91" />
                    <SPLIT distance="250" swimtime="00:03:22.56" />
                    <SPLIT distance="300" swimtime="00:04:04.92" />
                    <SPLIT distance="350" swimtime="00:04:47.43" />
                    <SPLIT distance="400" swimtime="00:05:29.93" />
                    <SPLIT distance="450" swimtime="00:06:13.04" />
                    <SPLIT distance="500" swimtime="00:06:56.19" />
                    <SPLIT distance="550" swimtime="00:07:38.59" />
                    <SPLIT distance="600" swimtime="00:08:21.74" />
                    <SPLIT distance="650" swimtime="00:09:05.71" />
                    <SPLIT distance="700" swimtime="00:09:49.37" />
                    <SPLIT distance="750" swimtime="00:10:32.84" />
                    <SPLIT distance="800" swimtime="00:11:16.67" />
                    <SPLIT distance="850" swimtime="00:12:01.04" />
                    <SPLIT distance="900" swimtime="00:12:45.31" />
                    <SPLIT distance="950" swimtime="00:13:29.90" />
                    <SPLIT distance="1000" swimtime="00:14:14.52" />
                    <SPLIT distance="1050" swimtime="00:14:59.29" />
                    <SPLIT distance="1100" swimtime="00:15:43.49" />
                    <SPLIT distance="1150" swimtime="00:16:28.68" />
                    <SPLIT distance="1200" swimtime="00:17:14.06" />
                    <SPLIT distance="1250" swimtime="00:17:58.97" />
                    <SPLIT distance="1300" swimtime="00:18:44.42" />
                    <SPLIT distance="1350" swimtime="00:19:29.86" />
                    <SPLIT distance="1400" swimtime="00:20:15.51" />
                    <SPLIT distance="1450" swimtime="00:21:00.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="320" swimtime="00:01:05.65" resultid="16051" heatid="19382" lane="0" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="228" reactiontime="+78" swimtime="00:02:57.47" resultid="16052" heatid="19416" lane="8" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.67" />
                    <SPLIT distance="100" swimtime="00:01:22.46" />
                    <SPLIT distance="150" swimtime="00:02:11.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="309" reactiontime="+79" swimtime="00:02:26.97" resultid="16053" heatid="19492" lane="1" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.30" />
                    <SPLIT distance="100" swimtime="00:01:11.31" />
                    <SPLIT distance="150" swimtime="00:01:49.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="251" reactiontime="+84" swimtime="00:06:12.98" resultid="16054" heatid="19509" lane="7" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.91" />
                    <SPLIT distance="100" swimtime="00:01:22.75" />
                    <SPLIT distance="150" swimtime="00:02:12.76" />
                    <SPLIT distance="200" swimtime="00:03:02.34" />
                    <SPLIT distance="250" swimtime="00:03:56.11" />
                    <SPLIT distance="300" swimtime="00:04:50.42" />
                    <SPLIT distance="350" swimtime="00:05:33.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="217" reactiontime="+76" swimtime="00:02:55.67" resultid="16055" heatid="19534" lane="7" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.44" />
                    <SPLIT distance="100" swimtime="00:01:25.90" />
                    <SPLIT distance="150" swimtime="00:02:12.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="290" reactiontime="+81" swimtime="00:05:20.31" resultid="16056" heatid="19705" lane="1" entrytime="00:05:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                    <SPLIT distance="100" swimtime="00:01:13.88" />
                    <SPLIT distance="150" swimtime="00:01:54.67" />
                    <SPLIT distance="200" swimtime="00:02:36.43" />
                    <SPLIT distance="250" swimtime="00:03:18.07" />
                    <SPLIT distance="300" swimtime="00:04:00.32" />
                    <SPLIT distance="350" swimtime="00:04:41.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-07-13" firstname="Piotr" gender="M" lastname="Hewelke" nation="POL" athleteid="16078">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="16079" heatid="19290" lane="9" entrytime="00:00:33.00" />
                <RESULT eventid="1205" points="251" reactiontime="+71" swimtime="00:00:35.20" resultid="16080" heatid="19347" lane="5" entrytime="00:00:37.00" />
                <RESULT eventid="1681" points="255" reactiontime="+81" swimtime="00:00:39.78" resultid="16081" heatid="19552" lane="5" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-04-24" firstname="Renata" gender="F" lastname="Osmala" nation="POL" athleteid="16006">
              <RESULTS>
                <RESULT eventid="1147" points="353" reactiontime="+91" swimtime="00:11:17.74" resultid="16007" heatid="19596" lane="0" entrytime="00:11:20.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                    <SPLIT distance="100" swimtime="00:01:17.67" />
                    <SPLIT distance="150" swimtime="00:01:59.75" />
                    <SPLIT distance="200" swimtime="00:02:42.07" />
                    <SPLIT distance="250" swimtime="00:03:24.87" />
                    <SPLIT distance="300" swimtime="00:04:07.72" />
                    <SPLIT distance="350" swimtime="00:04:50.66" />
                    <SPLIT distance="400" swimtime="00:05:33.64" />
                    <SPLIT distance="450" swimtime="00:06:16.63" />
                    <SPLIT distance="500" swimtime="00:06:59.75" />
                    <SPLIT distance="550" swimtime="00:07:42.73" />
                    <SPLIT distance="600" swimtime="00:08:26.03" />
                    <SPLIT distance="650" swimtime="00:09:09.68" />
                    <SPLIT distance="700" swimtime="00:09:53.30" />
                    <SPLIT distance="750" swimtime="00:10:36.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="290" reactiontime="+75" swimtime="00:00:38.77" resultid="16008" heatid="19339" lane="2" entrytime="00:00:38.95" />
                <RESULT eventid="1457" points="306" reactiontime="+73" swimtime="00:01:21.58" resultid="16009" heatid="19468" lane="9" entrytime="00:01:24.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="344" reactiontime="+89" swimtime="00:02:38.00" resultid="16010" heatid="19483" lane="6" entrytime="00:02:42.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                    <SPLIT distance="100" swimtime="00:01:16.55" />
                    <SPLIT distance="150" swimtime="00:01:57.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="330" reactiontime="+77" swimtime="00:02:52.46" resultid="16011" heatid="19529" lane="9" entrytime="00:02:56.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.72" />
                    <SPLIT distance="100" swimtime="00:01:23.97" />
                    <SPLIT distance="150" swimtime="00:02:08.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="353" reactiontime="+85" swimtime="00:05:31.83" resultid="16012" heatid="19698" lane="9" entrytime="00:05:40.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.62" />
                    <SPLIT distance="100" swimtime="00:01:19.18" />
                    <SPLIT distance="150" swimtime="00:02:01.38" />
                    <SPLIT distance="200" swimtime="00:02:44.00" />
                    <SPLIT distance="250" swimtime="00:03:26.28" />
                    <SPLIT distance="300" swimtime="00:04:08.96" />
                    <SPLIT distance="350" swimtime="00:04:51.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-03-30" firstname="Angelika" gender="F" lastname="Rozmus" nation="POL" athleteid="16057">
              <RESULTS>
                <RESULT eventid="1062" points="336" reactiontime="+91" swimtime="00:00:33.40" resultid="16058" heatid="19281" lane="1" entrytime="00:00:32.50" />
                <RESULT eventid="1096" points="316" reactiontime="+86" swimtime="00:02:58.79" resultid="16059" heatid="19308" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.16" />
                    <SPLIT distance="100" swimtime="00:01:25.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="292" reactiontime="+80" swimtime="00:03:22.71" resultid="16060" heatid="19358" lane="9" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.67" />
                    <SPLIT distance="100" swimtime="00:01:36.60" />
                    <SPLIT distance="150" swimtime="00:02:30.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" status="DNS" swimtime="00:00:00.00" resultid="16061" heatid="19394" lane="0" entrytime="00:01:21.50" />
                <RESULT eventid="1388" points="289" reactiontime="+88" swimtime="00:01:34.25" resultid="16062" heatid="19431" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="286" reactiontime="+94" swimtime="00:06:33.41" resultid="16063" heatid="19504" lane="7" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.66" />
                    <SPLIT distance="150" swimtime="00:02:23.42" />
                    <SPLIT distance="200" swimtime="00:03:13.61" />
                    <SPLIT distance="250" swimtime="00:04:09.10" />
                    <SPLIT distance="300" swimtime="00:05:04.85" />
                    <SPLIT distance="350" swimtime="00:05:50.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="250" reactiontime="+93" swimtime="00:01:26.61" resultid="16064" heatid="19514" lane="2" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="295" reactiontime="+90" swimtime="00:00:42.99" resultid="16065" heatid="19542" lane="2" entrytime="00:00:42.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-23" firstname="Krzysztof" gender="M" lastname="Ślęczka" nation="POL" athleteid="16021">
              <RESULTS>
                <RESULT eventid="1079" points="480" reactiontime="+86" swimtime="00:00:25.86" resultid="16022" heatid="19292" lane="1" entrytime="00:00:30.34" />
                <RESULT eventid="1113" points="409" reactiontime="+85" swimtime="00:02:27.64" resultid="16023" heatid="19315" lane="4" entrytime="00:02:34.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.40" />
                    <SPLIT distance="100" swimtime="00:01:10.01" />
                    <SPLIT distance="150" swimtime="00:01:53.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="473" reactiontime="+82" swimtime="00:00:57.64" resultid="16024" heatid="19382" lane="6" entrytime="00:01:04.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="436" reactiontime="+73" swimtime="00:01:06.32" resultid="16025" heatid="19405" lane="2" entrytime="00:01:12.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="439" reactiontime="+81" swimtime="00:01:13.13" resultid="16026" heatid="19440" lane="6" entrytime="00:01:18.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="465" reactiontime="+78" swimtime="00:02:08.21" resultid="16027" heatid="19494" lane="8" entrytime="00:02:14.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.20" />
                    <SPLIT distance="100" swimtime="00:01:01.37" />
                    <SPLIT distance="150" swimtime="00:01:34.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="407" reactiontime="+84" swimtime="00:01:04.86" resultid="16028" heatid="19521" lane="4" entrytime="00:01:11.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="456" reactiontime="+77" swimtime="00:00:32.80" resultid="16029" heatid="19555" lane="4" entrytime="00:00:35.28" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-25" firstname="Artur" gender="M" lastname="Szklarz" nation="POL" athleteid="16039">
              <RESULTS>
                <RESULT eventid="1079" points="371" reactiontime="+78" swimtime="00:00:28.18" resultid="16040" heatid="19294" lane="3" entrytime="00:00:29.04" />
                <RESULT eventid="1113" points="326" reactiontime="+77" swimtime="00:02:39.24" resultid="16041" heatid="19314" lane="8" entrytime="00:02:42.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                    <SPLIT distance="100" swimtime="00:01:17.53" />
                    <SPLIT distance="150" swimtime="00:02:01.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="346" reactiontime="+80" swimtime="00:02:51.51" resultid="16042" heatid="19363" lane="4" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                    <SPLIT distance="100" swimtime="00:01:23.12" />
                    <SPLIT distance="150" swimtime="00:02:07.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="327" reactiontime="+79" swimtime="00:01:12.99" resultid="16043" heatid="19405" lane="7" entrytime="00:01:12.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="359" reactiontime="+81" swimtime="00:01:18.20" resultid="16044" heatid="19439" lane="3" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="348" reactiontime="+78" swimtime="00:00:30.98" resultid="16045" heatid="19458" lane="5" entrytime="00:00:30.90" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="16046" heatid="19520" lane="4" entrytime="00:01:15.00" />
                <RESULT eventid="1681" points="366" reactiontime="+80" swimtime="00:00:35.27" resultid="16047" heatid="19555" lane="3" entrytime="00:00:35.69" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-03-28" firstname="Agata" gender="F" lastname="Meksuła" nation="POL" athleteid="16013">
              <RESULTS>
                <RESULT eventid="1062" points="387" reactiontime="+84" swimtime="00:00:31.89" resultid="16014" heatid="19279" lane="2" entrytime="00:00:35.40" />
                <RESULT eventid="1256" points="362" reactiontime="+81" swimtime="00:01:11.42" resultid="16015" heatid="19371" lane="2" entrytime="00:01:10.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="324" reactiontime="+79" swimtime="00:01:22.46" resultid="16016" heatid="19393" lane="5" entrytime="00:01:22.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="283" reactiontime="+76" swimtime="00:00:37.11" resultid="16017" heatid="19447" lane="7" entrytime="00:00:36.74" />
                <RESULT eventid="1491" points="302" reactiontime="+93" swimtime="00:02:45.09" resultid="16018" heatid="19483" lane="4" entrytime="00:02:38.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.72" />
                    <SPLIT distance="100" swimtime="00:01:17.73" />
                    <SPLIT distance="150" swimtime="00:02:01.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="246" reactiontime="+90" swimtime="00:01:27.11" resultid="16019" heatid="19514" lane="3" entrytime="00:01:25.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="272" reactiontime="+88" swimtime="00:00:44.15" resultid="16020" heatid="19542" lane="1" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-03-14" firstname="Maciej" gender="M" lastname="Kunicki" nation="POL" athleteid="16073">
              <RESULTS>
                <RESULT eventid="1113" points="285" reactiontime="+79" swimtime="00:02:46.52" resultid="16074" heatid="19312" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                    <SPLIT distance="100" swimtime="00:01:16.72" />
                    <SPLIT distance="150" swimtime="00:02:09.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="262" reactiontime="+94" swimtime="00:02:49.59" resultid="16075" heatid="19416" lane="7" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                    <SPLIT distance="100" swimtime="00:01:21.59" />
                    <SPLIT distance="150" swimtime="00:02:06.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="350" reactiontime="+87" swimtime="00:00:30.91" resultid="16076" heatid="19457" lane="9" entrytime="00:00:32.00" />
                <RESULT eventid="1613" points="315" reactiontime="+92" swimtime="00:01:10.59" resultid="16077" heatid="19520" lane="3" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-14" firstname="Piotr" gender="M" lastname="Darowski" nation="POL" athleteid="16066">
              <RESULTS>
                <RESULT eventid="1113" points="405" reactiontime="+79" swimtime="00:02:28.15" resultid="16067" heatid="19317" lane="7" entrytime="00:02:26.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.97" />
                    <SPLIT distance="100" swimtime="00:01:09.71" />
                    <SPLIT distance="150" swimtime="00:01:51.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="448" reactiontime="+78" swimtime="00:02:37.38" resultid="16068" heatid="19365" lane="7" entrytime="00:02:36.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                    <SPLIT distance="100" swimtime="00:01:13.46" />
                    <SPLIT distance="150" swimtime="00:01:54.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="449" reactiontime="+78" swimtime="00:01:12.62" resultid="16069" heatid="19441" lane="5" entrytime="00:01:12.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="384" reactiontime="+75" swimtime="00:05:23.95" resultid="16070" heatid="19512" lane="0" entrytime="00:05:20.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                    <SPLIT distance="100" swimtime="00:01:11.07" />
                    <SPLIT distance="150" swimtime="00:01:54.74" />
                    <SPLIT distance="200" swimtime="00:02:37.63" />
                    <SPLIT distance="250" swimtime="00:03:21.32" />
                    <SPLIT distance="300" swimtime="00:04:06.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="343" reactiontime="+85" swimtime="00:01:08.64" resultid="16071" heatid="19522" lane="5" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="437" reactiontime="+79" swimtime="00:00:33.25" resultid="16072" heatid="19557" lane="3" entrytime="00:00:33.04" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-17" firstname="Sławomir" gender="M" lastname="Kowalski" nation="POL" athleteid="16030">
              <RESULTS>
                <RESULT eventid="1079" points="397" reactiontime="+71" swimtime="00:00:27.56" resultid="16031" heatid="19292" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1113" points="357" reactiontime="+71" swimtime="00:02:34.49" resultid="16032" heatid="19313" lane="8" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.83" />
                    <SPLIT distance="100" swimtime="00:01:15.46" />
                    <SPLIT distance="150" swimtime="00:01:58.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="362" reactiontime="+74" swimtime="00:02:48.98" resultid="16033" heatid="19363" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                    <SPLIT distance="100" swimtime="00:01:20.05" />
                    <SPLIT distance="150" swimtime="00:02:04.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="366" reactiontime="+69" swimtime="00:01:10.29" resultid="16034" heatid="19405" lane="6" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="396" reactiontime="+68" swimtime="00:01:15.70" resultid="16035" heatid="19440" lane="9" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="316" reactiontime="+76" swimtime="00:00:31.98" resultid="16036" heatid="19460" lane="0" entrytime="00:00:30.00" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="16037" heatid="19520" lane="0" entrytime="00:01:20.00" />
                <RESULT eventid="1681" points="395" reactiontime="+66" swimtime="00:00:34.40" resultid="16038" heatid="19556" lane="9" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" points="419" reactiontime="+79" swimtime="00:01:50.36" resultid="16089" heatid="19502" lane="9" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.14" />
                    <SPLIT distance="100" swimtime="00:00:54.22" />
                    <SPLIT distance="150" swimtime="00:01:22.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16021" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="16039" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="16066" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="16030" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="337" reactiontime="+87" swimtime="00:01:58.63" resultid="16090" heatid="19500" lane="5" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                    <SPLIT distance="100" swimtime="00:00:58.40" />
                    <SPLIT distance="150" swimtime="00:01:29.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16082" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="16073" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="16078" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="16048" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" points="391" reactiontime="+66" swimtime="00:02:03.77" resultid="16091" heatid="19423" lane="6" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                    <SPLIT distance="100" swimtime="00:01:07.39" />
                    <SPLIT distance="150" swimtime="00:01:36.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16039" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="16066" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="16021" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="16030" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" points="287" reactiontime="+74" swimtime="00:02:17.14" resultid="16092" heatid="19423" lane="8" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                    <SPLIT distance="100" swimtime="00:01:16.68" />
                    <SPLIT distance="150" swimtime="00:01:48.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16048" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="16078" number="2" reactiontime="+54" />
                    <RELAYPOSITION athleteid="16073" number="3" reactiontime="+60" />
                    <RELAYPOSITION athleteid="16082" number="4" reactiontime="+63" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="424" reactiontime="+85" swimtime="00:01:57.81" resultid="16087" heatid="19322" lane="2" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.65" />
                    <SPLIT distance="100" swimtime="00:00:59.26" />
                    <SPLIT distance="150" swimtime="00:01:30.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16021" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="16057" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="16013" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="16030" number="4" reactiontime="+8" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="375" reactiontime="+80" swimtime="00:02:14.69" resultid="16088" heatid="19563" lane="3" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                    <SPLIT distance="100" swimtime="00:01:04.86" />
                    <SPLIT distance="150" swimtime="00:01:42.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16021" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="16066" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="16057" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="16013" number="4" reactiontime="+63" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="103810" nation="POL" region="10" clubid="14428" name="UKS Dwójka Tczew" name.en="MKS Sambor Tczew" shortname="Dwójka Tczew">
          <ATHLETES>
            <ATHLETE birthdate="1985-07-02" firstname="Jacek" gender="M" lastname="Śliwiński" nation="POL" license="103810700124" athleteid="14429">
              <RESULTS>
                <RESULT eventid="14189" points="534" reactiontime="+78" swimtime="00:09:06.24" resultid="14430" heatid="19618" lane="3" entrytime="00:09:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.60" />
                    <SPLIT distance="100" swimtime="00:01:04.36" />
                    <SPLIT distance="150" swimtime="00:01:38.51" />
                    <SPLIT distance="200" swimtime="00:02:12.51" />
                    <SPLIT distance="250" swimtime="00:02:46.50" />
                    <SPLIT distance="300" swimtime="00:03:20.70" />
                    <SPLIT distance="350" swimtime="00:03:54.97" />
                    <SPLIT distance="400" swimtime="00:04:28.80" />
                    <SPLIT distance="450" swimtime="00:05:02.95" />
                    <SPLIT distance="500" swimtime="00:05:37.61" />
                    <SPLIT distance="550" swimtime="00:06:12.37" />
                    <SPLIT distance="600" swimtime="00:06:47.18" />
                    <SPLIT distance="650" swimtime="00:07:22.00" />
                    <SPLIT distance="700" swimtime="00:07:56.90" />
                    <SPLIT distance="750" swimtime="00:08:31.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00501" nation="POL" region="DOL" clubid="14653" name="UKS Energetyk Zgorzelec">
          <CONTACT city="Zgorzelec" email="biuro@plywanie-zgorzelec.pl" internet="www.plywanie-zgorzelec.pl" name="Kondracki Łukasz" phone="693852488" state="DOL" street="Maratońska" street2="2" zip="59-900" />
          <ATHLETES>
            <ATHLETE birthdate="1948-11-29" firstname="Andrzej" gender="M" lastname="Daszyński" nation="POL" athleteid="14654">
              <RESULTS>
                <RESULT eventid="1113" points="76" reactiontime="+90" swimtime="00:04:18.56" resultid="14655" heatid="19311" lane="9" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.54" />
                    <SPLIT distance="100" swimtime="00:02:04.49" />
                    <SPLIT distance="150" swimtime="00:03:22.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14189" points="91" reactiontime="+89" swimtime="00:16:25.60" resultid="14656" heatid="19614" lane="5" entrytime="00:17:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.62" />
                    <SPLIT distance="100" swimtime="00:01:53.99" />
                    <SPLIT distance="150" swimtime="00:02:54.18" />
                    <SPLIT distance="200" swimtime="00:03:56.37" />
                    <SPLIT distance="250" swimtime="00:04:56.83" />
                    <SPLIT distance="300" swimtime="00:05:57.84" />
                    <SPLIT distance="350" swimtime="00:07:00.64" />
                    <SPLIT distance="400" swimtime="00:08:02.65" />
                    <SPLIT distance="450" swimtime="00:09:05.20" />
                    <SPLIT distance="500" swimtime="00:10:07.96" />
                    <SPLIT distance="550" swimtime="00:11:10.24" />
                    <SPLIT distance="600" swimtime="00:12:12.40" />
                    <SPLIT distance="650" swimtime="00:13:16.03" />
                    <SPLIT distance="700" swimtime="00:14:19.30" />
                    <SPLIT distance="750" swimtime="00:15:23.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="74" reactiontime="+82" swimtime="00:04:46.18" resultid="14657" heatid="19360" lane="0" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.22" />
                    <SPLIT distance="100" swimtime="00:02:19.44" />
                    <SPLIT distance="150" swimtime="00:03:33.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="50" reactiontime="+102" swimtime="00:04:54.41" resultid="14658" heatid="19414" lane="1" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.96" />
                    <SPLIT distance="100" swimtime="00:02:22.86" />
                    <SPLIT distance="150" swimtime="00:03:41.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="82" reactiontime="+85" swimtime="00:01:52.30" resultid="14659" heatid="19472" lane="9" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="79" reactiontime="+105" swimtime="00:09:07.14" resultid="14660" heatid="19507" lane="2" entrytime="00:08:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.35" />
                    <SPLIT distance="100" swimtime="00:02:20.81" />
                    <SPLIT distance="150" swimtime="00:04:32.93" />
                    <SPLIT distance="200" swimtime="00:05:51.86" />
                    <SPLIT distance="250" swimtime="00:07:11.86" />
                    <SPLIT distance="350" swimtime="00:08:10.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="48" reactiontime="+97" swimtime="00:02:11.92" resultid="14661" heatid="19517" lane="8" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="86" reactiontime="+78" swimtime="00:03:58.54" resultid="14662" heatid="19532" lane="5" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.22" />
                    <SPLIT distance="100" swimtime="00:01:57.28" />
                    <SPLIT distance="150" swimtime="00:02:59.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="026" nation="POL" clubid="18474" name="UKS FREGATA Kolbuszowa">
          <CONTACT name="Pietryka" phone="604620876" />
          <ATHLETES>
            <ATHLETE birthdate="1986-07-20" firstname="Bartosz" gender="M" lastname="Pietryka" nation="POL" license="102608700019" athleteid="18475">
              <RESULTS>
                <RESULT eventid="1205" points="331" reactiontime="+80" swimtime="00:00:32.11" resultid="18476" heatid="19352" lane="7" entrytime="00:00:29.20" entrycourse="SCM" />
                <RESULT eventid="1440" points="484" reactiontime="+77" swimtime="00:00:27.75" resultid="18477" heatid="19463" lane="0" entrytime="00:00:27.09" entrycourse="SCM" />
                <RESULT eventid="1613" points="496" reactiontime="+77" swimtime="00:01:00.73" resultid="18478" heatid="19525" lane="0" entrytime="00:01:00.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="MAL" clubid="14435" name="UKS Sp 8 Chrzanów">
          <CONTACT city="Chrzanów" email="abalp@poczta.onet.pl" name="Zabrzański" phone="692076808" state="MAŁ" street="Niepodległości" zip="32 500" />
          <ATHLETES>
            <ATHLETE birthdate="1954-05-12" firstname="Alfred" gender="M" lastname="Zabrzański" nation="POL" athleteid="14436">
              <RESULTS>
                <RESULT eventid="1079" points="270" reactiontime="+93" swimtime="00:00:31.34" resultid="14437" heatid="19291" lane="1" entrytime="00:00:31.60" />
                <RESULT eventid="14189" points="179" reactiontime="+109" swimtime="00:13:05.38" resultid="14438" heatid="19615" lane="4" entrytime="00:13:30.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                    <SPLIT distance="100" swimtime="00:01:27.59" />
                    <SPLIT distance="150" swimtime="00:02:15.50" />
                    <SPLIT distance="200" swimtime="00:03:06.31" />
                    <SPLIT distance="250" swimtime="00:03:56.70" />
                    <SPLIT distance="300" swimtime="00:04:47.62" />
                    <SPLIT distance="350" swimtime="00:05:39.19" />
                    <SPLIT distance="400" swimtime="00:06:30.07" />
                    <SPLIT distance="450" swimtime="00:07:20.60" />
                    <SPLIT distance="500" swimtime="00:08:10.81" />
                    <SPLIT distance="550" swimtime="00:09:00.81" />
                    <SPLIT distance="600" swimtime="00:09:51.04" />
                    <SPLIT distance="650" swimtime="00:10:41.00" />
                    <SPLIT distance="700" swimtime="00:11:30.96" />
                    <SPLIT distance="750" swimtime="00:12:20.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="153" reactiontime="+80" swimtime="00:00:41.48" resultid="14439" heatid="19346" lane="1" entrytime="00:00:41.50" />
                <RESULT eventid="1273" points="245" reactiontime="+91" swimtime="00:01:11.75" resultid="14440" heatid="19379" lane="6" entrytime="00:01:11.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="151" reactiontime="+74" swimtime="00:01:31.69" resultid="14441" heatid="19473" lane="7" entrytime="00:01:30.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="14442" heatid="19489" lane="5" entrytime="00:02:49.00" />
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="14443" heatid="19533" lane="2" entrytime="00:03:29.50" />
                <RESULT eventid="1744" points="190" reactiontime="+104" swimtime="00:06:09.08" resultid="14444" heatid="19701" lane="4" entrytime="00:06:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                    <SPLIT distance="100" swimtime="00:01:22.71" />
                    <SPLIT distance="150" swimtime="00:02:08.71" />
                    <SPLIT distance="200" swimtime="00:02:56.34" />
                    <SPLIT distance="250" swimtime="00:03:44.71" />
                    <SPLIT distance="300" swimtime="00:04:33.41" />
                    <SPLIT distance="350" swimtime="00:05:22.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="1001-11" nation="POL" region="SLA" clubid="16577" name="UKS TRÓJKA Częstochowa">
          <CONTACT city="Częstochowa" email="trojkaczestochowa@o2.pl" name="Gawda" phone="511181791" state="ŚL" street="Schillera" zip="42-200" />
          <ATHLETES>
            <ATHLETE birthdate="1997-08-04" firstname="Wiktoria" gender="F" lastname="Musik" nation="POL" license="100111600053" athleteid="16578">
              <RESULTS>
                <RESULT eventid="1062" points="623" reactiontime="+84" swimtime="00:00:27.20" resultid="16579" heatid="19283" lane="4" entrytime="00:00:27.44" />
                <RESULT eventid="1256" points="632" reactiontime="+83" swimtime="00:00:59.31" resultid="16580" heatid="19372" lane="3" entrytime="00:00:59.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="524" reactiontime="+80" swimtime="00:01:10.28" resultid="16581" heatid="19396" lane="8" entrytime="00:01:11.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="534" reactiontime="+83" swimtime="00:00:30.05" resultid="16582" heatid="19449" lane="6" entrytime="00:00:30.15" />
                <RESULT eventid="1491" points="567" reactiontime="+86" swimtime="00:02:13.83" resultid="16583" heatid="19484" lane="1" entrytime="00:02:28.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.18" />
                    <SPLIT distance="100" swimtime="00:01:04.38" />
                    <SPLIT distance="150" swimtime="00:01:39.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02914" nation="POL" region="MAZ" clubid="18545" name="UKS Victoria Józefów">
          <CONTACT email="ali90@o2.pl" name="kowalczyk alicja" />
          <ATHLETES>
            <ATHLETE birthdate="1966-03-01" firstname="Jan" gender="M" lastname="Kośmider" nation="POL" athleteid="18546">
              <RESULTS>
                <RESULT eventid="1079" points="295" reactiontime="+87" swimtime="00:00:30.41" resultid="18547" heatid="19289" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="18548" heatid="19379" lane="4" entrytime="00:01:10.00" />
                <RESULT eventid="14243" points="283" reactiontime="+82" swimtime="00:01:16.53" resultid="18549" heatid="19402" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="290" reactiontime="+83" swimtime="00:01:23.95" resultid="18550" heatid="19438" lane="9" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="18551" heatid="19552" lane="6" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03311" nation="POL" region="SLA" clubid="17690" name="UKS Wodnik 29 Katowice">
          <CONTACT name="Skoczylas Tomasz" />
          <ATHLETES>
            <ATHLETE birthdate="1958-03-01" firstname="Jan" gender="M" lastname="Wilczek" nation="POL" athleteid="18317">
              <RESULTS>
                <RESULT eventid="1079" points="310" reactiontime="+97" swimtime="00:00:29.93" resultid="18318" heatid="19295" lane="6" entrytime="00:00:29.00" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="18319" heatid="19380" lane="3" entrytime="00:01:08.00" />
                <RESULT eventid="1440" points="313" reactiontime="+105" swimtime="00:00:32.09" resultid="18320" heatid="19456" lane="7" entrytime="00:00:32.50" />
                <RESULT eventid="1613" points="242" reactiontime="+108" swimtime="00:01:17.10" resultid="18321" heatid="19520" lane="2" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-28" firstname="Jerzy" gender="M" lastname="Mroziński" nation="POL" athleteid="18282">
              <RESULTS>
                <RESULT eventid="1239" points="304" reactiontime="+85" swimtime="00:02:59.05" resultid="18283" heatid="19363" lane="3" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.21" />
                    <SPLIT distance="100" swimtime="00:01:24.83" />
                    <SPLIT distance="150" swimtime="00:02:11.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" status="DNS" swimtime="00:00:00.00" resultid="18284" heatid="19403" lane="6" entrytime="00:01:16.00" />
                <RESULT eventid="1406" points="354" reactiontime="+87" swimtime="00:01:18.56" resultid="18285" heatid="19440" lane="7" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="369" reactiontime="+91" swimtime="00:00:35.19" resultid="18286" heatid="19556" lane="2" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-05-08" firstname="Bartłomiej" gender="M" lastname="Kulaga" nation="POL" athleteid="17704">
              <RESULTS>
                <RESULT eventid="1341" points="290" reactiontime="+80" swimtime="00:02:43.95" resultid="17705" heatid="19418" lane="8" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                    <SPLIT distance="100" swimtime="00:01:12.14" />
                    <SPLIT distance="150" swimtime="00:01:54.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="409" reactiontime="+81" swimtime="00:02:13.79" resultid="17706" heatid="19496" lane="1" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.44" />
                    <SPLIT distance="100" swimtime="00:01:04.20" />
                    <SPLIT distance="150" swimtime="00:01:39.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-05-05" firstname="Marek" gender="M" lastname="Mróz" nation="POL" athleteid="17695">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="17696" heatid="19302" lane="6" entrytime="00:00:25.50" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="17697" heatid="19388" lane="0" entrytime="00:00:55.00" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="17698" heatid="19463" lane="5" entrytime="00:00:26.50" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="17699" heatid="19494" lane="4" entrytime="00:02:10.00" />
                <RESULT eventid="14189" status="DNS" swimtime="00:00:00.00" resultid="18952" heatid="19617" lane="1" entrytime="00:10:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-03-09" firstname="Aleksandra" gender="F" lastname="Morkisz" nation="POL" athleteid="17700">
              <RESULTS>
                <RESULT eventid="14225" points="277" reactiontime="+93" swimtime="00:01:26.89" resultid="17701" heatid="19395" lane="1" entrytime="00:01:14.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="312" reactiontime="+92" swimtime="00:01:31.92" resultid="17702" heatid="19431" lane="3" entrytime="00:01:26.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="297" reactiontime="+97" swimtime="00:00:42.89" resultid="17703" heatid="19545" lane="0" entrytime="00:00:37.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-05-16" firstname="Michał" gender="M" lastname="Spławiński" nation="POL" athleteid="17691">
              <RESULTS>
                <RESULT eventid="1079" points="484" reactiontime="+70" swimtime="00:00:25.79" resultid="17692" heatid="19302" lane="8" entrytime="00:00:25.90" />
                <RESULT eventid="1440" points="514" reactiontime="+74" swimtime="00:00:27.20" resultid="17693" heatid="19462" lane="8" entrytime="00:00:27.50" />
                <RESULT eventid="1681" points="561" reactiontime="+80" swimtime="00:00:30.60" resultid="17694" heatid="19558" lane="6" entrytime="00:00:32.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1932-05-18" firstname="Urszula" gender="F" lastname="Walkowicz" nation="POL" athleteid="18308">
              <RESULTS>
                <RESULT eventid="1062" points="25" reactiontime="+136" swimtime="00:01:18.74" resultid="18309" heatid="19275" lane="3" />
                <RESULT eventid="1147" points="29" reactiontime="+119" swimtime="00:25:55.85" resultid="18310" heatid="19594" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.60" />
                    <SPLIT distance="100" swimtime="00:03:03.90" />
                    <SPLIT distance="250" swimtime="00:07:56.37" />
                    <SPLIT distance="450" swimtime="00:14:22.54" />
                    <SPLIT distance="500" swimtime="00:16:05.20" />
                    <SPLIT distance="550" swimtime="00:17:45.21" />
                    <SPLIT distance="600" swimtime="00:19:24.94" />
                    <SPLIT distance="650" swimtime="00:21:02.03" />
                    <SPLIT distance="700" swimtime="00:22:46.14" />
                    <SPLIT distance="750" swimtime="00:24:20.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="35" swimtime="00:01:18.23" resultid="18311" heatid="19336" lane="0" />
                <RESULT eventid="1256" points="24" swimtime="00:02:54.34" resultid="18312" heatid="19367" lane="9" />
                <RESULT eventid="1457" points="29" reactiontime="+98" swimtime="00:02:57.66" resultid="18313" heatid="19465" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:27.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="18314" heatid="19479" lane="6" />
                <RESULT eventid="1630" points="33" reactiontime="+83" swimtime="00:06:08.63" resultid="18315" heatid="19526" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:27.38" />
                    <SPLIT distance="100" swimtime="00:03:02.13" />
                    <SPLIT distance="150" swimtime="00:04:39.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="30" swimtime="00:12:28.44" resultid="18316" heatid="19694" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.72" />
                    <SPLIT distance="100" swimtime="00:02:59.86" />
                    <SPLIT distance="150" swimtime="00:04:33.59" />
                    <SPLIT distance="200" swimtime="00:06:07.98" />
                    <SPLIT distance="250" swimtime="00:07:40.04" />
                    <SPLIT distance="300" swimtime="00:09:11.23" />
                    <SPLIT distance="350" swimtime="00:10:51.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-07-09" firstname="Krystyna" gender="F" lastname="Nicpoń" nation="POL" athleteid="18287">
              <RESULTS>
                <RESULT eventid="1187" points="91" reactiontime="+77" swimtime="00:00:57.04" resultid="18288" heatid="19337" lane="9" entrytime="00:00:55.00" />
                <RESULT eventid="14225" points="69" reactiontime="+109" swimtime="00:02:17.79" resultid="18289" heatid="19390" lane="7" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="85" reactiontime="+95" swimtime="00:02:05.12" resultid="18290" heatid="19466" lane="0" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="94" reactiontime="+77" swimtime="00:04:21.78" resultid="18291" heatid="19527" lane="8" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.43" />
                    <SPLIT distance="100" swimtime="00:02:06.32" />
                    <SPLIT distance="150" swimtime="00:03:15.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-11-14" firstname="Aleksander" gender="M" lastname="Aleksandrowicz" nation="POL" athleteid="18296">
              <RESULTS>
                <RESULT eventid="1079" points="77" reactiontime="+108" swimtime="00:00:47.62" resultid="18297" heatid="19285" lane="0" entrytime="00:00:45.00" />
                <RESULT eventid="1205" points="43" reactiontime="+82" swimtime="00:01:03.08" resultid="18298" heatid="19343" lane="5" entrytime="00:00:56.99" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="18299" heatid="19359" lane="5" entrytime="00:05:32.73" />
                <RESULT comment="K2 - Brak wynurzenia głowy po rozpoczęciu ruchu ramion do wewnątrz z jego najszerszego położenia w drugim cyklu ruchu ramion po starcie lub nawrocie (Time: 16:38)" eventid="1406" reactiontime="+115" status="DSQ" swimtime="00:02:32.83" resultid="18300" heatid="19433" lane="4" entrytime="00:02:36.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="48" reactiontime="+99" swimtime="00:02:14.23" resultid="18301" heatid="19471" lane="6" entrytime="00:02:08.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="50" reactiontime="+78" swimtime="00:04:46.62" resultid="18302" heatid="19532" lane="7" entrytime="00:04:33.15">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:03:34.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="50" reactiontime="+114" swimtime="00:01:08.40" resultid="18303" heatid="19547" lane="1" entrytime="00:01:10.15" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1934-02-02" firstname="Maria" gender="F" lastname="Śmiglewska" nation="POL" athleteid="18304">
              <RESULTS>
                <RESULT eventid="1187" points="29" reactiontime="+148" swimtime="00:01:22.67" resultid="18305" heatid="19336" lane="2" entrytime="00:01:15.00" />
                <RESULT eventid="1388" points="17" swimtime="00:03:58.23" resultid="18306" heatid="19427" lane="6" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:59.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="18" swimtime="00:01:49.21" resultid="18307" heatid="19539" lane="8" entrytime="00:01:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-12-05" firstname="Mariusz" gender="M" lastname="Grelewicz" nation="POL" athleteid="18292">
              <RESULTS>
                <RESULT eventid="1079" points="342" reactiontime="+93" swimtime="00:00:28.95" resultid="18293" heatid="19295" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="1440" points="313" reactiontime="+102" swimtime="00:00:32.08" resultid="18294" heatid="19459" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1681" points="351" reactiontime="+102" swimtime="00:00:35.78" resultid="18295" heatid="19556" lane="3" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-05-15" firstname="Jessica" gender="F" lastname="Thorpe" nation="GBR" athleteid="17707">
              <RESULTS>
                <RESULT eventid="1096" points="381" reactiontime="+111" swimtime="00:02:47.96" resultid="17708" heatid="19309" lane="0" entrytime="00:02:42.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                    <SPLIT distance="100" swimtime="00:01:19.22" />
                    <SPLIT distance="150" swimtime="00:02:07.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="469" reactiontime="+95" swimtime="00:10:16.71" resultid="17709" heatid="19596" lane="4" entrytime="00:09:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.22" />
                    <SPLIT distance="100" swimtime="00:01:11.34" />
                    <SPLIT distance="150" swimtime="00:01:49.44" />
                    <SPLIT distance="200" swimtime="00:02:28.28" />
                    <SPLIT distance="250" swimtime="00:03:07.36" />
                    <SPLIT distance="300" swimtime="00:03:46.52" />
                    <SPLIT distance="350" swimtime="00:04:26.25" />
                    <SPLIT distance="400" swimtime="00:05:05.77" />
                    <SPLIT distance="450" swimtime="00:05:44.39" />
                    <SPLIT distance="500" swimtime="00:06:23.43" />
                    <SPLIT distance="550" swimtime="00:07:02.65" />
                    <SPLIT distance="600" swimtime="00:07:41.73" />
                    <SPLIT distance="650" swimtime="00:08:20.68" />
                    <SPLIT distance="700" swimtime="00:08:59.71" />
                    <SPLIT distance="750" swimtime="00:09:38.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="353" reactiontime="+96" swimtime="00:03:10.27" resultid="17710" heatid="19357" lane="4" entrytime="00:03:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                    <SPLIT distance="100" swimtime="00:01:28.44" />
                    <SPLIT distance="150" swimtime="00:02:18.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" status="DNS" swimtime="00:00:00.00" resultid="17711" heatid="19394" lane="5" entrytime="00:01:15.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-04-22" firstname="Tomasz" gender="M" lastname="Skoczylas" nation="POL" athleteid="18273">
              <RESULTS>
                <RESULT eventid="1079" points="339" reactiontime="+97" swimtime="00:00:29.03" resultid="18274" heatid="19295" lane="2" entrytime="00:00:29.00" />
                <RESULT eventid="14207" points="286" reactiontime="+117" swimtime="00:21:26.06" resultid="18275" heatid="19622" lane="3" entrytime="00:21:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                    <SPLIT distance="100" swimtime="00:01:14.76" />
                    <SPLIT distance="150" swimtime="00:01:55.74" />
                    <SPLIT distance="200" swimtime="00:02:36.98" />
                    <SPLIT distance="250" swimtime="00:03:19.11" />
                    <SPLIT distance="300" swimtime="00:04:01.52" />
                    <SPLIT distance="350" swimtime="00:04:44.48" />
                    <SPLIT distance="400" swimtime="00:05:29.61" />
                    <SPLIT distance="450" swimtime="00:06:12.94" />
                    <SPLIT distance="500" swimtime="00:06:55.89" />
                    <SPLIT distance="550" swimtime="00:07:38.44" />
                    <SPLIT distance="600" swimtime="00:08:21.56" />
                    <SPLIT distance="650" swimtime="00:09:04.12" />
                    <SPLIT distance="700" swimtime="00:09:47.07" />
                    <SPLIT distance="750" swimtime="00:10:30.11" />
                    <SPLIT distance="800" swimtime="00:11:13.32" />
                    <SPLIT distance="850" swimtime="00:11:56.47" />
                    <SPLIT distance="900" swimtime="00:12:39.83" />
                    <SPLIT distance="950" swimtime="00:13:22.96" />
                    <SPLIT distance="1000" swimtime="00:14:06.60" />
                    <SPLIT distance="1050" swimtime="00:14:49.76" />
                    <SPLIT distance="1100" swimtime="00:15:33.23" />
                    <SPLIT distance="1150" swimtime="00:16:17.08" />
                    <SPLIT distance="1200" swimtime="00:17:00.78" />
                    <SPLIT distance="1250" swimtime="00:17:44.32" />
                    <SPLIT distance="1300" swimtime="00:18:28.25" />
                    <SPLIT distance="1350" swimtime="00:19:12.70" />
                    <SPLIT distance="1400" swimtime="00:19:57.33" />
                    <SPLIT distance="1450" swimtime="00:20:41.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="238" reactiontime="+90" swimtime="00:00:35.83" resultid="18276" heatid="19348" lane="0" entrytime="00:00:36.00" />
                <RESULT eventid="1273" points="331" reactiontime="+93" swimtime="00:01:04.93" resultid="18277" heatid="19382" lane="3" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="249" reactiontime="+94" swimtime="00:01:17.68" resultid="18278" heatid="19474" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="294" reactiontime="+97" swimtime="00:02:29.42" resultid="18279" heatid="19492" lane="8" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.98" />
                    <SPLIT distance="100" swimtime="00:01:11.21" />
                    <SPLIT distance="150" swimtime="00:01:49.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="229" reactiontime="+95" swimtime="00:02:52.52" resultid="18280" heatid="19534" lane="3" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                    <SPLIT distance="100" swimtime="00:01:24.50" />
                    <SPLIT distance="150" swimtime="00:02:09.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="319" reactiontime="+100" swimtime="00:05:10.56" resultid="18281" heatid="19704" lane="4" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.51" />
                    <SPLIT distance="100" swimtime="00:01:11.75" />
                    <SPLIT distance="150" swimtime="00:01:50.39" />
                    <SPLIT distance="200" swimtime="00:02:29.57" />
                    <SPLIT distance="250" swimtime="00:03:08.93" />
                    <SPLIT distance="300" swimtime="00:03:48.93" />
                    <SPLIT distance="350" swimtime="00:04:29.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-02-23" firstname="Paweł" gender="M" lastname="Bobeł" nation="POL" athleteid="17712">
              <RESULTS>
                <RESULT eventid="1205" points="277" reactiontime="+63" swimtime="00:00:34.05" resultid="17713" heatid="19347" lane="6" entrytime="00:00:37.15" />
                <RESULT eventid="14243" points="278" reactiontime="+82" swimtime="00:01:17.03" resultid="17714" heatid="19405" lane="9" entrytime="00:01:13.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="295" reactiontime="+84" swimtime="00:01:23.49" resultid="17715" heatid="19440" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="278" reactiontime="+67" swimtime="00:01:14.90" resultid="17716" heatid="19476" lane="0" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-19" firstname="Krzysztof" gender="M" lastname="Kulczyk" nation="POL" athleteid="18264">
              <RESULTS>
                <RESULT eventid="1079" points="211" reactiontime="+120" swimtime="00:00:34.03" resultid="18265" heatid="19289" lane="1" entrytime="00:00:33.50" />
                <RESULT eventid="1113" points="145" reactiontime="+102" swimtime="00:03:28.25" resultid="18266" heatid="19311" lane="3" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.23" />
                    <SPLIT distance="100" swimtime="00:01:31.64" />
                    <SPLIT distance="150" swimtime="00:02:40.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="153" reactiontime="+94" swimtime="00:00:41.49" resultid="18267" heatid="19345" lane="5" entrytime="00:00:43.00" />
                <RESULT eventid="1341" points="116" reactiontime="+108" swimtime="00:03:41.98" resultid="18268" heatid="19415" lane="8" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.60" />
                    <SPLIT distance="100" swimtime="00:01:42.85" />
                    <SPLIT distance="150" swimtime="00:02:43.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="244" reactiontime="+103" swimtime="00:00:34.88" resultid="18269" heatid="19453" lane="5" entrytime="00:00:36.50" />
                <RESULT eventid="1474" points="155" reactiontime="+88" swimtime="00:01:30.97" resultid="18270" heatid="19473" lane="0" entrytime="00:01:34.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="155" reactiontime="+107" swimtime="00:01:29.44" resultid="18271" heatid="19519" lane="0" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="141" reactiontime="+88" swimtime="00:03:22.88" resultid="18272" heatid="19533" lane="6" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.06" />
                    <SPLIT distance="100" swimtime="00:01:38.59" />
                    <SPLIT distance="150" swimtime="00:02:32.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" points="350" reactiontime="+98" swimtime="00:01:57.17" resultid="18322" heatid="19500" lane="6" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.26" />
                    <SPLIT distance="100" swimtime="00:00:59.90" />
                    <SPLIT distance="150" swimtime="00:01:29.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18292" number="1" reactiontime="+98" />
                    <RELAYPOSITION athleteid="18282" number="2" reactiontime="+43" />
                    <RELAYPOSITION athleteid="18317" number="3" reactiontime="+29" />
                    <RELAYPOSITION athleteid="18273" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1548" status="DNS" swimtime="00:00:00.00" resultid="17719" heatid="19501" lane="7" entrytime="00:01:55.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17712" number="1" />
                    <RELAYPOSITION athleteid="17695" number="2" />
                    <RELAYPOSITION athleteid="17691" number="3" />
                    <RELAYPOSITION athleteid="17704" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" status="DNS" swimtime="00:00:00.00" resultid="17717" heatid="19321" lane="6" entrytime="00:02:00.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17700" number="1" />
                    <RELAYPOSITION athleteid="17691" number="2" />
                    <RELAYPOSITION athleteid="17695" number="3" />
                    <RELAYPOSITION athleteid="17707" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1698" status="DNS" swimtime="00:00:00.00" resultid="17718" heatid="19562" lane="2" entrytime="00:02:30.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17704" number="1" />
                    <RELAYPOSITION athleteid="17700" number="2" />
                    <RELAYPOSITION athleteid="17712" number="3" />
                    <RELAYPOSITION athleteid="17707" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="01711" nation="POL" region="11" clubid="14346" name="UKS WODNIK Siemianowice Ślaskie" shortname="UKS WODNIK Siemianowice Ślaski">
          <CONTACT city="Siemianowice Śląskie" email="vivisektor@interia.pl" name="Małyszek Leszek" phone="534033934" state="ŚLĄSK" street="Mikołaja 3" zip="41-106" />
          <ATHLETES>
            <ATHLETE birthdate="1960-02-18" firstname="Piotr" gender="M" lastname="Szymik" nation="POL" athleteid="14347">
              <RESULTS>
                <RESULT eventid="1113" points="204" reactiontime="+88" swimtime="00:03:06.00" resultid="14348" heatid="19311" lane="4" entrytime="00:03:12.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.89" />
                    <SPLIT distance="100" swimtime="00:01:28.30" />
                    <SPLIT distance="150" swimtime="00:02:22.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14207" points="237" reactiontime="+86" swimtime="00:22:49.58" resultid="14349" heatid="19621" lane="3" entrytime="00:23:10.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                    <SPLIT distance="100" swimtime="00:01:21.82" />
                    <SPLIT distance="150" swimtime="00:02:07.51" />
                    <SPLIT distance="200" swimtime="00:02:53.42" />
                    <SPLIT distance="250" swimtime="00:03:39.82" />
                    <SPLIT distance="300" swimtime="00:04:26.14" />
                    <SPLIT distance="350" swimtime="00:05:12.59" />
                    <SPLIT distance="400" swimtime="00:05:58.89" />
                    <SPLIT distance="450" swimtime="00:06:45.40" />
                    <SPLIT distance="500" swimtime="00:07:31.23" />
                    <SPLIT distance="550" swimtime="00:08:17.31" />
                    <SPLIT distance="600" swimtime="00:09:03.06" />
                    <SPLIT distance="650" swimtime="00:09:49.01" />
                    <SPLIT distance="700" swimtime="00:10:34.11" />
                    <SPLIT distance="750" swimtime="00:11:19.85" />
                    <SPLIT distance="800" swimtime="00:12:06.02" />
                    <SPLIT distance="850" swimtime="00:12:52.97" />
                    <SPLIT distance="900" swimtime="00:13:39.39" />
                    <SPLIT distance="950" swimtime="00:14:25.42" />
                    <SPLIT distance="1000" swimtime="00:15:11.87" />
                    <SPLIT distance="1050" swimtime="00:15:58.11" />
                    <SPLIT distance="1100" swimtime="00:16:44.38" />
                    <SPLIT distance="1150" swimtime="00:17:31.09" />
                    <SPLIT distance="1200" swimtime="00:18:17.27" />
                    <SPLIT distance="1250" swimtime="00:19:02.70" />
                    <SPLIT distance="1300" swimtime="00:19:49.38" />
                    <SPLIT distance="1350" swimtime="00:20:36.04" />
                    <SPLIT distance="1400" swimtime="00:21:21.83" />
                    <SPLIT distance="1450" swimtime="00:22:06.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="128" reactiontime="+77" swimtime="00:03:35.01" resultid="14350" heatid="19415" lane="7" entrytime="00:03:21.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.84" />
                    <SPLIT distance="100" swimtime="00:01:39.16" />
                    <SPLIT distance="150" swimtime="00:02:38.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="203" reactiontime="+85" swimtime="00:00:37.06" resultid="14351" heatid="19453" lane="4" entrytime="00:00:36.23" />
                <RESULT eventid="1578" points="202" reactiontime="+89" swimtime="00:06:40.84" resultid="14352" heatid="19509" lane="1" entrytime="00:06:30.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.25" />
                    <SPLIT distance="100" swimtime="00:01:37.02" />
                    <SPLIT distance="150" swimtime="00:02:27.52" />
                    <SPLIT distance="200" swimtime="00:03:18.56" />
                    <SPLIT distance="250" swimtime="00:04:16.35" />
                    <SPLIT distance="300" swimtime="00:05:14.73" />
                    <SPLIT distance="350" swimtime="00:05:59.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="14353" heatid="19519" lane="2" entrytime="00:01:28.30" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="14354" heatid="19703" lane="2" entrytime="00:05:51.12" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01006" nation="POL" region="06" clubid="14596" name="Unia Oświęcim Masters">
          <ATHLETES>
            <ATHLETE birthdate="1961-03-16" firstname="Tomasz" gender="M" lastname="Dorywalski" nation="POL" license="101006700340" athleteid="14597">
              <RESULTS>
                <RESULT eventid="1205" points="201" reactiontime="+77" swimtime="00:00:37.92" resultid="14598" heatid="19346" lane="2" entrytime="00:00:40.50" />
                <RESULT eventid="1474" points="205" reactiontime="+75" swimtime="00:01:22.90" resultid="14599" heatid="19474" lane="2" entrytime="00:01:22.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="201" reactiontime="+81" swimtime="00:03:00.17" resultid="14600" heatid="19534" lane="2" entrytime="00:03:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.54" />
                    <SPLIT distance="100" swimtime="00:01:25.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="URWAR" nation="POL" region="WAR" clubid="17561" name="Ursynów Masters">
          <CONTACT city="WARSZAWA" name="MICHAŁ NOWAK" />
          <ATHLETES>
            <ATHLETE birthdate="1970-01-23" firstname="Michał" gender="M" lastname="Rybarczyk" nation="POL" athleteid="17562">
              <RESULTS>
                <RESULT eventid="1079" points="351" reactiontime="+87" swimtime="00:00:28.70" resultid="17563" heatid="19295" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="1205" points="124" reactiontime="+80" swimtime="00:00:44.51" resultid="17564" heatid="19346" lane="0" entrytime="00:00:42.00" />
                <RESULT eventid="1273" points="335" reactiontime="+80" swimtime="00:01:04.68" resultid="17565" heatid="19382" lane="9" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="274" reactiontime="+77" swimtime="00:00:33.55" resultid="17566" heatid="19456" lane="9" entrytime="00:00:33.00" />
                <RESULT eventid="1508" points="287" reactiontime="+85" swimtime="00:02:30.57" resultid="17567" heatid="19491" lane="7" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                    <SPLIT distance="100" swimtime="00:01:12.23" />
                    <SPLIT distance="150" swimtime="00:01:52.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="17568" heatid="19519" lane="4" entrytime="00:01:25.00" />
                <RESULT eventid="1744" points="275" reactiontime="+80" swimtime="00:05:26.07" resultid="17569" heatid="19704" lane="9" entrytime="00:05:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="100" swimtime="00:01:14.28" />
                    <SPLIT distance="150" swimtime="00:01:55.91" />
                    <SPLIT distance="200" swimtime="00:02:39.17" />
                    <SPLIT distance="250" swimtime="00:03:22.56" />
                    <SPLIT distance="300" swimtime="00:04:04.37" />
                    <SPLIT distance="350" swimtime="00:04:47.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="031/05" nation="POL" region="LOD" clubid="15072" name="UTW&quot;Masters&quot;Zgierz">
          <CONTACT city="ZGIERZ" email="roman.wiczel@gmail.com" name="WICZEL" phone="691-928-922" state="ŁÓDZK" street="ŁĘCZYCKA 24" zip="95-100" />
          <ATHLETES>
            <ATHLETE birthdate="1955-03-16" firstname="Janusz" gender="M" lastname="Błasiak" nation="POL" license="503105700050" athleteid="15253">
              <RESULTS>
                <RESULT eventid="1079" points="132" swimtime="00:00:39.76" resultid="15254" heatid="19286" lane="1" entrytime="00:00:39.88" entrycourse="SCM" />
                <RESULT eventid="1113" points="81" reactiontime="+94" swimtime="00:04:12.67" resultid="15255" heatid="19310" lane="7" entrytime="00:04:20.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.20" />
                    <SPLIT distance="100" swimtime="00:02:05.83" />
                    <SPLIT distance="150" swimtime="00:03:23.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="121" reactiontime="+102" swimtime="00:01:30.77" resultid="15256" heatid="19375" lane="4" entrytime="00:01:31.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="44" reactiontime="+108" swimtime="00:05:07.49" resultid="15257" heatid="19414" lane="9" entrytime="00:04:58.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.46" />
                    <SPLIT distance="100" swimtime="00:02:25.94" />
                    <SPLIT distance="150" swimtime="00:03:50.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="101" reactiontime="+99" swimtime="00:03:33.03" resultid="15258" heatid="19487" lane="8" entrytime="00:03:32.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.50" />
                    <SPLIT distance="100" swimtime="00:01:44.37" />
                    <SPLIT distance="150" swimtime="00:02:42.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="81" reactiontime="+104" swimtime="00:09:04.21" resultid="15259" heatid="19507" lane="7" entrytime="00:09:09.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.46" />
                    <SPLIT distance="100" swimtime="00:02:17.38" />
                    <SPLIT distance="150" swimtime="00:03:29.33" />
                    <SPLIT distance="200" swimtime="00:06:00.31" />
                    <SPLIT distance="250" swimtime="00:07:19.28" />
                    <SPLIT distance="350" swimtime="00:08:13.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="51" reactiontime="+102" swimtime="00:02:08.88" resultid="15260" heatid="19517" lane="7" entrytime="00:02:06.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="61" reactiontime="+92" swimtime="00:04:27.09" resultid="15261" heatid="19532" lane="9" entrytime="00:04:47.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.43" />
                    <SPLIT distance="100" swimtime="00:02:13.71" />
                    <SPLIT distance="150" swimtime="00:03:22.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-07-28" firstname="Natalia" gender="F" lastname="Szczęsnowicz" nation="POL" license="503105600052" athleteid="15300">
              <RESULTS>
                <RESULT eventid="1664" points="462" reactiontime="+81" swimtime="00:00:37.03" resultid="15301" heatid="19544" lane="4" entrytime="00:00:38.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-18" firstname="Daria" gender="F" lastname="Fajkowska" nation="POL" license="503105600018" athleteid="15281">
              <RESULTS>
                <RESULT eventid="1096" points="463" reactiontime="+102" swimtime="00:02:37.43" resultid="15282" heatid="19306" lane="3" entrytime="00:03:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.80" />
                    <SPLIT distance="100" swimtime="00:01:12.31" />
                    <SPLIT distance="150" swimtime="00:01:58.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="470" reactiontime="+83" swimtime="00:00:33.00" resultid="15283" heatid="19341" lane="8" entrytime="00:00:33.10" entrycourse="SCM" />
                <RESULT eventid="14225" points="499" reactiontime="+91" swimtime="00:01:11.42" resultid="15284" heatid="19395" lane="4" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="421" reactiontime="+76" swimtime="00:02:38.97" resultid="15285" heatid="19529" lane="1" entrytime="00:02:43.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.72" />
                    <SPLIT distance="100" swimtime="00:01:16.94" />
                    <SPLIT distance="150" swimtime="00:01:57.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-12" firstname="Małgorzata" gender="F" lastname="Ścibiorek" nation="POL" license="503105600028" athleteid="15235">
              <RESULTS>
                <RESULT eventid="1096" points="441" reactiontime="+86" swimtime="00:02:40.07" resultid="15236" heatid="19308" lane="2" entrytime="00:02:53.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                    <SPLIT distance="100" swimtime="00:01:14.50" />
                    <SPLIT distance="150" swimtime="00:02:02.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="368" reactiontime="+73" swimtime="00:00:35.79" resultid="15237" heatid="19340" lane="6" entrytime="00:00:35.40" entrycourse="SCM" />
                <RESULT eventid="14225" points="448" reactiontime="+83" swimtime="00:01:14.05" resultid="15238" heatid="19395" lane="6" entrytime="00:01:13.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="437" reactiontime="+81" swimtime="00:00:32.12" resultid="15239" heatid="19449" lane="9" entrytime="00:00:32.20" entrycourse="SCM" />
                <RESULT eventid="1457" points="338" reactiontime="+77" swimtime="00:01:18.99" resultid="15240" heatid="19468" lane="5" entrytime="00:01:14.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="459" swimtime="00:01:10.77" resultid="15241" heatid="19515" lane="6" entrytime="00:01:14.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-09" firstname="Włodzimierz" gender="M" lastname="Przytulski" nation="POL" license="503105700027" athleteid="15246">
              <RESULTS>
                <RESULT eventid="1205" points="237" reactiontime="+72" swimtime="00:00:35.89" resultid="15247" heatid="19348" lane="7" entrytime="00:00:36.00" entrycourse="SCM" />
                <RESULT eventid="1341" points="200" reactiontime="+92" swimtime="00:03:05.59" resultid="15248" heatid="19416" lane="9" entrytime="00:03:08.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.31" />
                    <SPLIT distance="100" swimtime="00:01:28.61" />
                    <SPLIT distance="150" swimtime="00:02:17.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="288" reactiontime="+90" swimtime="00:00:32.98" resultid="15249" heatid="19456" lane="2" entrytime="00:00:32.50" entrycourse="SCM" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="15250" heatid="19509" lane="0" entrytime="00:06:35.00" entrycourse="SCM" />
                <RESULT eventid="1613" points="218" reactiontime="+100" swimtime="00:01:19.79" resultid="15251" heatid="19520" lane="1" entrytime="00:01:18.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="15252" heatid="19703" lane="4" entrytime="00:05:40.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-04-16" firstname="Krzysztof" gender="M" lastname="Gawłowicz" nation="POL" license="503105700049" athleteid="15274">
              <RESULTS>
                <RESULT eventid="1079" points="503" reactiontime="+71" swimtime="00:00:25.47" resultid="15275" heatid="19303" lane="7" entrytime="00:00:24.99" entrycourse="SCM" />
                <RESULT eventid="1440" points="528" reactiontime="+74" swimtime="00:00:26.96" resultid="15276" heatid="19463" lane="3" entrytime="00:00:26.50" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-05-12" firstname="Tadeusz" gender="M" lastname="Obiedziński" nation="POL" license="503105700038" athleteid="15277">
              <RESULTS>
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="15278" heatid="19360" lane="5" entrytime="00:03:40.00" entrycourse="SCM" />
                <RESULT eventid="1406" points="188" reactiontime="+111" swimtime="00:01:37.04" resultid="15279" heatid="19436" lane="3" entrytime="00:01:33.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="223" reactiontime="+94" swimtime="00:00:41.58" resultid="15280" heatid="19551" lane="9" entrytime="00:00:42.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-07" firstname="Ewa" gender="F" lastname="Stępień" nation="POL" license="503105600029" athleteid="15242">
              <RESULTS>
                <RESULT eventid="1256" points="278" reactiontime="+83" swimtime="00:01:18.00" resultid="15243" heatid="19371" lane="1" entrytime="00:01:14.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="315" reactiontime="+75" swimtime="00:01:31.65" resultid="15244" heatid="19430" lane="4" entrytime="00:01:31.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="333" reactiontime="+75" swimtime="00:00:41.30" resultid="15245" heatid="19543" lane="8" entrytime="00:00:40.40" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-03" firstname="Urszula" gender="F" lastname="Mróz" nation="POL" license="503105600030" athleteid="15222">
              <RESULTS>
                <RESULT eventid="1062" points="360" reactiontime="+92" swimtime="00:00:32.66" resultid="15223" heatid="19281" lane="6" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1187" points="318" reactiontime="+77" swimtime="00:00:37.60" resultid="15224" heatid="19339" lane="5" entrytime="00:00:38.00" entrycourse="SCM" />
                <RESULT eventid="1324" points="226" reactiontime="+101" swimtime="00:03:16.35" resultid="15225" heatid="19412" lane="7" entrytime="00:03:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.73" />
                    <SPLIT distance="100" swimtime="00:01:38.33" />
                    <SPLIT distance="150" swimtime="00:02:29.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="346" reactiontime="+92" swimtime="00:00:34.70" resultid="15226" heatid="19447" lane="6" entrytime="00:00:36.30" entrycourse="SCM" />
                <RESULT eventid="1457" points="261" reactiontime="+78" swimtime="00:01:26.08" resultid="15227" heatid="19467" lane="5" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="283" reactiontime="+94" swimtime="00:01:23.11" resultid="15228" heatid="19515" lane="7" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-05-03" firstname="Stanisław" gender="M" lastname="Sikorski" nation="POL" license="503105700054" athleteid="15286">
              <RESULTS>
                <RESULT eventid="1205" points="64" reactiontime="+105" swimtime="00:00:55.31" resultid="15287" heatid="19344" lane="3" entrytime="00:00:50.00" entrycourse="SCM" />
                <RESULT eventid="1406" points="82" reactiontime="+123" swimtime="00:02:07.83" resultid="15288" heatid="19434" lane="8" entrytime="00:02:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="15289" heatid="19471" lane="0" entrytime="00:02:20.00" entrycourse="SCM" />
                <RESULT eventid="1681" points="112" reactiontime="+137" swimtime="00:00:52.32" resultid="15290" heatid="19548" lane="2" entrytime="00:00:54.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-06-10" firstname="Sonia" gender="F" lastname="Bochyńska" nation="POL" license="503105600046" athleteid="15229">
              <RESULTS>
                <RESULT eventid="1062" points="585" reactiontime="+79" swimtime="00:00:27.78" resultid="15230" heatid="19283" lane="2" entrytime="00:00:28.00" entrycourse="SCM" />
                <RESULT eventid="1187" points="562" reactiontime="+65" swimtime="00:00:31.10" resultid="15231" heatid="19341" lane="2" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1256" points="564" reactiontime="+70" swimtime="00:01:01.60" resultid="15232" heatid="19372" lane="7" entrytime="00:01:01.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" status="DNS" swimtime="00:00:00.00" resultid="15233" heatid="19449" lane="2" entrytime="00:00:30.50" entrycourse="SCM" />
                <RESULT eventid="1457" points="536" reactiontime="+69" swimtime="00:01:07.71" resultid="15234" heatid="19469" lane="5" entrytime="00:01:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-22" firstname="Roman" gender="M" lastname="Wiczel" nation="POL" license="503105700034" athleteid="15214">
              <RESULTS>
                <RESULT eventid="14189" points="112" reactiontime="+106" swimtime="00:15:18.39" resultid="15215" heatid="19614" lane="4" entrytime="00:16:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.93" />
                    <SPLIT distance="100" swimtime="00:01:45.15" />
                    <SPLIT distance="150" swimtime="00:02:44.58" />
                    <SPLIT distance="200" swimtime="00:03:42.50" />
                    <SPLIT distance="300" swimtime="00:05:38.13" />
                    <SPLIT distance="350" swimtime="00:06:35.52" />
                    <SPLIT distance="400" swimtime="00:08:31.16" />
                    <SPLIT distance="500" swimtime="00:09:30.50" />
                    <SPLIT distance="550" swimtime="00:10:29.35" />
                    <SPLIT distance="700" swimtime="00:13:27.76" />
                    <SPLIT distance="750" swimtime="00:14:28.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="130" swimtime="00:00:43.78" resultid="15216" heatid="19345" lane="0" entrytime="00:00:45.00" entrycourse="SCM" />
                <RESULT eventid="1239" points="195" reactiontime="+99" swimtime="00:03:27.53" resultid="15217" heatid="19361" lane="8" entrytime="00:03:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.27" />
                    <SPLIT distance="100" swimtime="00:01:42.22" />
                    <SPLIT distance="150" swimtime="00:02:37.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="209" reactiontime="+100" swimtime="00:01:33.68" resultid="15218" heatid="19436" lane="4" entrytime="00:01:31.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="129" reactiontime="+80" swimtime="00:01:36.63" resultid="15219" heatid="19472" lane="3" entrytime="00:01:39.00" entrycourse="SCM" />
                <RESULT eventid="1681" points="230" reactiontime="+95" swimtime="00:00:41.17" resultid="15220" heatid="19551" lane="7" entrytime="00:00:41.00" entrycourse="SCM" />
                <RESULT eventid="1744" points="116" reactiontime="+100" swimtime="00:07:14.96" resultid="15221" heatid="19700" lane="8" entrytime="00:07:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.49" />
                    <SPLIT distance="100" swimtime="00:01:41.95" />
                    <SPLIT distance="150" swimtime="00:02:38.59" />
                    <SPLIT distance="200" swimtime="00:03:34.42" />
                    <SPLIT distance="250" swimtime="00:04:30.86" />
                    <SPLIT distance="300" swimtime="00:05:26.09" />
                    <SPLIT distance="350" swimtime="00:06:20.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-03-01" firstname="Waldemar" gender="M" lastname="Jagiełło" nation="POL" license="503105700036" athleteid="15291">
              <RESULTS>
                <RESULT eventid="1079" points="493" reactiontime="+83" swimtime="00:00:25.63" resultid="15292" heatid="19300" lane="9" entrytime="00:00:26.70" entrycourse="SCM" />
                <RESULT eventid="1113" points="427" reactiontime="+92" swimtime="00:02:25.50" resultid="15293" heatid="19315" lane="3" entrytime="00:02:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.07" />
                    <SPLIT distance="100" swimtime="00:01:09.04" />
                    <SPLIT distance="150" swimtime="00:01:51.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="376" reactiontime="+46" swimtime="00:00:30.77" resultid="15294" heatid="19350" lane="7" entrytime="00:00:32.10" entrycourse="SCM" />
                <RESULT eventid="14243" points="478" reactiontime="+83" swimtime="00:01:04.31" resultid="15295" heatid="19409" lane="9" entrytime="00:01:04.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="458" reactiontime="+90" swimtime="00:01:12.14" resultid="15296" heatid="19441" lane="1" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="423" reactiontime="+86" swimtime="00:00:29.02" resultid="15297" heatid="19461" lane="3" entrytime="00:00:28.50" entrycourse="SCM" />
                <RESULT eventid="1613" points="343" reactiontime="+95" swimtime="00:01:08.65" resultid="15298" heatid="19522" lane="4" entrytime="00:01:09.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="488" reactiontime="+80" swimtime="00:00:32.07" resultid="15299" heatid="19559" lane="9" entrytime="00:00:32.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-12-03" firstname="Zbigniew" gender="M" lastname="Maciejczyk" nation="POL" license="503105700026" athleteid="15262">
              <RESULTS>
                <RESULT eventid="1079" points="223" swimtime="00:00:33.40" resultid="15263" heatid="19289" lane="9" entrytime="00:00:34.00" entrycourse="SCM" />
                <RESULT eventid="1273" points="189" reactiontime="+96" swimtime="00:01:18.29" resultid="15264" heatid="19378" lane="9" entrytime="00:01:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="70" reactiontime="+107" swimtime="00:04:22.59" resultid="15265" heatid="19414" lane="7" entrytime="00:04:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.77" />
                    <SPLIT distance="100" swimtime="00:02:15.41" />
                    <SPLIT distance="150" swimtime="00:03:28.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="174" reactiontime="+105" swimtime="00:00:38.99" resultid="15266" heatid="19453" lane="0" entrytime="00:00:38.00" entrycourse="SCM" />
                <RESULT eventid="1613" points="108" reactiontime="+103" swimtime="00:01:40.89" resultid="15267" heatid="19518" lane="7" entrytime="00:01:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="127" reactiontime="+101" swimtime="00:07:01.32" resultid="15268" heatid="19700" lane="3" entrytime="00:07:14.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.28" />
                    <SPLIT distance="100" swimtime="00:01:40.11" />
                    <SPLIT distance="150" swimtime="00:02:35.72" />
                    <SPLIT distance="200" swimtime="00:03:32.50" />
                    <SPLIT distance="250" swimtime="00:04:27.79" />
                    <SPLIT distance="300" swimtime="00:05:22.17" />
                    <SPLIT distance="350" swimtime="00:06:15.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-03-23" firstname="Tomasz" gender="M" lastname="Cajdler" nation="POL" license="503105700035" athleteid="15269">
              <RESULTS>
                <RESULT eventid="1079" points="244" reactiontime="+107" swimtime="00:00:32.39" resultid="15270" heatid="19289" lane="3" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1273" points="188" reactiontime="+109" swimtime="00:01:18.37" resultid="15271" heatid="19378" lane="2" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="167" reactiontime="+100" swimtime="00:01:40.92" resultid="15272" heatid="19436" lane="7" entrytime="00:01:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="192" reactiontime="+91" swimtime="00:00:43.70" resultid="15273" heatid="19551" lane="6" entrytime="00:00:40.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" points="234" reactiontime="+88" swimtime="00:02:13.99" resultid="15307" heatid="19500" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.73" />
                    <SPLIT distance="100" swimtime="00:01:05.25" />
                    <SPLIT distance="150" swimtime="00:01:49.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15291" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="15214" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="15286" number="3" reactiontime="+94" />
                    <RELAYPOSITION athleteid="15274" number="4" reactiontime="+12" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" status="DNS" swimtime="00:00:00.00" resultid="15308" heatid="19422" lane="2" entrytime="00:02:18.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15291" number="1" />
                    <RELAYPOSITION athleteid="15214" number="2" />
                    <RELAYPOSITION athleteid="15274" number="3" />
                    <RELAYPOSITION athleteid="15253" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1548" points="223" reactiontime="+87" swimtime="00:02:16.16" resultid="15309" heatid="19500" lane="8" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                    <SPLIT distance="100" swimtime="00:01:10.77" />
                    <SPLIT distance="150" swimtime="00:01:45.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15269" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="15277" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="15262" number="3" reactiontime="+83" />
                    <RELAYPOSITION athleteid="15246" number="4" reactiontime="+68" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" points="200" reactiontime="+75" swimtime="00:02:34.54" resultid="15310" heatid="19422" lane="8" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.57" />
                    <SPLIT distance="100" swimtime="00:01:19.01" />
                    <SPLIT distance="150" swimtime="00:01:59.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15246" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="15277" number="2" reactiontime="+75" />
                    <RELAYPOSITION athleteid="15262" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="15269" number="4" reactiontime="+117" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1525" points="411" reactiontime="+87" swimtime="00:02:06.74" resultid="15305" heatid="19498" lane="7" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                    <SPLIT distance="100" swimtime="00:01:03.78" />
                    <SPLIT distance="150" swimtime="00:01:37.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15235" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="15222" number="2" reactiontime="+80" />
                    <RELAYPOSITION athleteid="15242" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="15281" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1358" points="415" reactiontime="+86" swimtime="00:02:18.35" resultid="15306" heatid="19420" lane="5" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                    <SPLIT distance="100" swimtime="00:01:13.44" />
                    <SPLIT distance="150" swimtime="00:01:47.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15281" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="15242" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="15222" number="3" reactiontime="+75" />
                    <RELAYPOSITION athleteid="15235" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="442" reactiontime="+83" swimtime="00:01:56.23" resultid="15302" heatid="19322" lane="1" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.40" />
                    <SPLIT distance="100" swimtime="00:01:01.32" />
                    <SPLIT distance="150" swimtime="00:01:30.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15229" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="15269" number="2" reactiontime="+68" />
                    <RELAYPOSITION athleteid="15281" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="15291" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="398" reactiontime="+69" swimtime="00:02:12.04" resultid="15311" heatid="19564" lane="9" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                    <SPLIT distance="100" swimtime="00:01:05.55" />
                    <SPLIT distance="150" swimtime="00:01:37.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15281" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="15291" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="15235" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="15269" number="4" reactiontime="+109" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1130" points="279" reactiontime="+98" swimtime="00:02:15.43" resultid="15303" heatid="19320" lane="3" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.85" />
                    <SPLIT distance="100" swimtime="00:01:12.18" />
                    <SPLIT distance="150" swimtime="00:01:44.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15222" number="1" reactiontime="+98" />
                    <RELAYPOSITION athleteid="15214" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="15262" number="3" reactiontime="+19" />
                    <RELAYPOSITION athleteid="15235" number="4" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="282" reactiontime="+78" swimtime="00:02:28.01" resultid="15304" heatid="19562" lane="4" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.41" />
                    <SPLIT distance="100" swimtime="00:01:20.30" />
                    <SPLIT distance="150" swimtime="00:01:53.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15222" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="15242" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="15246" number="3" reactiontime="+60" />
                    <RELAYPOSITION athleteid="15262" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="WAR" clubid="18421" name="Vctory Masters Elbląg">
          <CONTACT email="lateccy@o2.pl" name="Latecki Grzegorz" street="Łokietka 45" />
          <ATHLETES>
            <ATHLETE birthdate="1954-02-04" firstname="Ewa" gender="M" lastname="Kerner-Mateusiak" nation="POL" athleteid="18436">
              <RESULTS>
                <RESULT eventid="14189" status="DNS" swimtime="00:00:00.00" resultid="18437" heatid="19615" lane="1" entrytime="00:16:00.00" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="18438" heatid="19359" lane="4" entrytime="00:05:00.00" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="18439" heatid="19434" lane="1" entrytime="00:02:20.00" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="18440" heatid="19470" lane="4" entrytime="00:02:22.00" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="18441" heatid="19486" lane="2" entrytime="00:04:40.00" />
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="18442" heatid="19531" lane="5" entrytime="00:05:00.00" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="18443" heatid="19699" lane="4" entrytime="00:08:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-05-05" firstname="Beata" gender="F" lastname="Karaś" nation="POL" athleteid="18428">
              <RESULTS>
                <RESULT eventid="1096" points="112" reactiontime="+118" swimtime="00:04:12.18" resultid="18429" heatid="19305" lane="3" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.43" />
                    <SPLIT distance="100" swimtime="00:02:01.82" />
                    <SPLIT distance="150" swimtime="00:03:19.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="155" reactiontime="+122" swimtime="00:28:29.02" resultid="18430" heatid="19624" lane="2" entrytime="00:27:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.73" />
                    <SPLIT distance="100" swimtime="00:01:45.32" />
                    <SPLIT distance="150" swimtime="00:02:40.75" />
                    <SPLIT distance="200" swimtime="00:03:37.20" />
                    <SPLIT distance="250" swimtime="00:04:34.21" />
                    <SPLIT distance="300" swimtime="00:05:31.78" />
                    <SPLIT distance="350" swimtime="00:06:29.55" />
                    <SPLIT distance="400" swimtime="00:07:27.25" />
                    <SPLIT distance="450" swimtime="00:08:24.61" />
                    <SPLIT distance="500" swimtime="00:09:22.41" />
                    <SPLIT distance="550" swimtime="00:10:20.37" />
                    <SPLIT distance="600" swimtime="00:11:17.86" />
                    <SPLIT distance="650" swimtime="00:12:15.22" />
                    <SPLIT distance="700" swimtime="00:13:12.30" />
                    <SPLIT distance="750" swimtime="00:14:10.52" />
                    <SPLIT distance="800" swimtime="00:15:08.03" />
                    <SPLIT distance="850" swimtime="00:16:06.48" />
                    <SPLIT distance="900" swimtime="00:17:03.64" />
                    <SPLIT distance="950" swimtime="00:18:00.99" />
                    <SPLIT distance="1000" swimtime="00:18:59.07" />
                    <SPLIT distance="1050" swimtime="00:19:56.71" />
                    <SPLIT distance="1100" swimtime="00:20:54.54" />
                    <SPLIT distance="1150" swimtime="00:21:51.69" />
                    <SPLIT distance="1200" swimtime="00:22:50.11" />
                    <SPLIT distance="1250" swimtime="00:23:47.32" />
                    <SPLIT distance="1300" swimtime="00:24:44.89" />
                    <SPLIT distance="1350" swimtime="00:25:14.07" />
                    <SPLIT distance="1400" swimtime="00:25:42.01" />
                    <SPLIT distance="1450" swimtime="00:27:35.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="92" reactiontime="+118" swimtime="00:04:24.42" resultid="18431" heatid="19411" lane="4" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.18" />
                    <SPLIT distance="100" swimtime="00:02:04.88" />
                    <SPLIT distance="150" swimtime="00:03:14.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="146" reactiontime="+114" swimtime="00:03:29.96" resultid="18432" heatid="19481" lane="7" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.45" />
                    <SPLIT distance="100" swimtime="00:01:40.80" />
                    <SPLIT distance="150" swimtime="00:02:35.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="111" reactiontime="+118" swimtime="00:08:59.39" resultid="18433" heatid="19503" lane="3" entrytime="00:08:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.75" />
                    <SPLIT distance="100" swimtime="00:02:05.98" />
                    <SPLIT distance="150" swimtime="00:03:19.59" />
                    <SPLIT distance="200" swimtime="00:04:29.47" />
                    <SPLIT distance="250" swimtime="00:05:48.54" />
                    <SPLIT distance="300" swimtime="00:07:08.72" />
                    <SPLIT distance="350" swimtime="00:08:05.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="87" reactiontime="+118" swimtime="00:02:02.84" resultid="18434" heatid="19513" lane="2" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="147" reactiontime="+113" swimtime="00:07:24.08" resultid="18435" heatid="19696" lane="8" entrytime="00:07:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.95" />
                    <SPLIT distance="100" swimtime="00:01:45.77" />
                    <SPLIT distance="150" swimtime="00:02:43.18" />
                    <SPLIT distance="200" swimtime="00:03:40.11" />
                    <SPLIT distance="250" swimtime="00:04:37.06" />
                    <SPLIT distance="300" swimtime="00:05:34.10" />
                    <SPLIT distance="350" swimtime="00:06:30.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-08-31" firstname="Karolina" gender="F" lastname="Karaś" nation="POL" athleteid="18422">
              <RESULTS>
                <RESULT eventid="1062" points="136" reactiontime="+109" swimtime="00:00:45.14" resultid="18423" heatid="19277" lane="0" entrytime="00:00:45.00" />
                <RESULT eventid="1147" reactiontime="+95" status="OTL" swimtime="00:14:48.63" resultid="18424" heatid="19596" lane="9" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.04" />
                    <SPLIT distance="100" swimtime="00:01:43.10" />
                    <SPLIT distance="150" swimtime="00:02:38.61" />
                    <SPLIT distance="200" swimtime="00:03:34.20" />
                    <SPLIT distance="250" swimtime="00:04:31.22" />
                    <SPLIT distance="300" swimtime="00:05:27.68" />
                    <SPLIT distance="350" swimtime="00:06:24.00" />
                    <SPLIT distance="400" swimtime="00:07:19.86" />
                    <SPLIT distance="450" swimtime="00:08:15.53" />
                    <SPLIT distance="500" swimtime="00:09:11.21" />
                    <SPLIT distance="550" swimtime="00:10:08.91" />
                    <SPLIT distance="600" swimtime="00:11:05.66" />
                    <SPLIT distance="650" swimtime="00:12:01.71" />
                    <SPLIT distance="700" swimtime="00:12:58.14" />
                    <SPLIT distance="750" swimtime="00:13:55.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="146" reactiontime="+101" swimtime="00:01:36.57" resultid="18425" heatid="19368" lane="2" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="154" reactiontime="+104" swimtime="00:03:26.61" resultid="18426" heatid="19481" lane="0" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.91" />
                    <SPLIT distance="100" swimtime="00:01:39.73" />
                    <SPLIT distance="150" swimtime="00:02:33.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="158" reactiontime="+109" swimtime="00:07:13.40" resultid="18427" heatid="19695" lane="4" entrytime="00:07:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.50" />
                    <SPLIT distance="100" swimtime="00:01:41.74" />
                    <SPLIT distance="150" swimtime="00:02:37.48" />
                    <SPLIT distance="200" swimtime="00:03:33.68" />
                    <SPLIT distance="250" swimtime="00:04:30.10" />
                    <SPLIT distance="300" swimtime="00:05:26.41" />
                    <SPLIT distance="350" swimtime="00:06:22.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-02-04" firstname="Ewa" gender="F" lastname="Kerner-Mateusiak" nation="POL" athleteid="19741">
              <RESULTS>
                <RESULT eventid="1147" reactiontime="+138" status="DNF" swimtime="00:00:00.00" resultid="19742" heatid="19594" lane="9" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.53" />
                    <SPLIT distance="100" swimtime="00:02:22.75" />
                    <SPLIT distance="150" swimtime="00:03:41.66" />
                    <SPLIT distance="200" swimtime="00:05:01.05" />
                    <SPLIT distance="250" swimtime="00:06:20.45" />
                    <SPLIT distance="300" swimtime="00:07:43.25" />
                    <SPLIT distance="350" swimtime="00:09:09.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="58" reactiontime="+116" swimtime="00:05:47.18" resultid="19743" heatid="19354" lane="6" late="yes" />
                <RESULT comment="K14 - Praca nóg w płaszczyźnie pionowej w dół (z wyjątkiem jednego ruchu po starcie i nawrocie) (Time: 16:11)" eventid="1388" reactiontime="+119" status="DSQ" swimtime="00:02:48.52" resultid="19744" heatid="19426" lane="7" late="yes" />
                <RESULT eventid="1457" points="47" reactiontime="+115" swimtime="00:02:31.94" resultid="19745" heatid="19465" lane="8" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="56" reactiontime="+118" swimtime="00:10:12.92" resultid="19747" heatid="19694" lane="6" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.79" />
                    <SPLIT distance="100" swimtime="00:02:22.07" />
                    <SPLIT distance="150" swimtime="00:03:41.02" />
                    <SPLIT distance="200" swimtime="00:05:02.10" />
                    <SPLIT distance="250" swimtime="00:06:21.33" />
                    <SPLIT distance="300" swimtime="00:07:40.08" />
                    <SPLIT distance="350" swimtime="00:08:58.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="VSKUK" nation="SVK" region="BAO" clubid="18552" name="Vysokoskolsky klub Univerzity komenskeho" shortname="Vysokoskolsky klub Univerzity " shortname.en="Vskuk">
          <ATHLETES>
            <ATHLETE birthdate="1973-11-11" firstname="Martin" gender="M" lastname="Hlavatý" nation="SVK" license="SVK11444" athleteid="18553">
              <RESULTS>
                <RESULT eventid="1113" points="464" reactiontime="+74" swimtime="00:02:21.60" resultid="18554" heatid="19317" lane="5" entrytime="00:02:23.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.83" />
                    <SPLIT distance="100" swimtime="00:01:08.08" />
                    <SPLIT distance="150" swimtime="00:01:48.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="441" reactiontime="+77" swimtime="00:02:38.23" resultid="18555" heatid="19365" lane="0" entrytime="00:02:38.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                    <SPLIT distance="100" swimtime="00:01:15.66" />
                    <SPLIT distance="150" swimtime="00:01:57.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="523" reactiontime="+68" swimtime="00:01:02.40" resultid="18556" heatid="19409" lane="7" entrytime="00:01:03.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="572" reactiontime="+76" swimtime="00:01:06.99" resultid="18557" heatid="19443" lane="1" entrytime="00:01:06.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="510" reactiontime="+69" swimtime="00:00:27.28" resultid="18558" heatid="19462" lane="7" entrytime="00:00:27.50" entrycourse="SCM" />
                <RESULT eventid="1681" points="607" reactiontime="+70" swimtime="00:00:29.81" resultid="18559" heatid="19560" lane="3" entrytime="00:00:29.60" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-11-07" firstname="Marian" gender="M" lastname="Horínek" nation="SVK" license="SVK11041" athleteid="18560">
              <RESULTS>
                <RESULT eventid="1113" points="452" reactiontime="+83" swimtime="00:02:22.78" resultid="18561" heatid="19317" lane="3" entrytime="00:02:23.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.53" />
                    <SPLIT distance="100" swimtime="00:01:08.52" />
                    <SPLIT distance="150" swimtime="00:01:50.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="511" reactiontime="+78" swimtime="00:00:56.20" resultid="18562" heatid="19387" lane="6" entrytime="00:00:56.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="507" reactiontime="+79" swimtime="00:02:04.57" resultid="18563" heatid="19496" lane="7" entrytime="00:02:03.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                    <SPLIT distance="100" swimtime="00:01:00.91" />
                    <SPLIT distance="150" swimtime="00:01:32.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="489" reactiontime="+85" swimtime="00:04:29.26" resultid="18564" heatid="19708" lane="3" entrytime="00:04:25.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.25" />
                    <SPLIT distance="100" swimtime="00:01:05.35" />
                    <SPLIT distance="150" swimtime="00:01:39.92" />
                    <SPLIT distance="200" swimtime="00:02:14.49" />
                    <SPLIT distance="250" swimtime="00:02:48.56" />
                    <SPLIT distance="300" swimtime="00:03:22.45" />
                    <SPLIT distance="350" swimtime="00:03:56.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WMT" nation="POL" region="MAZ" clubid="17300" name="Warsaw Masters Team">
          <CONTACT email="agnieszka.z.mazurkiewicz@gmail.com" name="Agnieszka Mazurkiewicz" phone="882 185 766" state="MAZ" zip="WAW" />
          <ATHLETES>
            <ATHLETE birthdate="1975-01-05" firstname="Bartłomiej" gender="M" lastname="Pawłowski" nation="POL" athleteid="17402">
              <RESULTS>
                <RESULT eventid="1079" points="342" reactiontime="+78" swimtime="00:00:28.95" resultid="17403" heatid="19293" lane="9" entrytime="00:00:30.00" />
                <RESULT eventid="1239" points="289" reactiontime="+93" swimtime="00:03:01.97" resultid="17404" heatid="19362" lane="2" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.63" />
                    <SPLIT distance="100" swimtime="00:01:26.67" />
                    <SPLIT distance="150" swimtime="00:02:14.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" status="DNS" swimtime="00:00:00.00" resultid="17405" heatid="19403" lane="7" entrytime="00:01:17.00" />
                <RESULT eventid="1406" points="350" reactiontime="+81" swimtime="00:01:18.86" resultid="17406" heatid="19438" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="379" reactiontime="+75" swimtime="00:00:34.89" resultid="17407" heatid="19555" lane="7" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-10-04" firstname="Maciej" gender="M" lastname="Szymański" nation="POL" athleteid="17472">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="17473" heatid="19303" lane="2" entrytime="00:00:24.85" />
                <RESULT eventid="1205" points="439" reactiontime="+73" swimtime="00:00:29.22" resultid="17474" heatid="19352" lane="5" entrytime="00:00:28.50" />
                <RESULT eventid="14243" points="537" reactiontime="+76" swimtime="00:01:01.85" resultid="17475" heatid="19409" lane="5" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="519" reactiontime="+73" swimtime="00:00:27.11" resultid="17476" heatid="19450" lane="6" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="17477" heatid="19478" lane="6" entrytime="00:01:02.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-09-13" firstname="Michał" gender="M" lastname="Jabłoński" nation="POL" athleteid="17455">
              <RESULTS>
                <RESULT eventid="1273" points="326" reactiontime="+76" swimtime="00:01:05.26" resultid="17456" heatid="19381" lane="4" entrytime="00:01:05.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="251" reactiontime="+87" swimtime="00:02:52.07" resultid="17457" heatid="19416" lane="1" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.51" />
                    <SPLIT distance="100" swimtime="00:01:23.12" />
                    <SPLIT distance="150" swimtime="00:02:08.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="17458" heatid="19457" lane="5" entrytime="00:00:31.40" />
                <RESULT eventid="1613" points="293" reactiontime="+81" swimtime="00:01:12.37" resultid="17459" heatid="19521" lane="6" entrytime="00:01:12.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-06-10" firstname="Łukasz" gender="M" lastname="Rybiński" nation="POL" athleteid="17500">
              <RESULTS>
                <RESULT eventid="1239" points="233" reactiontime="+95" swimtime="00:03:15.60" resultid="17501" heatid="19362" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.93" />
                    <SPLIT distance="100" swimtime="00:01:30.67" />
                    <SPLIT distance="150" swimtime="00:02:21.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="273" reactiontime="+97" swimtime="00:01:09.25" resultid="17502" heatid="19380" lane="5" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="17503" heatid="19437" lane="4" entrytime="00:01:28.00" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="17504" heatid="19490" lane="9" entrytime="00:02:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-07-26" firstname="Anna" gender="F" lastname="Szemberg" nation="POL" athleteid="17434">
              <RESULTS>
                <RESULT eventid="1147" points="108" reactiontime="+104" swimtime="00:16:44.23" resultid="17435" heatid="19594" lane="4" entrytime="00:16:21.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.46" />
                    <SPLIT distance="100" swimtime="00:02:01.61" />
                    <SPLIT distance="150" swimtime="00:03:04.61" />
                    <SPLIT distance="200" swimtime="00:04:08.52" />
                    <SPLIT distance="250" swimtime="00:05:14.63" />
                    <SPLIT distance="300" swimtime="00:06:19.24" />
                    <SPLIT distance="350" swimtime="00:07:21.64" />
                    <SPLIT distance="400" swimtime="00:08:24.31" />
                    <SPLIT distance="450" swimtime="00:09:28.12" />
                    <SPLIT distance="500" swimtime="00:10:30.39" />
                    <SPLIT distance="550" swimtime="00:11:33.39" />
                    <SPLIT distance="600" swimtime="00:12:37.34" />
                    <SPLIT distance="650" swimtime="00:13:39.90" />
                    <SPLIT distance="700" swimtime="00:14:42.92" />
                    <SPLIT distance="750" swimtime="00:15:44.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="87" reactiontime="+95" swimtime="00:01:54.88" resultid="17436" heatid="19367" lane="4" entrytime="00:01:54.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" status="DNS" swimtime="00:00:00.00" resultid="17437" heatid="19389" lane="5" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="17438" heatid="19480" lane="8" entrytime="00:04:01.55" />
                <RESULT eventid="1721" points="103" reactiontime="+101" swimtime="00:08:19.93" resultid="17439" heatid="19695" lane="2" entrytime="00:08:18.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.89" />
                    <SPLIT distance="100" swimtime="00:02:00.59" />
                    <SPLIT distance="150" swimtime="00:03:06.35" />
                    <SPLIT distance="200" swimtime="00:06:17.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-06-07" firstname="Olga" gender="F" lastname="Krysiak" nation="POL" athleteid="17376">
              <RESULTS>
                <RESULT eventid="1062" points="519" reactiontime="+77" swimtime="00:00:28.91" resultid="17377" heatid="19283" lane="1" entrytime="00:00:28.21" />
                <RESULT eventid="1256" points="536" reactiontime="+72" swimtime="00:01:02.64" resultid="17378" heatid="19372" lane="8" entrytime="00:01:02.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" status="DNS" swimtime="00:00:00.00" resultid="17379" heatid="19448" lane="7" entrytime="00:00:33.40" />
                <RESULT eventid="1491" points="491" reactiontime="+79" swimtime="00:02:20.39" resultid="17380" heatid="19484" lane="2" entrytime="00:02:21.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                    <SPLIT distance="100" swimtime="00:01:06.44" />
                    <SPLIT distance="150" swimtime="00:01:43.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="378" reactiontime="+75" swimtime="00:05:24.30" resultid="17381" heatid="19698" lane="7" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                    <SPLIT distance="100" swimtime="00:01:15.72" />
                    <SPLIT distance="150" swimtime="00:01:57.64" />
                    <SPLIT distance="200" swimtime="00:02:39.87" />
                    <SPLIT distance="250" swimtime="00:03:22.51" />
                    <SPLIT distance="300" swimtime="00:04:04.05" />
                    <SPLIT distance="350" swimtime="00:04:45.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-06-10" firstname="Tomasz" gender="M" lastname="Porada" nation="POL" athleteid="17301">
              <RESULTS>
                <RESULT eventid="1079" points="401" reactiontime="+69" swimtime="00:00:27.46" resultid="17302" heatid="19299" lane="9" entrytime="00:00:27.50" />
                <RESULT eventid="1113" points="399" reactiontime="+81" swimtime="00:02:28.81" resultid="17303" heatid="19316" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.49" />
                    <SPLIT distance="100" swimtime="00:01:12.26" />
                    <SPLIT distance="150" swimtime="00:01:53.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="475" reactiontime="+76" swimtime="00:02:34.27" resultid="17304" heatid="19364" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.03" />
                    <SPLIT distance="100" swimtime="00:01:14.19" />
                    <SPLIT distance="150" swimtime="00:01:53.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="454" reactiontime="+75" swimtime="00:01:12.31" resultid="17305" heatid="19441" lane="6" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="465" reactiontime="+82" swimtime="00:00:32.57" resultid="17306" heatid="19557" lane="1" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-24" firstname="Jan" gender="M" lastname="Pfitzner" nation="POL" athleteid="17440">
              <RESULTS>
                <RESULT eventid="1205" points="351" reactiontime="+73" swimtime="00:00:31.48" resultid="17441" heatid="19352" lane="8" entrytime="00:00:29.50" />
                <RESULT eventid="1440" points="396" reactiontime="+86" swimtime="00:00:29.67" resultid="17442" heatid="19462" lane="2" entrytime="00:00:27.50" />
                <RESULT eventid="1681" points="363" reactiontime="+75" swimtime="00:00:35.38" resultid="17443" heatid="19555" lane="5" entrytime="00:00:35.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-28" firstname="Karol" gender="M" lastname="Dzięcioł" nation="POL" athleteid="17491">
              <RESULTS>
                <RESULT eventid="1079" points="476" reactiontime="+66" swimtime="00:00:25.93" resultid="17492" heatid="19302" lane="0" entrytime="00:00:25.90" />
                <RESULT eventid="1273" points="497" reactiontime="+77" swimtime="00:00:56.72" resultid="17493" heatid="19386" lane="6" entrytime="00:00:57.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="448" reactiontime="+84" swimtime="00:01:05.73" resultid="17494" heatid="19408" lane="2" entrytime="00:01:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="353" reactiontime="+86" swimtime="00:05:00.19" resultid="17495" heatid="19706" lane="4" entrytime="00:04:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.31" />
                    <SPLIT distance="100" swimtime="00:01:07.80" />
                    <SPLIT distance="150" swimtime="00:01:45.14" />
                    <SPLIT distance="200" swimtime="00:02:23.47" />
                    <SPLIT distance="250" swimtime="00:03:02.21" />
                    <SPLIT distance="300" swimtime="00:03:41.96" />
                    <SPLIT distance="350" swimtime="00:04:21.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-10-03" firstname="Ryszard" gender="M" lastname="Sielski" nation="POL" athleteid="17344">
              <RESULTS>
                <RESULT eventid="1205" points="27" reactiontime="+82" swimtime="00:01:13.20" resultid="17345" heatid="19342" lane="5" entrytime="00:01:15.00" />
                <RESULT eventid="14243" points="38" reactiontime="+138" swimtime="00:02:28.86" resultid="17346" heatid="19397" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="57" reactiontime="+133" swimtime="00:02:23.87" resultid="17347" heatid="19435" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="25" reactiontime="+130" swimtime="00:01:14.20" resultid="17348" heatid="19450" lane="5" entrytime="00:01:35.00" />
                <RESULT eventid="1647" points="27" reactiontime="+85" swimtime="00:05:50.99" resultid="17349" heatid="19531" lane="7" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.96" />
                    <SPLIT distance="100" swimtime="00:02:56.68" />
                    <SPLIT distance="150" swimtime="00:04:29.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="75" reactiontime="+127" swimtime="00:00:59.87" resultid="17350" heatid="19547" lane="7" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-07-13" firstname="Sebastian" gender="M" lastname="Ostapczuk" nation="POL" athleteid="17364">
              <RESULTS>
                <RESULT eventid="1239" points="189" swimtime="00:03:29.75" resultid="17365" heatid="19361" lane="9" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.92" />
                    <SPLIT distance="100" swimtime="00:01:41.00" />
                    <SPLIT distance="150" swimtime="00:02:36.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="175" reactiontime="+109" swimtime="00:01:20.34" resultid="17366" heatid="19375" lane="8" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="191" reactiontime="+105" swimtime="00:01:36.50" resultid="17367" heatid="19435" lane="7" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-12-11" firstname="Igor" gender="M" lastname="Rębas" nation="POL" athleteid="17484">
              <RESULTS>
                <RESULT eventid="1079" points="446" reactiontime="+73" swimtime="00:00:26.50" resultid="17485" heatid="19300" lane="4" entrytime="00:00:26.00" />
                <RESULT eventid="1273" points="556" reactiontime="+78" swimtime="00:00:54.63" resultid="17486" heatid="19385" lane="0" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="491" reactiontime="+74" swimtime="00:01:03.75" resultid="17487" heatid="19409" lane="3" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="543" reactiontime="+78" swimtime="00:00:26.72" resultid="17488" heatid="19464" lane="0" entrytime="00:00:26.00" />
                <RESULT eventid="1508" points="503" reactiontime="+74" swimtime="00:02:04.89" resultid="17489" heatid="19495" lane="9" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.93" />
                    <SPLIT distance="100" swimtime="00:01:01.03" />
                    <SPLIT distance="150" swimtime="00:01:34.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="17490" heatid="19525" lane="6" entrytime="00:00:58.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-06-16" firstname="Paweł" gender="M" lastname="Witkowski" nation="POL" athleteid="17415">
              <RESULTS>
                <RESULT eventid="1406" points="482" reactiontime="+86" swimtime="00:01:10.88" resultid="17416" heatid="19440" lane="5" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="497" reactiontime="+87" swimtime="00:00:31.87" resultid="17417" heatid="19557" lane="6" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-10" firstname="Michał" gender="M" lastname="Rudziński" nation="POL" athleteid="17390">
              <RESULTS>
                <RESULT eventid="1239" points="218" reactiontime="+108" swimtime="00:03:20.09" resultid="17391" heatid="19361" lane="4" entrytime="00:03:18.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.71" />
                    <SPLIT distance="100" swimtime="00:01:34.24" />
                    <SPLIT distance="150" swimtime="00:02:25.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="126" reactiontime="+106" swimtime="00:03:36.13" resultid="17392" heatid="19414" lane="4" entrytime="00:03:52.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.24" />
                    <SPLIT distance="100" swimtime="00:01:39.88" />
                    <SPLIT distance="150" swimtime="00:02:36.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="206" reactiontime="+108" swimtime="00:01:34.06" resultid="17393" heatid="19436" lane="5" entrytime="00:01:31.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="131" reactiontime="+112" swimtime="00:01:34.52" resultid="17394" heatid="19518" lane="3" entrytime="00:01:37.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="215" reactiontime="+105" swimtime="00:00:42.13" resultid="17395" heatid="19551" lane="8" entrytime="00:00:41.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-20" firstname="Robert" gender="M" lastname="Budek" nation="POL" athleteid="17396">
              <RESULTS>
                <RESULT eventid="1079" points="246" reactiontime="+82" swimtime="00:00:32.33" resultid="17397" heatid="19290" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1273" points="193" reactiontime="+79" swimtime="00:01:17.68" resultid="17398" heatid="19378" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" status="DNS" swimtime="00:00:00.00" resultid="17399" heatid="19400" lane="2" entrytime="00:01:30.00" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="17400" heatid="19451" lane="2" entrytime="00:00:50.00" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="17401" heatid="19549" lane="4" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-08-12" firstname="Jakub" gender="M" lastname="Szulc" nation="POL" athleteid="17465">
              <RESULTS>
                <RESULT eventid="1079" points="383" reactiontime="+83" swimtime="00:00:27.89" resultid="17466" heatid="19298" lane="3" entrytime="00:00:27.50" />
                <RESULT eventid="1205" points="293" reactiontime="+88" swimtime="00:00:33.43" resultid="17467" heatid="19348" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="14243" points="346" reactiontime="+77" swimtime="00:01:11.62" resultid="17468" heatid="19405" lane="5" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="379" reactiontime="+83" swimtime="00:00:30.11" resultid="17469" heatid="19458" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="1508" points="403" reactiontime="+81" swimtime="00:02:14.43" resultid="17470" heatid="19493" lane="3" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.70" />
                    <SPLIT distance="100" swimtime="00:01:06.11" />
                    <SPLIT distance="150" swimtime="00:01:40.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="369" reactiontime="+78" swimtime="00:04:55.72" resultid="17471" heatid="19706" lane="8" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.14" />
                    <SPLIT distance="100" swimtime="00:01:08.96" />
                    <SPLIT distance="150" swimtime="00:01:45.61" />
                    <SPLIT distance="200" swimtime="00:02:22.74" />
                    <SPLIT distance="250" swimtime="00:03:00.51" />
                    <SPLIT distance="300" swimtime="00:03:39.20" />
                    <SPLIT distance="350" swimtime="00:04:17.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-02-23" firstname="Joanna" gender="F" lastname="Gołębiowska" nation="POL" athleteid="17444">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="14225" points="598" reactiontime="+74" swimtime="00:01:07.25" resultid="17445" heatid="19396" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="550" reactiontime="+75" swimtime="00:00:29.74" resultid="17446" heatid="19449" lane="4" entrytime="00:00:29.50" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1595" points="568" reactiontime="+79" swimtime="00:01:05.92" resultid="17447" heatid="19515" lane="4" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-10-06" firstname="Mateusz" gender="M" lastname="Bednarz" nation="POL" athleteid="17351">
              <RESULTS>
                <RESULT eventid="1079" points="356" reactiontime="+79" swimtime="00:00:28.57" resultid="17352" heatid="19296" lane="7" entrytime="00:00:28.76" />
                <RESULT comment="K15 - Brak dotknięcia ściany obydwoma rozłączonymi dłońmi przy nawrocie lub na zakończenie wyścigu (Time: 16:34), Z-2" eventid="1113" reactiontime="+107" status="DSQ" swimtime="00:02:35.98" resultid="17353" heatid="19314" lane="2" entrytime="00:02:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                    <SPLIT distance="100" swimtime="00:01:13.70" />
                    <SPLIT distance="150" swimtime="00:02:00.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="258" reactiontime="+76" swimtime="00:00:34.88" resultid="17354" heatid="19347" lane="7" entrytime="00:00:37.27" />
                <RESULT eventid="14243" points="349" reactiontime="+82" swimtime="00:01:11.38" resultid="17355" heatid="19404" lane="5" entrytime="00:01:13.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="364" reactiontime="+89" swimtime="00:00:30.53" resultid="17356" heatid="19456" lane="5" entrytime="00:00:32.01" />
                <RESULT eventid="1508" points="369" reactiontime="+73" swimtime="00:02:18.50" resultid="17357" heatid="19493" lane="0" entrytime="00:02:20.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                    <SPLIT distance="100" swimtime="00:01:07.87" />
                    <SPLIT distance="150" swimtime="00:01:44.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="328" reactiontime="+87" swimtime="00:01:09.67" resultid="17358" heatid="19521" lane="9" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="373" reactiontime="+97" swimtime="00:04:54.85" resultid="17359" heatid="19706" lane="1" entrytime="00:05:01.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                    <SPLIT distance="100" swimtime="00:01:09.20" />
                    <SPLIT distance="150" swimtime="00:02:24.25" />
                    <SPLIT distance="250" swimtime="00:03:02.73" />
                    <SPLIT distance="300" swimtime="00:03:41.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-12-06" firstname="Mateusz" gender="M" lastname="Grula" nation="POL" athleteid="17430">
              <RESULTS>
                <RESULT eventid="14243" points="635" reactiontime="+72" swimtime="00:00:58.51" resultid="17431" heatid="19410" lane="0" entrytime="00:01:00.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="638" reactiontime="+65" swimtime="00:01:04.57" resultid="17432" heatid="19443" lane="9" entrytime="00:01:07.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="617" reactiontime="+65" swimtime="00:00:29.65" resultid="17433" heatid="19560" lane="6" entrytime="00:00:29.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-13" firstname="Agnieszka" gender="F" lastname="Mazurkiewicz" nation="POL" athleteid="17496">
              <RESULTS>
                <RESULT eventid="1256" points="267" reactiontime="+92" swimtime="00:01:19.03" resultid="17497" heatid="19369" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="262" reactiontime="+96" swimtime="00:02:52.91" resultid="17498" heatid="19482" lane="3" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.61" />
                    <SPLIT distance="100" swimtime="00:01:22.54" />
                    <SPLIT distance="150" swimtime="00:02:07.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="236" reactiontime="+95" swimtime="00:06:19.14" resultid="17499" heatid="19697" lane="1" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.14" />
                    <SPLIT distance="100" swimtime="00:01:27.79" />
                    <SPLIT distance="150" swimtime="00:02:16.51" />
                    <SPLIT distance="200" swimtime="00:03:04.77" />
                    <SPLIT distance="250" swimtime="00:03:53.21" />
                    <SPLIT distance="300" swimtime="00:04:42.40" />
                    <SPLIT distance="350" swimtime="00:05:32.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-08-01" firstname="Edyta" gender="F" lastname="Olszewska" nation="POL" athleteid="17418">
              <RESULTS>
                <RESULT eventid="1222" points="356" reactiontime="+87" swimtime="00:03:09.87" resultid="17419" heatid="19358" lane="1" entrytime="00:03:09.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.93" />
                    <SPLIT distance="100" swimtime="00:01:32.63" />
                    <SPLIT distance="150" swimtime="00:02:20.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="340" reactiontime="+79" swimtime="00:01:29.31" resultid="17420" heatid="19431" lane="6" entrytime="00:01:27.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="268" reactiontime="+78" swimtime="00:02:51.63" resultid="17421" heatid="19483" lane="8" entrytime="00:02:47.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                    <SPLIT distance="100" swimtime="00:01:23.40" />
                    <SPLIT distance="150" swimtime="00:02:06.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="354" reactiontime="+81" swimtime="00:00:40.45" resultid="17422" heatid="19543" lane="0" entrytime="00:00:40.53" />
                <RESULT eventid="1721" points="277" reactiontime="+83" swimtime="00:05:59.43" resultid="17423" heatid="19697" lane="6" entrytime="00:05:56.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.60" />
                    <SPLIT distance="100" swimtime="00:01:24.79" />
                    <SPLIT distance="150" swimtime="00:02:10.48" />
                    <SPLIT distance="200" swimtime="00:02:56.05" />
                    <SPLIT distance="250" swimtime="00:03:40.99" />
                    <SPLIT distance="300" swimtime="00:04:26.12" />
                    <SPLIT distance="350" swimtime="00:05:12.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-05-31" firstname="Katharina" gender="F" lastname="Szymańska" nation="POL" athleteid="17478">
              <RESULTS>
                <RESULT eventid="1096" points="166" reactiontime="+96" swimtime="00:03:41.40" resultid="17479" heatid="19305" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.63" />
                    <SPLIT distance="100" swimtime="00:01:49.20" />
                    <SPLIT distance="150" swimtime="00:02:48.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="177" reactiontime="+94" swimtime="00:01:40.88" resultid="17480" heatid="19389" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="108" reactiontime="+96" swimtime="00:04:10.85" resultid="17481" heatid="19411" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.25" />
                    <SPLIT distance="100" swimtime="00:01:54.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" status="DNS" swimtime="00:00:00.00" resultid="17482" heatid="19444" lane="4" />
                <RESULT eventid="1595" status="DNS" swimtime="00:00:00.00" resultid="17483" heatid="19513" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-03" firstname="Robert" gender="M" lastname="Sutowski" nation="POL" athleteid="17307">
              <RESULTS>
                <RESULT eventid="1079" points="136" reactiontime="+104" swimtime="00:00:39.38" resultid="17308" heatid="19286" lane="6" entrytime="00:00:39.10" />
                <RESULT eventid="14189" points="162" reactiontime="+107" swimtime="00:13:33.41" resultid="17309" heatid="19615" lane="5" entrytime="00:14:05.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.30" />
                    <SPLIT distance="100" swimtime="00:01:35.93" />
                    <SPLIT distance="150" swimtime="00:02:28.03" />
                    <SPLIT distance="200" swimtime="00:03:19.59" />
                    <SPLIT distance="250" swimtime="00:04:11.18" />
                    <SPLIT distance="300" swimtime="00:05:03.19" />
                    <SPLIT distance="350" swimtime="00:05:54.94" />
                    <SPLIT distance="400" swimtime="00:06:47.25" />
                    <SPLIT distance="450" swimtime="00:07:38.72" />
                    <SPLIT distance="500" swimtime="00:08:30.23" />
                    <SPLIT distance="550" swimtime="00:09:21.08" />
                    <SPLIT distance="600" swimtime="00:10:13.55" />
                    <SPLIT distance="650" swimtime="00:11:05.78" />
                    <SPLIT distance="700" swimtime="00:11:57.30" />
                    <SPLIT distance="750" swimtime="00:12:46.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="57" reactiontime="+136" swimtime="00:00:57.43" resultid="17310" heatid="19344" lane="9" entrytime="00:00:55.01" />
                <RESULT eventid="1273" points="143" reactiontime="+110" swimtime="00:01:25.90" resultid="17311" heatid="19376" lane="2" entrytime="00:01:25.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="101" reactiontime="+108" swimtime="00:00:46.68" resultid="17312" heatid="19451" lane="3" entrytime="00:00:46.76" />
                <RESULT eventid="1508" points="154" reactiontime="+109" swimtime="00:03:05.08" resultid="17313" heatid="19488" lane="0" entrytime="00:03:09.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.94" />
                    <SPLIT distance="100" swimtime="00:01:31.22" />
                    <SPLIT distance="150" swimtime="00:02:19.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="77" reactiontime="+109" swimtime="00:01:52.96" resultid="17314" heatid="19518" lane="9" entrytime="00:01:53.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="17315" heatid="19701" lane="7" entrytime="00:06:38.19" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-05-04" firstname="Ewa" gender="F" lastname="Matlak" nation="POL" athleteid="17382">
              <RESULTS>
                <RESULT eventid="1423" points="282" reactiontime="+90" swimtime="00:00:37.14" resultid="17383" heatid="19447" lane="3" entrytime="00:00:36.00" />
                <RESULT eventid="1491" points="302" reactiontime="+84" swimtime="00:02:45.04" resultid="17384" heatid="19483" lane="2" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                    <SPLIT distance="100" swimtime="00:01:18.09" />
                    <SPLIT distance="150" swimtime="00:02:01.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="257" reactiontime="+83" swimtime="00:01:25.81" resultid="17385" heatid="19514" lane="7" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="310" reactiontime="+88" swimtime="00:05:46.19" resultid="17386" heatid="19697" lane="5" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.16" />
                    <SPLIT distance="100" swimtime="00:01:20.84" />
                    <SPLIT distance="150" swimtime="00:02:04.57" />
                    <SPLIT distance="200" swimtime="00:02:48.55" />
                    <SPLIT distance="250" swimtime="00:03:33.30" />
                    <SPLIT distance="300" swimtime="00:04:17.83" />
                    <SPLIT distance="350" swimtime="00:05:02.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-22" firstname="Timea" gender="F" lastname="Balajcza" nation="POL" athleteid="17327">
              <RESULTS>
                <RESULT eventid="1096" points="258" reactiontime="+92" swimtime="00:03:11.24" resultid="17328" heatid="19306" lane="2" entrytime="00:03:20.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.63" />
                    <SPLIT distance="100" swimtime="00:01:32.93" />
                    <SPLIT distance="150" swimtime="00:02:23.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="253" reactiontime="+98" swimtime="00:12:37.31" resultid="17329" heatid="19595" lane="2" entrytime="00:13:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.04" />
                    <SPLIT distance="100" swimtime="00:01:27.72" />
                    <SPLIT distance="150" swimtime="00:02:14.85" />
                    <SPLIT distance="200" swimtime="00:03:02.94" />
                    <SPLIT distance="250" swimtime="00:03:51.01" />
                    <SPLIT distance="300" swimtime="00:04:38.87" />
                    <SPLIT distance="350" swimtime="00:05:27.19" />
                    <SPLIT distance="400" swimtime="00:06:15.47" />
                    <SPLIT distance="450" swimtime="00:07:03.38" />
                    <SPLIT distance="500" swimtime="00:07:50.60" />
                    <SPLIT distance="550" swimtime="00:08:38.45" />
                    <SPLIT distance="600" swimtime="00:09:26.72" />
                    <SPLIT distance="650" swimtime="00:10:14.96" />
                    <SPLIT distance="700" swimtime="00:11:03.46" />
                    <SPLIT distance="750" swimtime="00:11:51.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="301" reactiontime="+95" swimtime="00:03:20.62" resultid="17330" heatid="19357" lane="3" entrytime="00:03:20.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.85" />
                    <SPLIT distance="100" swimtime="00:01:36.44" />
                    <SPLIT distance="150" swimtime="00:02:28.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="256" reactiontime="+95" swimtime="00:01:29.21" resultid="17331" heatid="19392" lane="2" entrytime="00:01:28.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="297" reactiontime="+89" swimtime="00:01:33.41" resultid="17332" heatid="19430" lane="6" entrytime="00:01:33.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="233" reactiontime="+99" swimtime="00:02:59.85" resultid="17333" heatid="19481" lane="4" entrytime="00:03:02.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.16" />
                    <SPLIT distance="100" swimtime="00:01:26.90" />
                    <SPLIT distance="150" swimtime="00:02:13.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="303" reactiontime="+89" swimtime="00:00:42.64" resultid="17334" heatid="19542" lane="4" entrytime="00:00:41.81" />
                <RESULT eventid="1721" points="245" reactiontime="+92" swimtime="00:06:14.70" resultid="17335" heatid="19696" lane="4" entrytime="00:06:18.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.61" />
                    <SPLIT distance="100" swimtime="00:01:29.01" />
                    <SPLIT distance="150" swimtime="00:02:17.40" />
                    <SPLIT distance="200" swimtime="00:03:05.75" />
                    <SPLIT distance="250" swimtime="00:03:52.92" />
                    <SPLIT distance="300" swimtime="00:04:39.59" />
                    <SPLIT distance="350" swimtime="00:05:27.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-05-25" firstname="Patryk" gender="M" lastname="Gąsior" nation="POL" athleteid="17322">
              <RESULTS>
                <RESULT eventid="1113" points="633" reactiontime="+78" swimtime="00:02:07.68" resultid="17323" heatid="19318" lane="3" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.60" />
                    <SPLIT distance="100" swimtime="00:01:00.83" />
                    <SPLIT distance="150" swimtime="00:01:37.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="630" reactiontime="+82" swimtime="00:02:06.60" resultid="17324" heatid="19418" lane="4" entrytime="00:02:05.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.31" />
                    <SPLIT distance="100" swimtime="00:01:00.92" />
                    <SPLIT distance="150" swimtime="00:01:33.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="616" reactiontime="+79" swimtime="00:04:36.72" resultid="17325" heatid="19512" lane="4" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.47" />
                    <SPLIT distance="100" swimtime="00:01:04.22" />
                    <SPLIT distance="150" swimtime="00:01:38.39" />
                    <SPLIT distance="200" swimtime="00:02:12.48" />
                    <SPLIT distance="250" swimtime="00:02:51.67" />
                    <SPLIT distance="300" swimtime="00:03:31.19" />
                    <SPLIT distance="350" swimtime="00:04:05.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="522" reactiontime="+76" swimtime="00:02:11.14" resultid="17326" heatid="19537" lane="4" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.86" />
                    <SPLIT distance="100" swimtime="00:01:03.11" />
                    <SPLIT distance="150" swimtime="00:01:37.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-20" firstname="Katarzyna" gender="F" lastname="Dziedzic" nation="POL" athleteid="17360">
              <RESULTS>
                <RESULT eventid="14225" points="326" reactiontime="+84" swimtime="00:01:22.30" resultid="17361" heatid="19389" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" status="DNS" swimtime="00:00:00.00" resultid="17362" heatid="19430" lane="9" entrytime="00:01:37.00" />
                <RESULT eventid="1423" points="327" reactiontime="+71" swimtime="00:00:35.36" resultid="17363" heatid="19448" lane="9" entrytime="00:00:35.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-06-17" firstname="Leszek" gender="M" lastname="Madej" nation="POL" athleteid="17316">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="17317" heatid="19299" lane="8" entrytime="00:00:27.11" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="17318" heatid="19386" lane="8" entrytime="00:00:58.21" />
                <RESULT eventid="14243" status="DNS" swimtime="00:00:00.00" resultid="17319" heatid="19407" lane="2" entrytime="00:01:08.32" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="17320" heatid="19459" lane="7" entrytime="00:00:30.11" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="17321" heatid="19552" lane="4" entrytime="00:00:36.82" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-10-19" firstname="Emilia" gender="F" lastname="Sączyńska" nation="POL" athleteid="17505">
              <RESULTS>
                <RESULT eventid="1096" status="DNS" swimtime="00:00:00.00" resultid="17506" heatid="19307" lane="0" entrytime="00:03:08.50" />
                <RESULT eventid="1187" points="356" reactiontime="+81" swimtime="00:00:36.21" resultid="17507" heatid="19339" lane="4" entrytime="00:00:37.50" />
                <RESULT eventid="14225" points="326" reactiontime="+95" swimtime="00:01:22.28" resultid="17508" heatid="19394" lane="9" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="302" reactiontime="+94" swimtime="00:00:36.31" resultid="17509" heatid="19447" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="1457" points="318" reactiontime="+82" swimtime="00:01:20.60" resultid="17510" heatid="19468" lane="1" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="358" reactiontime="+75" swimtime="00:02:47.78" resultid="17511" heatid="19528" lane="5" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.87" />
                    <SPLIT distance="100" swimtime="00:01:19.51" />
                    <SPLIT distance="150" swimtime="00:02:03.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-12-17" firstname="Michał" gender="M" lastname="Nowak" nation="POL" athleteid="17448">
              <RESULTS>
                <RESULT eventid="1113" points="198" reactiontime="+83" swimtime="00:03:07.86" resultid="17449" heatid="19312" lane="2" entrytime="00:03:02.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.45" />
                    <SPLIT distance="100" swimtime="00:01:35.61" />
                    <SPLIT distance="150" swimtime="00:02:25.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="265" reactiontime="+85" swimtime="00:03:07.43" resultid="17450" heatid="19362" lane="6" entrytime="00:03:08.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.00" />
                    <SPLIT distance="100" swimtime="00:01:30.55" />
                    <SPLIT distance="150" swimtime="00:02:19.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="255" reactiontime="+86" swimtime="00:01:19.27" resultid="17451" heatid="19402" lane="6" entrytime="00:01:19.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="302" reactiontime="+81" swimtime="00:01:22.87" resultid="17452" heatid="19439" lane="8" entrytime="00:01:22.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="162" reactiontime="+102" swimtime="00:07:11.46" resultid="17453" heatid="19508" lane="3" entrytime="00:06:57.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.44" />
                    <SPLIT distance="100" swimtime="00:01:50.93" />
                    <SPLIT distance="150" swimtime="00:02:47.05" />
                    <SPLIT distance="200" swimtime="00:03:47.66" />
                    <SPLIT distance="250" swimtime="00:04:41.86" />
                    <SPLIT distance="300" swimtime="00:05:36.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="333" reactiontime="+87" swimtime="00:00:36.42" resultid="17454" heatid="19554" lane="6" entrytime="00:00:36.82" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-30" firstname="Monika" gender="F" lastname="Jarecka-Skorykow" nation="POL" athleteid="17460">
              <RESULTS>
                <RESULT eventid="1062" points="355" reactiontime="+84" swimtime="00:00:32.81" resultid="17461" heatid="19280" lane="7" entrytime="00:00:33.50" />
                <RESULT eventid="14225" points="290" reactiontime="+92" swimtime="00:01:25.53" resultid="17462" heatid="19393" lane="0" entrytime="00:01:25.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="304" reactiontime="+94" swimtime="00:01:32.65" resultid="17463" heatid="19430" lane="1" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="349" reactiontime="+82" swimtime="00:00:40.64" resultid="17464" heatid="19542" lane="7" entrytime="00:00:42.78" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-05-10" firstname="Katarzyna" gender="F" lastname="Czarnecka" nation="POL" athleteid="17424">
              <RESULTS>
                <RESULT eventid="1062" points="449" reactiontime="+62" swimtime="00:00:30.34" resultid="17425" heatid="19282" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="1222" status="DNS" swimtime="00:00:00.00" resultid="17426" heatid="19357" lane="7" entrytime="00:03:25.00" />
                <RESULT eventid="14225" points="322" reactiontime="+69" swimtime="00:01:22.60" resultid="17427" heatid="19389" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="364" reactiontime="+64" swimtime="00:01:27.31" resultid="17428" heatid="19431" lane="7" entrytime="00:01:28.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="390" reactiontime="+57" swimtime="00:00:39.17" resultid="17429" heatid="19544" lane="8" entrytime="00:00:38.66" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-20" firstname="Magdalena" gender="F" lastname="Mostowska" nation="POL" athleteid="17387">
              <RESULTS>
                <RESULT eventid="1165" points="287" reactiontime="+106" swimtime="00:23:13.73" resultid="17388" heatid="19624" lane="6" entrytime="00:25:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.91" />
                    <SPLIT distance="100" swimtime="00:01:27.33" />
                    <SPLIT distance="150" swimtime="00:02:12.44" />
                    <SPLIT distance="200" swimtime="00:02:58.09" />
                    <SPLIT distance="250" swimtime="00:03:44.07" />
                    <SPLIT distance="300" swimtime="00:04:30.36" />
                    <SPLIT distance="350" swimtime="00:05:16.51" />
                    <SPLIT distance="400" swimtime="00:06:02.53" />
                    <SPLIT distance="450" swimtime="00:06:49.28" />
                    <SPLIT distance="500" swimtime="00:07:35.87" />
                    <SPLIT distance="550" swimtime="00:08:22.92" />
                    <SPLIT distance="600" swimtime="00:09:10.01" />
                    <SPLIT distance="650" swimtime="00:09:56.53" />
                    <SPLIT distance="700" swimtime="00:10:43.10" />
                    <SPLIT distance="750" swimtime="00:11:29.94" />
                    <SPLIT distance="800" swimtime="00:12:16.91" />
                    <SPLIT distance="850" swimtime="00:13:03.74" />
                    <SPLIT distance="900" swimtime="00:13:50.80" />
                    <SPLIT distance="950" swimtime="00:14:37.97" />
                    <SPLIT distance="1000" swimtime="00:15:24.93" />
                    <SPLIT distance="1050" swimtime="00:16:12.04" />
                    <SPLIT distance="1100" swimtime="00:16:59.19" />
                    <SPLIT distance="1150" swimtime="00:17:46.40" />
                    <SPLIT distance="1200" swimtime="00:18:33.87" />
                    <SPLIT distance="1250" swimtime="00:19:21.20" />
                    <SPLIT distance="1300" swimtime="00:20:08.23" />
                    <SPLIT distance="1350" swimtime="00:20:55.34" />
                    <SPLIT distance="1400" swimtime="00:21:42.60" />
                    <SPLIT distance="1450" swimtime="00:22:29.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14225" points="195" reactiontime="+105" swimtime="00:01:37.68" resultid="17389" heatid="19391" lane="0" entrytime="00:01:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-10-07" firstname="Daniel" gender="M" lastname="Julian Aguilar" nation="POL" athleteid="17368">
              <RESULTS>
                <RESULT eventid="1079" points="473" reactiontime="+69" swimtime="00:00:26.00" resultid="17369" heatid="19299" lane="1" entrytime="00:00:27.00" />
                <RESULT eventid="1113" points="425" reactiontime="+80" swimtime="00:02:25.80" resultid="17370" heatid="19315" lane="0" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                    <SPLIT distance="100" swimtime="00:01:10.45" />
                    <SPLIT distance="150" swimtime="00:01:52.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="417" reactiontime="+67" swimtime="00:00:29.72" resultid="17371" heatid="19351" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="14243" points="472" reactiontime="+74" swimtime="00:01:04.60" resultid="17372" heatid="19406" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="374" reactiontime="+75" swimtime="00:01:17.17" resultid="17373" heatid="19440" lane="0" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="403" reactiontime="+77" swimtime="00:02:22.92" resultid="17374" heatid="19536" lane="8" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                    <SPLIT distance="100" swimtime="00:01:09.84" />
                    <SPLIT distance="150" swimtime="00:01:46.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="419" reactiontime="+71" swimtime="00:00:33.73" resultid="17375" heatid="19556" lane="8" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-05" firstname="Rafał" gender="M" lastname="Skośkiewicz" nation="POL" athleteid="17336">
              <RESULTS>
                <RESULT eventid="1079" points="398" reactiontime="+80" swimtime="00:00:27.54" resultid="17337" heatid="19295" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="1113" points="405" reactiontime="+91" swimtime="00:02:28.16" resultid="17338" heatid="19316" lane="1" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="100" swimtime="00:01:09.10" />
                    <SPLIT distance="150" swimtime="00:01:54.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="372" reactiontime="+77" swimtime="00:00:30.88" resultid="17339" heatid="19350" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="14243" points="413" reactiontime="+87" swimtime="00:01:07.53" resultid="17340" heatid="19406" lane="3" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="398" reactiontime="+78" swimtime="00:01:06.46" resultid="17341" heatid="19470" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="415" reactiontime="+78" swimtime="00:02:13.20" resultid="17342" heatid="19494" lane="0" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.00" />
                    <SPLIT distance="100" swimtime="00:01:04.96" />
                    <SPLIT distance="150" swimtime="00:01:39.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="363" reactiontime="+80" swimtime="00:02:28.04" resultid="17343" heatid="19536" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.50" />
                    <SPLIT distance="100" swimtime="00:01:10.89" />
                    <SPLIT distance="150" swimtime="00:01:50.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-08-30" firstname="Mirosław" gender="M" lastname="Warchoł" nation="POL" athleteid="17408">
              <RESULTS>
                <RESULT eventid="1079" points="351" reactiontime="+97" swimtime="00:00:28.72" resultid="17409" heatid="19284" lane="1" />
                <RESULT eventid="1113" points="292" reactiontime="+86" swimtime="00:02:45.07" resultid="17410" heatid="19313" lane="6" entrytime="00:02:45.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.86" />
                    <SPLIT distance="100" swimtime="00:01:16.45" />
                    <SPLIT distance="150" swimtime="00:02:08.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="361" reactiontime="+90" swimtime="00:01:03.07" resultid="17411" heatid="19382" lane="2" entrytime="00:01:04.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="308" reactiontime="+72" swimtime="00:01:12.41" resultid="17412" heatid="19470" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="348" reactiontime="+84" swimtime="00:02:21.24" resultid="17413" heatid="19492" lane="6" entrytime="00:02:24.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                    <SPLIT distance="100" swimtime="00:01:08.00" />
                    <SPLIT distance="150" swimtime="00:02:20.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="300" reactiontime="+79" swimtime="00:02:37.71" resultid="17414" heatid="19535" lane="3" entrytime="00:02:44.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                    <SPLIT distance="100" swimtime="00:01:16.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="WMT Meteoryty" number="3">
              <RESULTS>
                <RESULT eventid="1381" points="447" reactiontime="+63" swimtime="00:01:58.37" resultid="17514" heatid="19424" lane="7" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.26" />
                    <SPLIT distance="150" swimtime="00:01:30.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17368" number="1" reactiontime="+63" />
                    <RELAYPOSITION athleteid="17301" number="2" />
                    <RELAYPOSITION athleteid="17440" number="3" reactiontime="+23" />
                    <RELAYPOSITION athleteid="17465" number="4" reactiontime="+65" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="WMT Wielki Wóz" number="4">
              <RESULTS>
                <RESULT eventid="1381" points="493" reactiontime="+79" swimtime="00:01:54.57" resultid="17515" heatid="19424" lane="3" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.85" />
                    <SPLIT distance="100" swimtime="00:01:02.41" />
                    <SPLIT distance="150" swimtime="00:01:29.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17336" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="17415" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="17472" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="17491" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="WMT Kometa Halleya" number="6">
              <RESULTS>
                <RESULT eventid="1548" points="554" reactiontime="+75" swimtime="00:01:40.57" resultid="17517" heatid="19502" lane="5" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.80" />
                    <SPLIT distance="100" swimtime="00:00:49.87" />
                    <SPLIT distance="150" swimtime="00:01:15.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17472" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="17368" number="2" reactiontime="+19" />
                    <RELAYPOSITION athleteid="17440" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="17491" number="4" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="WMT Czarna Dziura" number="7">
              <RESULTS>
                <RESULT eventid="1548" points="377" reactiontime="+74" swimtime="00:01:54.32" resultid="17518" heatid="19501" lane="6" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.90" />
                    <SPLIT distance="100" swimtime="00:00:59.33" />
                    <SPLIT distance="150" swimtime="00:01:27.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17465" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="17396" number="2" reactiontime="+20" />
                    <RELAYPOSITION athleteid="17351" number="3" reactiontime="+5" />
                    <RELAYPOSITION athleteid="17301" number="4" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="WMT Stella Timea" number="5">
              <RESULTS>
                <RESULT eventid="1358" points="297" reactiontime="+83" swimtime="00:02:34.74" resultid="17516" heatid="19420" lane="1" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.91" />
                    <SPLIT distance="100" swimtime="00:01:35.68" />
                    <SPLIT distance="150" swimtime="00:02:10.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17327" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="17478" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="17360" number="3" />
                    <RELAYPOSITION athleteid="17496" number="4" reactiontime="+63" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="WMT Droga Mleczna" number="8">
              <RESULTS>
                <RESULT eventid="1525" points="433" reactiontime="+70" swimtime="00:02:04.53" resultid="17519" heatid="19498" lane="1" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.87" />
                    <SPLIT distance="100" swimtime="00:01:06.47" />
                    <SPLIT distance="150" swimtime="00:01:37.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17424" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="17382" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="17460" number="3" />
                    <RELAYPOSITION athleteid="17444" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="WMT Zorza Polarna" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="544" reactiontime="+77" swimtime="00:01:48.47" resultid="17512" heatid="19322" lane="4" entrytime="00:01:47.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.81" />
                    <SPLIT distance="100" swimtime="00:00:53.29" />
                    <SPLIT distance="150" swimtime="00:01:24.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17484" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="17376" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="17424" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="17472" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="WMT Kasjopea" number="2">
              <RESULTS>
                <RESULT eventid="1130" points="361" reactiontime="+87" swimtime="00:02:04.29" resultid="17513" heatid="19321" lane="2" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                    <SPLIT distance="100" swimtime="00:01:08.35" />
                    <SPLIT distance="150" swimtime="00:01:36.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17460" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="17327" number="2" reactiontime="+38" />
                    <RELAYPOSITION athleteid="17465" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="17402" number="4" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" name="WMT Totalny Kosmos" number="9">
              <RESULTS>
                <RESULT eventid="1698" points="592" reactiontime="+76" swimtime="00:01:55.68" resultid="17520" heatid="19564" lane="4" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.19" />
                    <SPLIT distance="100" swimtime="00:01:01.66" />
                    <SPLIT distance="150" swimtime="00:01:27.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17472" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="17444" number="2" reactiontime="+22" />
                    <RELAYPOSITION athleteid="17484" number="3" reactiontime="+18" />
                    <RELAYPOSITION athleteid="17376" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="WMT Asteroidy" number="10">
              <RESULTS>
                <RESULT eventid="1698" points="382" reactiontime="+78" swimtime="00:02:13.87" resultid="17521" heatid="19563" lane="5" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.20" />
                    <SPLIT distance="100" swimtime="00:01:10.26" />
                    <SPLIT distance="150" swimtime="00:01:41.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17336" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="17424" number="2" reactiontime="+29" />
                    <RELAYPOSITION athleteid="17455" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="17460" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="WMT Galaktyka Andromedy" number="11">
              <RESULTS>
                <RESULT eventid="1698" points="285" reactiontime="+67" swimtime="00:02:27.50" resultid="17522" heatid="19562" lane="6" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                    <SPLIT distance="100" swimtime="00:01:06.46" />
                    <SPLIT distance="150" swimtime="00:01:51.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17368" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="17448" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="17478" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="17327" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="SLA" clubid="14451" name="Weteran Zabrze">
          <CONTACT city="ZABRZE" email="weteranzabrze@op.pl" name="BOSOWSKI  WŁODZIMIERZ" street="ŚW.  JANA" zip="41803" />
          <ATHLETES>
            <ATHLETE birthdate="1943-12-02" firstname="Renata" gender="F" lastname="Bastek" nation="POL" license="102611600023" athleteid="14456">
              <RESULTS>
                <RESULT eventid="1062" points="217" reactiontime="+86" swimtime="00:00:38.64" resultid="14457" heatid="19278" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1187" points="146" reactiontime="+78" swimtime="00:00:48.66" resultid="14458" heatid="19338" lane="0" entrytime="00:00:46.00" />
                <RESULT eventid="1256" points="197" swimtime="00:01:27.49" resultid="14459" heatid="19369" lane="9" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="101" reactiontime="+87" swimtime="00:00:52.34" resultid="14460" heatid="19445" lane="2" entrytime="00:00:50.00" />
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="14461" heatid="19695" lane="3" entrytime="00:07:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-07-16" firstname="Ewald" gender="M" lastname="Bastek" nation="POL" license="102611700022" athleteid="14452">
              <RESULTS>
                <RESULT eventid="1113" points="111" reactiontime="+104" swimtime="00:03:47.65" resultid="14453" heatid="19310" lane="5" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.58" />
                    <SPLIT distance="100" swimtime="00:01:55.39" />
                    <SPLIT distance="150" swimtime="00:02:59.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="111" reactiontime="+105" swimtime="00:01:44.62" resultid="14454" heatid="19399" lane="9" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="127" reactiontime="+104" swimtime="00:03:17.20" resultid="14455" heatid="19487" lane="7" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-07-27" firstname="Danuta" gender="F" lastname="Skorupa" nation="POL" license="102611600020" athleteid="14518">
              <RESULTS>
                <RESULT eventid="1187" points="53" reactiontime="+94" swimtime="00:01:08.14" resultid="14519" heatid="19336" lane="4" entrytime="00:00:59.98" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-29" firstname="Wiesław" gender="M" lastname="Kornicki" nation="POL" license="102611700015" athleteid="14520">
              <RESULTS>
                <RESULT eventid="1079" points="198" swimtime="00:00:34.74" resultid="14521" heatid="19291" lane="9" entrytime="00:00:32.00" />
                <RESULT eventid="1273" points="187" reactiontime="+86" swimtime="00:01:18.45" resultid="14522" heatid="19378" lane="8" entrytime="00:01:16.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="148" reactiontime="+88" swimtime="00:01:35.05" resultid="14523" heatid="19400" lane="9" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="197" reactiontime="+90" swimtime="00:00:37.46" resultid="14524" heatid="19454" lane="8" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-08-23" firstname="Danuta" gender="F" lastname="Karczewska" nation="POL" athleteid="14485">
              <RESULTS>
                <RESULT eventid="1062" points="111" swimtime="00:00:48.27" resultid="14486" heatid="19277" lane="9" entrytime="00:00:45.80" />
                <RESULT eventid="1147" reactiontime="+121" status="OTL" swimtime="00:18:40.46" resultid="14487" heatid="19594" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.94" />
                    <SPLIT distance="100" swimtime="00:02:03.32" />
                    <SPLIT distance="150" swimtime="00:03:12.77" />
                    <SPLIT distance="200" swimtime="00:04:24.25" />
                    <SPLIT distance="250" swimtime="00:05:34.51" />
                    <SPLIT distance="300" swimtime="00:06:44.54" />
                    <SPLIT distance="350" swimtime="00:07:56.91" />
                    <SPLIT distance="400" swimtime="00:09:09.28" />
                    <SPLIT distance="450" swimtime="00:10:21.46" />
                    <SPLIT distance="500" swimtime="00:11:33.67" />
                    <SPLIT distance="550" swimtime="00:12:46.31" />
                    <SPLIT distance="600" swimtime="00:13:58.77" />
                    <SPLIT distance="650" swimtime="00:15:11.65" />
                    <SPLIT distance="700" swimtime="00:16:23.49" />
                    <SPLIT distance="750" swimtime="00:17:35.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="96" reactiontime="+109" swimtime="00:01:51.02" resultid="14488" heatid="19368" lane="1" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="74" reactiontime="+119" swimtime="00:04:23.31" resultid="14489" heatid="19479" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.00" />
                    <SPLIT distance="100" swimtime="00:02:03.15" />
                    <SPLIT distance="150" swimtime="00:03:15.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="87" reactiontime="+142" swimtime="00:08:48.38" resultid="14490" heatid="19694" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.43" />
                    <SPLIT distance="100" swimtime="00:02:02.79" />
                    <SPLIT distance="150" swimtime="00:03:09.45" />
                    <SPLIT distance="200" swimtime="00:04:17.71" />
                    <SPLIT distance="250" swimtime="00:05:26.16" />
                    <SPLIT distance="300" swimtime="00:06:34.69" />
                    <SPLIT distance="350" swimtime="00:07:43.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-11-02" firstname="Beata" gender="F" lastname="Sulewska" nation="POL" license="102611600016" athleteid="14525">
              <RESULTS>
                <RESULT comment="Wynik lepszy od Rekordu Polski na 800m i 400m" eventid="1147" points="492" reactiontime="+94" swimtime="00:10:07.02" resultid="14526" heatid="19596" lane="6" entrytime="00:10:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                    <SPLIT distance="100" swimtime="00:01:12.44" />
                    <SPLIT distance="150" swimtime="00:01:50.35" />
                    <SPLIT distance="200" swimtime="00:02:28.62" />
                    <SPLIT distance="250" swimtime="00:03:06.99" />
                    <SPLIT distance="300" swimtime="00:03:45.27" />
                    <SPLIT distance="350" swimtime="00:04:23.45" />
                    <SPLIT distance="400" swimtime="00:05:01.68" />
                    <SPLIT distance="450" swimtime="00:05:39.80" />
                    <SPLIT distance="500" swimtime="00:06:18.08" />
                    <SPLIT distance="550" swimtime="00:06:56.39" />
                    <SPLIT distance="600" swimtime="00:07:34.89" />
                    <SPLIT distance="650" swimtime="00:08:13.20" />
                    <SPLIT distance="700" swimtime="00:08:51.42" />
                    <SPLIT distance="750" swimtime="00:09:29.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="424" reactiontime="+90" swimtime="00:02:59.06" resultid="14527" heatid="19358" lane="6" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.13" />
                    <SPLIT distance="100" swimtime="00:01:25.39" />
                    <SPLIT distance="150" swimtime="00:02:11.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="438" reactiontime="+79" swimtime="00:01:22.11" resultid="14528" heatid="19432" lane="0" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.91" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1555" points="444" reactiontime="+92" swimtime="00:05:39.97" resultid="14529" heatid="19505" lane="6" entrytime="00:05:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                    <SPLIT distance="100" swimtime="00:01:17.06" />
                    <SPLIT distance="150" swimtime="00:02:03.00" />
                    <SPLIT distance="200" swimtime="00:02:48.60" />
                    <SPLIT distance="250" swimtime="00:03:35.60" />
                    <SPLIT distance="300" swimtime="00:04:22.33" />
                    <SPLIT distance="350" swimtime="00:05:02.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" status="DNS" swimtime="00:00:00.00" resultid="14530" heatid="19544" lane="9" entrytime="00:00:40.00" />
                <RESULT comment="Wynik lepszy od Rekordu Polski" eventid="1721" points="479" reactiontime="+88" swimtime="00:04:59.65" resultid="14531" heatid="19698" lane="6" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.24" />
                    <SPLIT distance="100" swimtime="00:01:10.66" />
                    <SPLIT distance="150" swimtime="00:01:48.00" />
                    <SPLIT distance="200" swimtime="00:02:25.90" />
                    <SPLIT distance="250" swimtime="00:03:04.34" />
                    <SPLIT distance="300" swimtime="00:03:43.45" />
                    <SPLIT distance="350" swimtime="00:04:22.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-02-25" firstname="Bernard" gender="M" lastname="Poloczek" nation="POL" athleteid="14496">
              <RESULTS>
                <RESULT eventid="1205" points="139" reactiontime="+70" swimtime="00:00:42.81" resultid="14497" heatid="19345" lane="7" entrytime="00:00:44.11" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="14498" heatid="19451" lane="5" entrytime="00:00:46.20" />
                <RESULT eventid="1474" points="130" reactiontime="+71" swimtime="00:01:36.37" resultid="14499" heatid="19473" lane="9" entrytime="00:01:35.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="114" reactiontime="+70" swimtime="00:03:37.61" resultid="14500" heatid="19533" lane="9" entrytime="00:03:46.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.82" />
                    <SPLIT distance="100" swimtime="00:01:46.57" />
                    <SPLIT distance="150" swimtime="00:02:42.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-11" firstname="Jan" gender="M" lastname="Barucha" nation="POL" license="102611700021" athleteid="14511">
              <RESULTS>
                <RESULT eventid="1079" points="273" reactiontime="+73" swimtime="00:00:31.20" resultid="14512" heatid="19291" lane="8" entrytime="00:00:31.68" />
                <RESULT eventid="1205" points="165" reactiontime="+76" swimtime="00:00:40.44" resultid="14513" heatid="19346" lane="6" entrytime="00:00:40.24" />
                <RESULT eventid="1273" points="237" reactiontime="+75" swimtime="00:01:12.56" resultid="14514" heatid="19379" lane="0" entrytime="00:01:12.60" />
                <RESULT eventid="1440" points="207" reactiontime="+77" swimtime="00:00:36.80" resultid="14515" heatid="19453" lane="9" entrytime="00:00:39.89" />
                <RESULT eventid="1474" points="175" reactiontime="+75" swimtime="00:01:27.45" resultid="14516" heatid="19473" lane="6" entrytime="00:01:28.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="155" reactiontime="+81" swimtime="00:03:16.62" resultid="14517" heatid="19534" lane="0" entrytime="00:03:15.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.71" />
                    <SPLIT distance="100" swimtime="00:01:32.34" />
                    <SPLIT distance="150" swimtime="00:02:24.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-03-12" firstname="Krystyna" gender="F" lastname="Fecica" nation="POL" license="102611600019" athleteid="14477">
              <RESULTS>
                <RESULT eventid="1165" points="112" reactiontime="+96" swimtime="00:31:47.16" resultid="14478" heatid="19624" lane="8" entrytime="00:34:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.52" />
                    <SPLIT distance="100" swimtime="00:01:52.47" />
                    <SPLIT distance="150" swimtime="00:02:54.77" />
                    <SPLIT distance="200" swimtime="00:03:56.90" />
                    <SPLIT distance="250" swimtime="00:04:58.76" />
                    <SPLIT distance="300" swimtime="00:06:02.42" />
                    <SPLIT distance="350" swimtime="00:07:07.44" />
                    <SPLIT distance="400" swimtime="00:08:12.81" />
                    <SPLIT distance="450" swimtime="00:10:21.07" />
                    <SPLIT distance="500" swimtime="00:11:25.34" />
                    <SPLIT distance="550" swimtime="00:12:32.40" />
                    <SPLIT distance="600" swimtime="00:13:36.53" />
                    <SPLIT distance="650" swimtime="00:14:39.41" />
                    <SPLIT distance="700" swimtime="00:17:54.71" />
                    <SPLIT distance="750" swimtime="00:20:02.13" />
                    <SPLIT distance="800" swimtime="00:21:07.81" />
                    <SPLIT distance="850" swimtime="00:23:17.68" />
                    <SPLIT distance="900" swimtime="00:24:22.03" />
                    <SPLIT distance="950" swimtime="00:25:27.12" />
                    <SPLIT distance="1000" swimtime="00:26:31.41" />
                    <SPLIT distance="1050" swimtime="00:27:34.60" />
                    <SPLIT distance="1100" swimtime="00:28:37.68" />
                    <SPLIT distance="1150" swimtime="00:30:46.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="91" reactiontime="+103" swimtime="00:04:25.16" resultid="14479" heatid="19411" lane="3" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.38" />
                    <SPLIT distance="100" swimtime="00:02:05.80" />
                    <SPLIT distance="150" swimtime="00:03:15.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-11-29" firstname="Daniel" gender="M" lastname="Fecica" nation="POL" license="102611700018" athleteid="14473">
              <RESULTS>
                <RESULT eventid="1239" points="167" reactiontime="+116" swimtime="00:03:38.64" resultid="14474" heatid="19360" lane="3" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.31" />
                    <SPLIT distance="100" swimtime="00:01:45.56" />
                    <SPLIT distance="150" swimtime="00:02:43.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="169" reactiontime="+108" swimtime="00:01:40.53" resultid="14475" heatid="19435" lane="5" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="177" reactiontime="+106" swimtime="00:00:44.97" resultid="14476" heatid="19549" lane="3" entrytime="00:00:45.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-03-11" firstname="Bartłomiej" gender="M" lastname="Bober" nation="POL" athleteid="14480">
              <RESULTS>
                <RESULT eventid="1079" points="449" reactiontime="+83" swimtime="00:00:26.44" resultid="14481" heatid="19302" lane="2" entrytime="00:00:25.50" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="14482" heatid="19387" lane="0" entrytime="00:00:56.50" />
                <RESULT eventid="1508" points="454" reactiontime="+79" swimtime="00:02:09.22" resultid="14483" heatid="19495" lane="7" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.59" />
                    <SPLIT distance="100" swimtime="00:01:02.07" />
                    <SPLIT distance="150" swimtime="00:01:35.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="442" reactiontime="+84" swimtime="00:04:38.46" resultid="14484" heatid="19707" lane="2" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                    <SPLIT distance="100" swimtime="00:01:07.73" />
                    <SPLIT distance="150" swimtime="00:01:43.39" />
                    <SPLIT distance="200" swimtime="00:02:19.01" />
                    <SPLIT distance="250" swimtime="00:02:54.58" />
                    <SPLIT distance="300" swimtime="00:03:30.33" />
                    <SPLIT distance="350" swimtime="00:04:05.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14189" points="477" swimtime="00:09:27.45" resultid="16545" heatid="19618" lane="0" entrytime="00:09:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.78" />
                    <SPLIT distance="100" swimtime="00:01:06.36" />
                    <SPLIT distance="150" swimtime="00:01:41.69" />
                    <SPLIT distance="200" swimtime="00:02:17.02" />
                    <SPLIT distance="250" swimtime="00:02:52.83" />
                    <SPLIT distance="300" swimtime="00:03:28.96" />
                    <SPLIT distance="350" swimtime="00:04:05.18" />
                    <SPLIT distance="400" swimtime="00:04:40.96" />
                    <SPLIT distance="450" swimtime="00:05:17.03" />
                    <SPLIT distance="500" swimtime="00:05:52.92" />
                    <SPLIT distance="550" swimtime="00:06:29.03" />
                    <SPLIT distance="600" swimtime="00:07:05.34" />
                    <SPLIT distance="650" swimtime="00:07:41.50" />
                    <SPLIT distance="700" swimtime="00:08:17.81" />
                    <SPLIT distance="750" swimtime="00:08:53.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="434" reactiontime="+90" swimtime="00:05:10.88" resultid="16546" heatid="19512" lane="2" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                    <SPLIT distance="100" swimtime="00:01:11.27" />
                    <SPLIT distance="150" swimtime="00:01:54.42" />
                    <SPLIT distance="200" swimtime="00:02:34.99" />
                    <SPLIT distance="250" swimtime="00:03:17.83" />
                    <SPLIT distance="300" swimtime="00:04:00.20" />
                    <SPLIT distance="350" swimtime="00:04:36.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="406" reactiontime="+81" swimtime="00:01:04.93" resultid="16547" heatid="19524" lane="3" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-04-14" firstname="Gabriela" gender="F" lastname="Molenda" nation="POL" athleteid="14507">
              <RESULTS>
                <RESULT eventid="1147" reactiontime="+108" status="OTL" swimtime="00:15:20.57" resultid="14508" heatid="19595" lane="7" entrytime="00:13:46.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.93" />
                    <SPLIT distance="100" swimtime="00:01:40.80" />
                    <SPLIT distance="150" swimtime="00:02:37.12" />
                    <SPLIT distance="200" swimtime="00:03:34.50" />
                    <SPLIT distance="250" swimtime="00:04:31.36" />
                    <SPLIT distance="300" swimtime="00:05:28.98" />
                    <SPLIT distance="350" swimtime="00:06:26.72" />
                    <SPLIT distance="400" swimtime="00:07:24.97" />
                    <SPLIT distance="450" swimtime="00:08:24.76" />
                    <SPLIT distance="500" swimtime="00:09:23.59" />
                    <SPLIT distance="550" swimtime="00:10:22.53" />
                    <SPLIT distance="600" swimtime="00:11:21.01" />
                    <SPLIT distance="650" swimtime="00:12:21.28" />
                    <SPLIT distance="700" swimtime="00:13:21.48" />
                    <SPLIT distance="750" swimtime="00:14:21.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="103" reactiontime="+75" swimtime="00:00:54.76" resultid="14509" heatid="19337" lane="5" entrytime="00:00:48.70" />
                <RESULT eventid="1721" points="150" reactiontime="+105" swimtime="00:07:20.89" resultid="14510" heatid="19697" lane="0" entrytime="00:06:42.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.54" />
                    <SPLIT distance="100" swimtime="00:01:41.15" />
                    <SPLIT distance="150" swimtime="00:02:36.96" />
                    <SPLIT distance="200" swimtime="00:03:33.24" />
                    <SPLIT distance="250" swimtime="00:04:29.83" />
                    <SPLIT distance="300" swimtime="00:05:26.66" />
                    <SPLIT distance="350" swimtime="00:06:24.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-05-22" firstname="Włodzimierz" gender="M" lastname="Bosowski" nation="POL" license="102611700014" athleteid="14462">
              <RESULTS>
                <RESULT eventid="1079" points="130" reactiontime="+109" swimtime="00:00:39.90" resultid="14463" heatid="19286" lane="3" entrytime="00:00:38.50" />
                <RESULT eventid="1440" points="81" reactiontime="+109" swimtime="00:00:50.31" resultid="14464" heatid="19452" lane="1" entrytime="00:00:43.00" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="14465" heatid="19518" lane="0" entrytime="00:01:53.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-02-18" firstname="Genowefa" gender="F" lastname="Drużyńska" nation="POL" athleteid="14469">
              <RESULTS>
                <RESULT eventid="1222" points="98" reactiontime="+100" swimtime="00:04:50.95" resultid="14470" heatid="19355" lane="7" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:19.18" />
                    <SPLIT distance="150" swimtime="00:03:37.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="104" reactiontime="+109" swimtime="00:02:12.25" resultid="14471" heatid="19427" lane="4" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="132" reactiontime="+104" swimtime="00:00:56.17" resultid="14472" heatid="19539" lane="6" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-05-23" firstname="Janina" gender="F" lastname="Bosowska" nation="POL" license="102611600024" athleteid="14466">
              <RESULTS>
                <RESULT eventid="14225" points="86" reactiontime="+106" swimtime="00:02:08.27" resultid="14467" heatid="19390" lane="2" entrytime="00:01:56.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="138" reactiontime="+106" swimtime="00:00:55.40" resultid="14468" heatid="19539" lane="4" entrytime="00:00:56.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-10-05" firstname="Barbara" gender="F" lastname="Brendler" nation="POL" license="102611600017" athleteid="14491">
              <RESULTS>
                <RESULT eventid="1062" points="182" reactiontime="+103" swimtime="00:00:40.96" resultid="14492" heatid="19277" lane="3" entrytime="00:00:41.00" />
                <RESULT eventid="1256" points="143" reactiontime="+115" swimtime="00:01:37.14" resultid="14493" heatid="19368" lane="3" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="116" reactiontime="+112" swimtime="00:03:47.04" resultid="14494" heatid="19480" lane="3" entrytime="00:03:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.27" />
                    <SPLIT distance="100" swimtime="00:01:49.21" />
                    <SPLIT distance="150" swimtime="00:02:48.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="66" reactiontime="+93" swimtime="00:04:54.02" resultid="14495" heatid="19526" lane="3" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.77" />
                    <SPLIT distance="100" swimtime="00:02:24.41" />
                    <SPLIT distance="150" swimtime="00:03:43.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-05-25" firstname="Wojciech" gender="M" lastname="Nowiński" nation="POL" athleteid="14501">
              <RESULTS>
                <RESULT eventid="1079" points="294" reactiontime="+73" swimtime="00:00:30.44" resultid="14502" heatid="19296" lane="9" entrytime="00:00:29.00" />
                <RESULT eventid="1205" points="230" reactiontime="+67" swimtime="00:00:36.26" resultid="14503" heatid="19350" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="1273" points="272" reactiontime="+92" swimtime="00:01:09.29" resultid="14504" heatid="19382" lane="1" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="14505" heatid="19454" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1474" points="214" swimtime="00:01:21.76" resultid="14506" heatid="19476" lane="9" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1381" points="173" reactiontime="+75" swimtime="00:02:42.28" resultid="14535" heatid="19421" lane="5" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                    <SPLIT distance="100" swimtime="00:01:26.06" />
                    <SPLIT distance="150" swimtime="00:02:03.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14511" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="14473" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="14520" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="14452" number="4" reactiontime="+71" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="6">
              <RESULTS>
                <RESULT eventid="1548" points="182" reactiontime="+103" swimtime="00:02:25.67" resultid="14537" heatid="19499" lane="5" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.25" />
                    <SPLIT distance="100" swimtime="00:01:18.51" />
                    <SPLIT distance="150" swimtime="00:01:53.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14473" number="1" reactiontime="+103" />
                    <RELAYPOSITION athleteid="14452" number="2" reactiontime="+75" />
                    <RELAYPOSITION athleteid="14520" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="14511" number="4" reactiontime="+14" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="F" number="3">
              <RESULTS>
                <RESULT eventid="1358" points="149" reactiontime="+70" swimtime="00:03:14.68" resultid="14534" heatid="19419" lane="5" entrytime="00:03:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.71" />
                    <SPLIT distance="100" swimtime="00:01:42.48" />
                    <SPLIT distance="150" swimtime="00:02:34.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14477" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="14466" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="14456" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="14491" number="4" reactiontime="+66" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="F" number="5">
              <RESULTS>
                <RESULT eventid="1525" points="140" reactiontime="+90" swimtime="00:03:01.29" resultid="14536" heatid="19498" lane="9" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.51" />
                    <SPLIT distance="100" swimtime="00:01:40.06" />
                    <SPLIT distance="150" swimtime="00:02:22.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14477" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="14466" number="2" reactiontime="+54" />
                    <RELAYPOSITION athleteid="14491" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="14456" number="4" reactiontime="+20" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="146" reactiontime="+89" swimtime="00:02:48.00" resultid="14532" heatid="19320" lane="0" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.99" />
                    <SPLIT distance="100" swimtime="00:01:25.79" />
                    <SPLIT distance="150" swimtime="00:02:07.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14473" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="14466" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="14491" number="3" />
                    <RELAYPOSITION athleteid="14462" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1130" points="278" reactiontime="+84" swimtime="00:02:15.56" resultid="14533" heatid="19320" lane="7" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.12" />
                    <SPLIT distance="150" swimtime="00:01:44.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14456" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="14520" number="2" />
                    <RELAYPOSITION athleteid="14525" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="14511" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" number="7">
              <RESULTS>
                <RESULT eventid="1698" points="180" reactiontime="+69" swimtime="00:02:51.99" resultid="14538" heatid="19562" lane="9" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.09" />
                    <SPLIT distance="100" swimtime="00:01:33.43" />
                    <SPLIT distance="150" swimtime="00:02:10.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14456" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="14473" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="14520" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="14491" number="4" reactiontime="+85" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="14734" name="WKS Śląsk Wrocław">
          <CONTACT email="marrot68@wp.pl" name="Rother Marek" />
          <ATHLETES>
            <ATHLETE birthdate="1968-05-21" firstname="Marek" gender="M" lastname="Rother" nation="POL" athleteid="14735">
              <RESULTS>
                <RESULT eventid="1205" points="433" reactiontime="+70" swimtime="00:00:29.36" resultid="14736" heatid="19350" lane="3" entrytime="00:00:31.50" />
                <RESULT eventid="14243" points="421" reactiontime="+74" swimtime="00:01:07.10" resultid="14737" heatid="19406" lane="9" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="425" reactiontime="+71" swimtime="00:01:05.03" resultid="14738" heatid="19477" lane="2" entrytime="00:01:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="415" reactiontime="+72" swimtime="00:02:21.54" resultid="14739" heatid="19537" lane="1" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                    <SPLIT distance="100" swimtime="00:01:07.92" />
                    <SPLIT distance="150" swimtime="00:01:44.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="18345" name="Wyższa Szkoła Biznesu w Dąbrowie Górniczej">
          <ATHLETES>
            <ATHLETE birthdate="1993-02-05" firstname="Kacper" gender="M" lastname="Kaproń" nation="SVK" athleteid="18565">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="18566" heatid="19297" lane="0" entrytime="00:00:28.00" />
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="18567" heatid="19312" lane="6" entrytime="00:03:00.00" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="18568" heatid="19349" lane="8" entrytime="00:00:34.00" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="18569" heatid="19363" lane="2" entrytime="00:03:00.00" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="18570" heatid="19438" lane="6" entrytime="00:01:25.00" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="18571" heatid="19474" lane="1" entrytime="00:01:25.00" />
                <RESULT eventid="1647" points="270" reactiontime="+64" swimtime="00:02:43.36" resultid="18572" heatid="19535" lane="9" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.87" />
                    <SPLIT distance="100" swimtime="00:01:19.29" />
                    <SPLIT distance="150" swimtime="00:02:01.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="406" reactiontime="+76" swimtime="00:00:34.08" resultid="18573" heatid="19557" lane="4" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="18344" name="Wyższa Szkoła Humanitas w Sosnowcu">
          <ATHLETES>
            <ATHLETE birthdate="1996-03-24" firstname="Kinga" gender="F" lastname="Pluta" nation="SVK" athleteid="18574">
              <RESULTS>
                <RESULT eventid="1062" status="DNS" swimtime="00:00:00.00" resultid="18575" heatid="19280" lane="0" entrytime="00:00:34.00" />
                <RESULT eventid="1096" status="DNS" swimtime="00:00:00.00" resultid="18576" heatid="19306" lane="4" entrytime="00:03:15.00" />
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="18577" heatid="19339" lane="3" entrytime="00:00:38.00" />
                <RESULT eventid="1222" points="395" reactiontime="+87" swimtime="00:03:03.34" resultid="18578" heatid="19358" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.72" />
                    <SPLIT distance="100" swimtime="00:01:26.46" />
                    <SPLIT distance="150" swimtime="00:02:14.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" status="DNS" swimtime="00:00:00.00" resultid="18579" heatid="19431" lane="8" entrytime="00:01:30.00" />
                <RESULT eventid="1457" status="DNS" swimtime="00:00:00.00" resultid="18580" heatid="19467" lane="1" entrytime="00:01:28.00" />
                <RESULT eventid="1630" points="302" reactiontime="+87" swimtime="00:02:57.71" resultid="18581" heatid="19529" lane="0" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.50" />
                    <SPLIT distance="100" swimtime="00:01:26.88" />
                    <SPLIT distance="150" swimtime="00:02:12.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="446" reactiontime="+88" swimtime="00:00:37.46" resultid="18582" heatid="19544" lane="5" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="SVK" clubid="14684" name="ŠPK Kúpele Piešťany">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1948-11-25" firstname="Karol" gender="M" lastname="Kantek" nation="SVK" license="SVK18954" athleteid="14699">
              <RESULTS>
                <RESULT eventid="1079" points="282" reactiontime="+74" swimtime="00:00:30.89" resultid="14700" heatid="19291" lane="6" entrytime="00:00:31.30" />
                <RESULT comment="O4 - Start wykonany przed sygnłem (przedwczesny start) (Time: 11:03)" eventid="1273" reactiontime="+65" status="DSQ" swimtime="00:01:11.55" resultid="14701" heatid="19378" lane="4" entrytime="00:01:13.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="230" reactiontime="+94" swimtime="00:00:35.56" resultid="14702" heatid="19455" lane="1" entrytime="00:00:34.30" />
                <RESULT eventid="1681" points="222" reactiontime="+93" swimtime="00:00:41.70" resultid="14703" heatid="19550" lane="4" entrytime="00:00:42.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-10-27" firstname="Pavol" gender="M" lastname="Škodný" nation="SVK" license="SVK12519" athleteid="14693">
              <RESULTS>
                <RESULT eventid="14207" points="310" reactiontime="+114" swimtime="00:20:52.08" resultid="14694" heatid="19622" lane="2" entrytime="00:21:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.54" />
                    <SPLIT distance="100" swimtime="00:01:14.86" />
                    <SPLIT distance="150" swimtime="00:01:55.37" />
                    <SPLIT distance="200" swimtime="00:02:36.58" />
                    <SPLIT distance="250" swimtime="00:03:18.24" />
                    <SPLIT distance="300" swimtime="00:04:00.32" />
                    <SPLIT distance="350" swimtime="00:04:42.68" />
                    <SPLIT distance="400" swimtime="00:05:24.47" />
                    <SPLIT distance="450" swimtime="00:06:06.95" />
                    <SPLIT distance="500" swimtime="00:07:30.91" />
                    <SPLIT distance="550" swimtime="00:08:13.16" />
                    <SPLIT distance="600" swimtime="00:09:38.13" />
                    <SPLIT distance="650" swimtime="00:10:20.49" />
                    <SPLIT distance="700" swimtime="00:11:02.78" />
                    <SPLIT distance="750" swimtime="00:11:44.98" />
                    <SPLIT distance="800" swimtime="00:12:28.05" />
                    <SPLIT distance="850" swimtime="00:13:10.68" />
                    <SPLIT distance="900" swimtime="00:13:53.34" />
                    <SPLIT distance="950" swimtime="00:14:35.80" />
                    <SPLIT distance="1000" swimtime="00:15:17.55" />
                    <SPLIT distance="1050" swimtime="00:16:00.14" />
                    <SPLIT distance="1100" swimtime="00:16:42.46" />
                    <SPLIT distance="1150" swimtime="00:17:24.88" />
                    <SPLIT distance="1200" swimtime="00:18:07.27" />
                    <SPLIT distance="1250" swimtime="00:18:49.62" />
                    <SPLIT distance="1300" swimtime="00:19:31.45" />
                    <SPLIT distance="1350" swimtime="00:20:13.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="274" reactiontime="+107" swimtime="00:02:47.05" resultid="14695" heatid="19416" lane="3" entrytime="00:02:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                    <SPLIT distance="100" swimtime="00:01:17.22" />
                    <SPLIT distance="150" swimtime="00:02:01.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="311" reactiontime="+75" swimtime="00:01:12.20" resultid="14696" heatid="19476" lane="6" entrytime="00:01:11.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="323" reactiontime="+107" swimtime="00:05:43.21" resultid="14697" heatid="19511" lane="7" entrytime="00:05:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.04" />
                    <SPLIT distance="100" swimtime="00:01:17.61" />
                    <SPLIT distance="150" swimtime="00:02:01.07" />
                    <SPLIT distance="200" swimtime="00:02:44.46" />
                    <SPLIT distance="250" swimtime="00:03:35.54" />
                    <SPLIT distance="300" swimtime="00:04:23.97" />
                    <SPLIT distance="350" swimtime="00:05:05.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="299" reactiontime="+77" swimtime="00:02:37.93" resultid="14698" heatid="19536" lane="6" entrytime="00:02:35.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                    <SPLIT distance="100" swimtime="00:01:15.90" />
                    <SPLIT distance="150" swimtime="00:01:57.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-04-03" firstname="Juraj" gender="M" lastname="Horil" nation="SVK" license="SVK14912" athleteid="14704">
              <RESULTS>
                <RESULT eventid="1079" points="294" swimtime="00:00:30.44" resultid="14705" heatid="19292" lane="0" entrytime="00:00:30.50" />
                <RESULT eventid="14189" points="215" reactiontime="+92" swimtime="00:12:19.99" resultid="14706" heatid="19616" lane="7" entrytime="00:11:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                    <SPLIT distance="100" swimtime="00:01:17.86" />
                    <SPLIT distance="150" swimtime="00:02:01.16" />
                    <SPLIT distance="200" swimtime="00:02:46.03" />
                    <SPLIT distance="250" swimtime="00:03:31.96" />
                    <SPLIT distance="300" swimtime="00:04:17.94" />
                    <SPLIT distance="350" swimtime="00:05:04.92" />
                    <SPLIT distance="400" swimtime="00:05:52.29" />
                    <SPLIT distance="450" swimtime="00:06:39.88" />
                    <SPLIT distance="500" swimtime="00:07:28.01" />
                    <SPLIT distance="550" swimtime="00:08:16.23" />
                    <SPLIT distance="600" swimtime="00:09:05.13" />
                    <SPLIT distance="650" swimtime="00:09:54.38" />
                    <SPLIT distance="700" swimtime="00:10:43.77" />
                    <SPLIT distance="750" swimtime="00:11:32.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="290" reactiontime="+93" swimtime="00:03:01.92" resultid="14707" heatid="19362" lane="5" entrytime="00:03:04.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.27" />
                    <SPLIT distance="100" swimtime="00:01:23.91" />
                    <SPLIT distance="150" swimtime="00:02:12.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14243" points="255" reactiontime="+86" swimtime="00:01:19.30" resultid="14708" heatid="19402" lane="5" entrytime="00:01:18.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="325" reactiontime="+88" swimtime="00:01:20.87" resultid="14709" heatid="19439" lane="6" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="320" reactiontime="+82" swimtime="00:00:36.90" resultid="14710" heatid="19554" lane="4" entrytime="00:00:36.60" />
                <RESULT eventid="1744" points="219" reactiontime="+94" swimtime="00:05:51.70" resultid="14711" heatid="19702" lane="4" entrytime="00:06:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.29" />
                    <SPLIT distance="100" swimtime="00:01:17.96" />
                    <SPLIT distance="150" swimtime="00:02:01.63" />
                    <SPLIT distance="200" swimtime="00:02:46.82" />
                    <SPLIT distance="250" swimtime="00:03:32.53" />
                    <SPLIT distance="300" swimtime="00:04:18.75" />
                    <SPLIT distance="350" swimtime="00:05:06.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-04-20" firstname="Anna" gender="F" lastname="Kičínová" nation="SVK" license="SVK13974" athleteid="14685">
              <RESULTS>
                <RESULT eventid="1096" points="229" reactiontime="+98" swimtime="00:03:19.15" resultid="14686" heatid="19306" lane="6" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.62" />
                    <SPLIT distance="100" swimtime="00:01:38.86" />
                    <SPLIT distance="150" swimtime="00:02:32.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="270" reactiontime="+91" swimtime="00:03:28.02" resultid="14687" heatid="19357" lane="6" entrytime="00:03:24.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.93" />
                    <SPLIT distance="100" swimtime="00:01:41.94" />
                    <SPLIT distance="150" swimtime="00:02:35.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="224" reactiontime="+99" swimtime="00:03:16.76" resultid="14688" heatid="19412" lane="2" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.94" />
                    <SPLIT distance="100" swimtime="00:01:32.28" />
                    <SPLIT distance="150" swimtime="00:02:24.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="269" reactiontime="+76" swimtime="00:01:36.52" resultid="14689" heatid="19430" lane="7" entrytime="00:01:34.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="197" reactiontime="+90" swimtime="00:00:41.85" resultid="14690" heatid="19446" lane="4" entrytime="00:00:38.20" />
                <RESULT eventid="1595" points="232" swimtime="00:01:28.82" resultid="14691" heatid="19514" lane="6" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="260" reactiontime="+96" swimtime="00:00:44.83" resultid="14692" heatid="19542" lane="0" entrytime="00:00:43.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-04-12" firstname="Zuzana" gender="F" lastname="Matúšová" nation="SVK" license="SVK21695" athleteid="14712">
              <RESULTS>
                <RESULT eventid="1062" points="502" reactiontime="+80" swimtime="00:00:29.24" resultid="14713" heatid="19282" lane="5" entrytime="00:00:29.80" />
                <RESULT eventid="1096" points="421" reactiontime="+88" swimtime="00:02:42.58" resultid="14714" heatid="19308" lane="5" entrytime="00:02:46.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                    <SPLIT distance="100" swimtime="00:01:18.02" />
                    <SPLIT distance="150" swimtime="00:02:05.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="347" reactiontime="+83" swimtime="00:00:36.50" resultid="14715" heatid="19340" lane="0" entrytime="00:00:36.80" />
                <RESULT eventid="14225" points="464" reactiontime="+77" swimtime="00:01:13.19" resultid="14716" heatid="19395" lane="8" entrytime="00:01:14.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="456" reactiontime="+84" swimtime="00:00:31.67" resultid="14717" heatid="19449" lane="1" entrytime="00:00:31.10" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" points="348" reactiontime="+86" swimtime="00:02:05.88" resultid="14718" heatid="19321" lane="1" entrytime="00:02:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                    <SPLIT distance="100" swimtime="00:01:12.62" />
                    <SPLIT distance="150" swimtime="00:01:38.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14699" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="14685" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="14712" number="3" />
                    <RELAYPOSITION athleteid="14693" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" points="340" reactiontime="+70" swimtime="00:02:19.18" resultid="14719" heatid="19563" lane="8" entrytime="00:02:20.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.93" />
                    <SPLIT distance="100" swimtime="00:01:17.06" />
                    <SPLIT distance="150" swimtime="00:01:48.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14693" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="14685" number="2" reactiontime="+33" />
                    <RELAYPOSITION athleteid="14712" number="3" reactiontime="+60" />
                    <RELAYPOSITION athleteid="14699" number="4" reactiontime="+64" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>

<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="SiKReT Gliwice" version="11.59270">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Gliwice" name="Letnie Mistrzostwa Polski w Pływaniu Masters" course="LCM" hostclub="SiKReT Gliwice" hostclub.url="http://www.sikret-plywanie.pl" organizer="Samorząd Miasta Gliwice, MZUK Gliwice, PZP,SLOZP,SiKReT Gliwice" reservecount="2" result.url="http://www.megatiming.pl" startmethod="1" timing="AUTOMATIC" nation="POL">
      <AGEDATE value="2019-05-31" type="YEAR" />
      <POOL name="Olimpijczyk Gliwice" lanemax="9" />
      <FACILITY city="Gliwice" name="Olimpijczyk Gliwice" nation="POL" />
      <POINTTABLE pointtableid="3012" name="FINA Point Scoring" version="2019" />
      <CONTACT email="wisniowicz@gmail.com" name="Wojciech Wiśniowicz" phone="500193225" />
      <SESSIONS>
        <SESSION date="2019-05-31" daytime="15:00" endtime="21:41" name="BLOK I" number="1" warmupfrom="13:30">
          <EVENTS>
            <EVENT eventid="19751" daytime="18:35" gender="F" number="8" order="11" round="FHT" preveventid="1165">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="24319" daytime="18:35" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="19749" daytime="16:30" gender="F" number="6" order="7" round="FHT" preveventid="1147">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="24312" daytime="16:30" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="14207" daytime="20:00" gender="M" number="9" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="24531" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19952" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24532" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22048" />
                    <RANKING order="2" place="2" resultid="20186" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24533" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19846" />
                    <RANKING order="2" place="2" resultid="21502" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24534" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="19781" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24535" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22069" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24536" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20414" />
                    <RANKING order="2" place="2" resultid="21400" />
                    <RANKING order="3" place="3" resultid="21591" />
                    <RANKING order="4" place="4" resultid="21218" />
                    <RANKING order="5" place="5" resultid="21827" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24537" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="20252" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24538" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22063" />
                    <RANKING order="2" place="2" resultid="20401" />
                    <RANKING order="3" place="-1" resultid="19802" />
                    <RANKING order="4" place="-1" resultid="22268" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24539" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21528" />
                    <RANKING order="2" place="2" resultid="22677" />
                    <RANKING order="3" place="3" resultid="21835" />
                    <RANKING order="4" place="4" resultid="22305" />
                    <RANKING order="5" place="5" resultid="21522" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24540" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20141" />
                    <RANKING order="2" place="2" resultid="20960" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24541" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="20159" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24542" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="21370" />
                    <RANKING order="2" place="-1" resultid="20938" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24543" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22647" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24544" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21494" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24545" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="24546" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24320" daytime="20:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24321" daytime="20:45" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="14189" daytime="17:30" gender="M" number="7" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="24499" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22318" />
                    <RANKING order="2" place="-1" resultid="21425" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24500" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21280" />
                    <RANKING order="2" place="-1" resultid="21095" />
                    <RANKING order="3" place="-1" resultid="21930" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24501" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21722" />
                    <RANKING order="2" place="2" resultid="20498" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24502" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22356" />
                    <RANKING order="2" place="2" resultid="20624" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24503" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20682" />
                    <RANKING order="2" place="2" resultid="19763" />
                    <RANKING order="3" place="3" resultid="20194" />
                    <RANKING order="4" place="4" resultid="21857" />
                    <RANKING order="5" place="-1" resultid="22488" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24504" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22031" />
                    <RANKING order="2" place="2" resultid="20285" />
                    <RANKING order="3" place="3" resultid="21871" />
                    <RANKING order="4" place="4" resultid="22039" />
                    <RANKING order="5" place="5" resultid="19973" />
                    <RANKING order="6" place="6" resultid="21476" />
                    <RANKING order="7" place="-1" resultid="22250" />
                    <RANKING order="8" place="-1" resultid="23367" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24505" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21980" />
                    <RANKING order="2" place="2" resultid="21352" />
                    <RANKING order="3" place="3" resultid="20931" />
                    <RANKING order="4" place="4" resultid="19982" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24506" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20917" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24507" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21120" />
                    <RANKING order="2" place="2" resultid="20692" />
                    <RANKING order="3" place="3" resultid="21468" />
                    <RANKING order="4" place="4" resultid="22394" />
                    <RANKING order="5" place="-1" resultid="20454" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24508" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20491" />
                    <RANKING order="2" place="2" resultid="23428" />
                    <RANKING order="3" place="3" resultid="19946" />
                    <RANKING order="4" place="-1" resultid="19773" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24509" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21325" />
                    <RANKING order="2" place="2" resultid="20385" />
                    <RANKING order="3" place="-1" resultid="20514" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24510" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22624" />
                    <RANKING order="2" place="2" resultid="19937" />
                    <RANKING order="3" place="3" resultid="22424" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24511" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="24512" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="24513" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="24514" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24313" daytime="17:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24314" daytime="17:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24315" daytime="18:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24316" daytime="18:25" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="19752" daytime="19:40" gender="M" number="9" order="13" round="FHT" preveventid="14207">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="24322" daytime="19:40" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1062" daytime="15:00" gender="F" number="1" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1064" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21288" />
                    <RANKING order="2" place="2" resultid="20780" />
                    <RANKING order="3" place="3" resultid="22663" />
                    <RANKING order="4" place="4" resultid="20767" />
                    <RANKING order="5" place="5" resultid="20750" />
                    <RANKING order="6" place="6" resultid="21441" />
                    <RANKING order="7" place="7" resultid="22917" />
                    <RANKING order="8" place="8" resultid="21197" />
                    <RANKING order="9" place="9" resultid="20764" />
                    <RANKING order="10" place="10" resultid="21952" />
                    <RANKING order="11" place="-1" resultid="23391" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21261" />
                    <RANKING order="2" place="2" resultid="21551" />
                    <RANKING order="3" place="3" resultid="23419" />
                    <RANKING order="4" place="4" resultid="21900" />
                    <RANKING order="5" place="5" resultid="21187" />
                    <RANKING order="6" place="6" resultid="22637" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22986" />
                    <RANKING order="2" place="2" resultid="20734" />
                    <RANKING order="3" place="3" resultid="21936" />
                    <RANKING order="4" place="4" resultid="22456" />
                    <RANKING order="5" place="5" resultid="21388" />
                    <RANKING order="6" place="6" resultid="20638" />
                    <RANKING order="7" place="7" resultid="21909" />
                    <RANKING order="8" place="8" resultid="21906" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20955" />
                    <RANKING order="2" place="2" resultid="22923" />
                    <RANKING order="3" place="3" resultid="22882" />
                    <RANKING order="4" place="4" resultid="20741" />
                    <RANKING order="5" place="-1" resultid="20165" />
                    <RANKING order="6" place="-1" resultid="21761" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1068" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21176" />
                    <RANKING order="2" place="1" resultid="22951" />
                    <RANKING order="3" place="3" resultid="23059" />
                    <RANKING order="4" place="4" resultid="21820" />
                    <RANKING order="5" place="5" resultid="22024" />
                    <RANKING order="6" place="6" resultid="21895" />
                    <RANKING order="7" place="-1" resultid="19906" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21171" />
                    <RANKING order="2" place="2" resultid="21747" />
                    <RANKING order="3" place="3" resultid="20215" />
                    <RANKING order="4" place="4" resultid="21839" />
                    <RANKING order="5" place="5" resultid="23351" />
                    <RANKING order="6" place="6" resultid="21360" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21297" />
                    <RANKING order="2" place="2" resultid="22888" />
                    <RANKING order="3" place="3" resultid="20202" />
                    <RANKING order="4" place="4" resultid="22900" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21112" />
                    <RANKING order="2" place="2" resultid="21315" />
                    <RANKING order="3" place="3" resultid="20445" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1072" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21376" />
                    <RANKING order="2" place="2" resultid="22282" />
                    <RANKING order="3" place="3" resultid="21605" />
                    <RANKING order="4" place="4" resultid="21614" />
                    <RANKING order="5" place="5" resultid="20481" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1073" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19868" />
                    <RANKING order="2" place="2" resultid="21484" />
                    <RANKING order="3" place="3" resultid="22275" />
                    <RANKING order="4" place="4" resultid="21629" />
                    <RANKING order="5" place="5" resultid="22691" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1074" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21228" />
                    <RANKING order="2" place="2" resultid="20116" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1075" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19882" />
                    <RANKING order="2" place="2" resultid="21224" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1076" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1077" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1078" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1063" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24275" daytime="15:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24276" daytime="15:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24277" daytime="15:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24278" daytime="15:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="24279" daytime="15:05" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="24280" daytime="15:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="24281" daytime="15:10" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1130" daytime="16:25" gender="X" number="5" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="12486" agemax="99" agemin="80" calculate="TOTAL" />
                <AGEGROUP agegroupid="1182" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21564" />
                    <RANKING order="2" place="2" resultid="22094" />
                    <RANKING order="3" place="-1" resultid="21959" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1183" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21958" />
                    <RANKING order="2" place="2" resultid="20655" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1184" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22088" />
                    <RANKING order="2" place="2" resultid="21891" />
                    <RANKING order="3" place="3" resultid="22511" />
                    <RANKING order="4" place="4" resultid="22983" />
                    <RANKING order="5" place="5" resultid="21212" />
                    <RANKING order="6" place="6" resultid="23377" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1185" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21214" />
                    <RANKING order="2" place="2" resultid="22371" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1186" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21395" />
                    <RANKING order="2" place="2" resultid="21640" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1145" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19921" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24308" daytime="16:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24309" daytime="16:25" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1147" daytime="16:45" gender="F" number="6" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="24483" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22296" />
                    <RANKING order="2" place="2" resultid="20751" />
                    <RANKING order="3" place="-1" resultid="22918" />
                    <RANKING order="4" place="-1" resultid="20759" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24484" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22056" />
                    <RANKING order="2" place="2" resultid="22018" />
                    <RANKING order="3" place="3" resultid="21201" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24485" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21389" />
                    <RANKING order="2" place="2" resultid="22010" />
                    <RANKING order="3" place="-1" resultid="21739" />
                    <RANKING order="4" place="-1" resultid="20639" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24486" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22494" />
                    <RANKING order="2" place="2" resultid="20739" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24487" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20258" />
                    <RANKING order="2" place="2" resultid="21409" />
                    <RANKING order="3" place="3" resultid="20898" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24488" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19899" />
                    <RANKING order="2" place="2" resultid="21748" />
                    <RANKING order="3" place="3" resultid="20216" />
                    <RANKING order="4" place="4" resultid="21684" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24489" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22287" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24490" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21316" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24491" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21606" />
                    <RANKING order="2" place="2" resultid="21615" />
                    <RANKING order="3" place="3" resultid="20716" />
                    <RANKING order="4" place="4" resultid="20482" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24492" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22692" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24493" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="24494" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19892" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24495" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="24496" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="24497" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="24498" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24310" daytime="16:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24311" daytime="17:05" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="19750" daytime="17:20" gender="M" number="7" order="9" round="FHT" preveventid="14189">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="24317" daytime="17:20" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1113" daytime="15:45" gender="M" number="4" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1114" agemax="24" agemin="20" />
                <AGEGROUP agegroupid="1115" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22047" />
                    <RANKING order="2" place="2" resultid="21279" />
                    <RANKING order="3" place="3" resultid="22967" />
                    <RANKING order="4" place="4" resultid="21884" />
                    <RANKING order="5" place="5" resultid="21094" />
                    <RANKING order="6" place="6" resultid="21929" />
                    <RANKING order="7" place="7" resultid="22680" />
                    <RANKING order="8" place="8" resultid="20946" />
                    <RANKING order="9" place="9" resultid="21508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1116" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21721" />
                    <RANKING order="2" place="2" resultid="21249" />
                    <RANKING order="3" place="3" resultid="22995" />
                    <RANKING order="4" place="4" resultid="22262" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1117" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="23004" />
                    <RANKING order="2" place="2" resultid="22330" />
                    <RANKING order="3" place="-1" resultid="20505" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1118" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20681" />
                    <RANKING order="2" place="2" resultid="22339" />
                    <RANKING order="3" place="3" resultid="22932" />
                    <RANKING order="4" place="4" resultid="21578" />
                    <RANKING order="5" place="5" resultid="19762" />
                    <RANKING order="6" place="6" resultid="21165" />
                    <RANKING order="7" place="7" resultid="21450" />
                    <RANKING order="8" place="8" resultid="22472" />
                    <RANKING order="9" place="9" resultid="22389" />
                    <RANKING order="10" place="10" resultid="19768" />
                    <RANKING order="11" place="-1" resultid="22322" />
                    <RANKING order="12" place="-1" resultid="23417" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1119" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20172" />
                    <RANKING order="2" place="2" resultid="20726" />
                    <RANKING order="3" place="3" resultid="21415" />
                    <RANKING order="4" place="4" resultid="19965" />
                    <RANKING order="5" place="5" resultid="21870" />
                    <RANKING order="6" place="6" resultid="20289" />
                    <RANKING order="7" place="7" resultid="22401" />
                    <RANKING order="8" place="-1" resultid="21878" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1120" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22876" />
                    <RANKING order="2" place="2" resultid="20909" />
                    <RANKING order="3" place="3" resultid="19815" />
                    <RANKING order="4" place="4" resultid="20225" />
                    <RANKING order="5" place="5" resultid="22894" />
                    <RANKING order="6" place="-1" resultid="21233" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1121" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21256" />
                    <RANKING order="2" place="2" resultid="20276" />
                    <RANKING order="3" place="3" resultid="20179" />
                    <RANKING order="4" place="4" resultid="20469" />
                    <RANKING order="5" place="5" resultid="22313" />
                    <RANKING order="6" place="-1" resultid="21343" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1122" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21150" />
                    <RANKING order="2" place="2" resultid="21467" />
                    <RANKING order="3" place="3" resultid="22445" />
                    <RANKING order="4" place="4" resultid="22304" />
                    <RANKING order="5" place="5" resultid="20453" />
                    <RANKING order="6" place="6" resultid="20461" />
                    <RANKING order="7" place="-1" resultid="21119" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1123" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21843" />
                    <RANKING order="2" place="2" resultid="22432" />
                    <RANKING order="3" place="3" resultid="20421" />
                    <RANKING order="4" place="4" resultid="20140" />
                    <RANKING order="5" place="5" resultid="21971" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1124" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21134" />
                    <RANKING order="2" place="2" resultid="19930" />
                    <RANKING order="3" place="3" resultid="21324" />
                    <RANKING order="4" place="4" resultid="20384" />
                    <RANKING order="5" place="5" resultid="20132" />
                    <RANKING order="6" place="6" resultid="20513" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1125" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21459" />
                    <RANKING order="2" place="2" resultid="19936" />
                    <RANKING order="3" place="3" resultid="20937" />
                    <RANKING order="4" place="-1" resultid="20149" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1126" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22650" />
                    <RANKING order="2" place="2" resultid="20889" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1127" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20700" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1128" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1129" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24300" daytime="15:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24301" daytime="15:55" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24302" daytime="16:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24303" daytime="16:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="24304" daytime="16:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="24305" daytime="16:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="24306" daytime="16:15" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="24307" daytime="16:20" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1096" daytime="15:35" gender="F" number="3" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1097" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21289" />
                    <RANKING order="2" place="2" resultid="22295" />
                    <RANKING order="3" place="3" resultid="21442" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20775" />
                    <RANKING order="2" place="2" resultid="21262" />
                    <RANKING order="3" place="3" resultid="23420" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1099" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22009" />
                    <RANKING order="2" place="2" resultid="22499" />
                    <RANKING order="3" place="3" resultid="21738" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1100" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20645" />
                    <RANKING order="2" place="-1" resultid="21762" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1101" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21408" />
                    <RANKING order="2" place="2" resultid="21144" />
                    <RANKING order="3" place="3" resultid="22256" />
                    <RANKING order="4" place="4" resultid="21534" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21128" />
                    <RANKING order="2" place="2" resultid="21730" />
                    <RANKING order="3" place="3" resultid="21683" />
                    <RANKING order="4" place="4" resultid="21361" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1103" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20203" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1104" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21333" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1105" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21515" />
                    <RANKING order="2" place="2" resultid="22632" />
                    <RANKING order="3" place="3" resultid="21377" />
                    <RANKING order="4" place="4" resultid="20707" />
                    <RANKING order="5" place="-1" resultid="20715" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1106" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1107" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1108" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19883" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1109" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1110" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1111" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1112" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24297" daytime="15:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24298" daytime="15:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24299" daytime="15:45" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1079" daytime="15:10" gender="M" number="2" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1080" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21427" />
                    <RANKING order="2" place="2" resultid="23397" />
                    <RANKING order="3" place="3" resultid="20307" />
                    <RANKING order="4" place="4" resultid="22962" />
                    <RANKING order="5" place="5" resultid="23379" />
                    <RANKING order="6" place="6" resultid="21436" />
                    <RANKING order="7" place="7" resultid="20968" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1081" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22667" />
                    <RANKING order="2" place="2" resultid="22441" />
                    <RANKING order="3" place="3" resultid="21541" />
                    <RANKING order="4" place="4" resultid="21883" />
                    <RANKING order="5" place="5" resultid="21662" />
                    <RANKING order="6" place="6" resultid="22973" />
                    <RANKING order="7" place="7" resultid="20302" />
                    <RANKING order="8" place="8" resultid="20773" />
                    <RANKING order="9" place="9" resultid="21507" />
                    <RANKING order="10" place="10" resultid="23357" />
                    <RANKING order="11" place="11" resultid="21940" />
                    <RANKING order="12" place="12" resultid="22679" />
                    <RANKING order="13" place="13" resultid="22658" />
                    <RANKING order="14" place="14" resultid="21944" />
                    <RANKING order="15" place="15" resultid="20631" />
                    <RANKING order="16" place="16" resultid="22642" />
                    <RANKING order="17" place="-1" resultid="21948" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1082" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21702" />
                    <RANKING order="2" place="2" resultid="21248" />
                    <RANKING order="3" place="3" resultid="21919" />
                    <RANKING order="4" place="4" resultid="22994" />
                    <RANKING order="5" place="5" resultid="22461" />
                    <RANKING order="6" place="6" resultid="21692" />
                    <RANKING order="7" place="7" resultid="22244" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1083" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22505" />
                    <RANKING order="2" place="2" resultid="22329" />
                    <RANKING order="3" place="3" resultid="23003" />
                    <RANKING order="4" place="4" resultid="20233" />
                    <RANKING order="5" place="5" resultid="19757" />
                    <RANKING order="6" place="6" resultid="22083" />
                    <RANKING order="7" place="7" resultid="21695" />
                    <RANKING order="8" place="8" resultid="22355" />
                    <RANKING order="9" place="9" resultid="19780" />
                    <RANKING order="10" place="10" resultid="20623" />
                    <RANKING order="11" place="11" resultid="20653" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1084" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22931" />
                    <RANKING order="2" place="2" resultid="22616" />
                    <RANKING order="3" place="3" resultid="22936" />
                    <RANKING order="4" place="4" resultid="22338" />
                    <RANKING order="5" place="5" resultid="21164" />
                    <RANKING order="6" place="6" resultid="22945" />
                    <RANKING order="7" place="7" resultid="22321" />
                    <RANKING order="8" place="8" resultid="22068" />
                    <RANKING order="9" place="9" resultid="22471" />
                    <RANKING order="10" place="10" resultid="21449" />
                    <RANKING order="11" place="11" resultid="22941" />
                    <RANKING order="12" place="12" resultid="21678" />
                    <RANKING order="13" place="13" resultid="21856" />
                    <RANKING order="14" place="14" resultid="20950" />
                    <RANKING order="15" place="15" resultid="21848" />
                    <RANKING order="16" place="16" resultid="20193" />
                    <RANKING order="17" place="17" resultid="20109" />
                    <RANKING order="18" place="18" resultid="22378" />
                    <RANKING order="19" place="19" resultid="21599" />
                    <RANKING order="20" place="20" resultid="22388" />
                    <RANKING order="21" place="21" resultid="21393" />
                    <RANKING order="22" place="-1" resultid="22487" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1085" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20171" />
                    <RANKING order="2" place="2" resultid="22030" />
                    <RANKING order="3" place="3" resultid="20725" />
                    <RANKING order="4" place="4" resultid="19964" />
                    <RANKING order="5" place="5" resultid="22956" />
                    <RANKING order="6" place="6" resultid="21475" />
                    <RANKING order="7" place="7" resultid="21877" />
                    <RANKING order="8" place="8" resultid="23091" />
                    <RANKING order="9" place="9" resultid="21590" />
                    <RANKING order="10" place="10" resultid="20284" />
                    <RANKING order="11" place="11" resultid="21826" />
                    <RANKING order="12" place="12" resultid="21421" />
                    <RANKING order="13" place="13" resultid="21399" />
                    <RANKING order="14" place="14" resultid="19972" />
                    <RANKING order="15" place="15" resultid="22400" />
                    <RANKING order="16" place="16" resultid="23366" />
                    <RANKING order="17" place="17" resultid="21182" />
                    <RANKING order="18" place="18" resultid="22038" />
                    <RANKING order="19" place="-1" resultid="20267" />
                    <RANKING order="20" place="-1" resultid="21217" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1086" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21099" />
                    <RANKING order="2" place="2" resultid="22875" />
                    <RANKING order="3" place="3" resultid="20908" />
                    <RANKING order="4" place="4" resultid="21572" />
                    <RANKING order="5" place="5" resultid="21979" />
                    <RANKING order="6" place="6" resultid="21192" />
                    <RANKING order="7" place="7" resultid="21351" />
                    <RANKING order="8" place="8" resultid="21139" />
                    <RANKING order="9" place="9" resultid="19810" />
                    <RANKING order="10" place="10" resultid="19981" />
                    <RANKING order="11" place="11" resultid="20923" />
                    <RANKING order="12" place="12" resultid="21671" />
                    <RANKING order="13" place="13" resultid="20224" />
                    <RANKING order="14" place="14" resultid="22893" />
                    <RANKING order="15" place="-1" resultid="20930" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1087" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22466" />
                    <RANKING order="2" place="2" resultid="21255" />
                    <RANKING order="3" place="3" resultid="20275" />
                    <RANKING order="4" place="4" resultid="20468" />
                    <RANKING order="5" place="5" resultid="21342" />
                    <RANKING order="6" place="6" resultid="20400" />
                    <RANKING order="7" place="-1" resultid="19801" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1088" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22002" />
                    <RANKING order="2" place="2" resultid="19858" />
                    <RANKING order="3" place="3" resultid="21264" />
                    <RANKING order="4" place="4" resultid="21149" />
                    <RANKING order="5" place="5" resultid="21622" />
                    <RANKING order="6" place="6" resultid="20691" />
                    <RANKING order="7" place="7" resultid="21240" />
                    <RANKING order="8" place="8" resultid="22393" />
                    <RANKING order="9" place="9" resultid="19795" />
                    <RANKING order="10" place="10" resultid="20460" />
                    <RANKING order="11" place="-1" resultid="22676" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1089" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22451" />
                    <RANKING order="2" place="2" resultid="19772" />
                    <RANKING order="3" place="3" resultid="20490" />
                    <RANKING order="4" place="4" resultid="21970" />
                    <RANKING order="5" place="5" resultid="23427" />
                    <RANKING order="6" place="6" resultid="20883" />
                    <RANKING order="7" place="7" resultid="19945" />
                    <RANKING order="8" place="-1" resultid="20959" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1090" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19874" />
                    <RANKING order="2" place="2" resultid="21133" />
                    <RANKING order="3" place="3" resultid="19929" />
                    <RANKING order="4" place="4" resultid="20158" />
                    <RANKING order="5" place="5" resultid="19916" />
                    <RANKING order="6" place="6" resultid="20131" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1091" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21636" />
                    <RANKING order="2" place="2" resultid="21458" />
                    <RANKING order="3" place="3" resultid="22423" />
                    <RANKING order="4" place="4" resultid="21369" />
                    <RANKING order="5" place="5" resultid="20437" />
                    <RANKING order="6" place="-1" resultid="22623" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1092" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22649" />
                    <RANKING order="2" place="2" resultid="20888" />
                    <RANKING order="3" place="3" resultid="21988" />
                    <RANKING order="4" place="4" resultid="22415" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1093" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20699" />
                    <RANKING order="2" place="2" resultid="21493" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1095" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24282" daytime="15:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24283" daytime="15:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24284" daytime="15:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24285" daytime="15:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="24286" daytime="15:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="24287" daytime="15:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="24288" daytime="15:20" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="24289" daytime="15:25" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="24290" daytime="15:25" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="24291" daytime="15:25" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="24292" daytime="15:25" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="24293" daytime="15:30" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="24294" daytime="15:30" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="24295" daytime="15:30" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="24296" daytime="15:30" number="15" order="15" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1165" daytime="19:05" gender="F" number="8" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="24515" agemax="24" agemin="20" />
                <AGEGROUP agegroupid="24516" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21585" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24517" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22500" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24518" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="22948" />
                    <RANKING order="2" place="-1" resultid="22911" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24519" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="24520" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="23363" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24521" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20394" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24522" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21862" />
                    <RANKING order="2" place="-1" resultid="21334" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24523" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21516" />
                    <RANKING order="2" place="-1" resultid="20708" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24524" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="24525" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22438" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24526" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="24527" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="24528" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="24529" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="24530" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24318" daytime="19:05" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2019-06-01" daytime="09:00" endtime="12:24" name="BLOK II" number="2" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="1187" daytime="09:00" gender="F" number="10" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1189" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21290" />
                    <RANKING order="2" place="2" resultid="21556" />
                    <RANKING order="3" place="3" resultid="21198" />
                    <RANKING order="4" place="4" resultid="23392" />
                    <RANKING order="5" place="5" resultid="22919" />
                    <RANKING order="6" place="6" resultid="20752" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1190" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21552" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1191" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21925" />
                    <RANKING order="2" place="2" resultid="22011" />
                    <RANKING order="3" place="3" resultid="21910" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1192" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20646" />
                    <RANKING order="2" place="2" resultid="22883" />
                    <RANKING order="3" place="-1" resultid="20166" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1193" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22025" />
                    <RANKING order="2" place="2" resultid="21177" />
                    <RANKING order="3" place="3" resultid="22257" />
                    <RANKING order="4" place="4" resultid="22952" />
                    <RANKING order="5" place="5" resultid="21821" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1194" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21172" />
                    <RANKING order="2" place="2" resultid="21749" />
                    <RANKING order="3" place="3" resultid="21731" />
                    <RANKING order="4" place="4" resultid="20217" />
                    <RANKING order="5" place="5" resultid="23352" />
                    <RANKING order="6" place="6" resultid="21362" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1195" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21298" />
                    <RANKING order="2" place="2" resultid="22889" />
                    <RANKING order="3" place="3" resultid="22288" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1196" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21113" />
                    <RANKING order="2" place="2" resultid="21863" />
                    <RANKING order="3" place="3" resultid="21335" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1197" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21607" />
                    <RANKING order="2" place="2" resultid="19909" />
                    <RANKING order="3" place="3" resultid="20717" />
                    <RANKING order="4" place="4" resultid="20483" />
                    <RANKING order="5" place="5" resultid="22906" />
                    <RANKING order="6" place="6" resultid="19865" />
                    <RANKING order="7" place="7" resultid="23856" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1198" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19869" />
                    <RANKING order="2" place="2" resultid="21485" />
                    <RANKING order="3" place="3" resultid="21630" />
                    <RANKING order="4" place="4" resultid="19838" />
                    <RANKING order="5" place="5" resultid="19853" />
                    <RANKING order="6" place="6" resultid="22693" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1199" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20117" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1200" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19884" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1201" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20427" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1202" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1203" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1204" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24323" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24324" daytime="09:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24325" daytime="09:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24326" daytime="09:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="24327" daytime="09:05" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1324" daytime="11:00" gender="F" number="16" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1325" agemax="24" agemin="20" />
                <AGEGROUP agegroupid="1326" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22057" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1327" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22012" />
                    <RANKING order="2" place="2" resultid="21741" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1328" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="1329" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21145" />
                    <RANKING order="2" place="2" resultid="21536" />
                    <RANKING order="3" place="3" resultid="21273" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1330" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21129" />
                    <RANKING order="2" place="2" resultid="21732" />
                    <RANKING order="3" place="3" resultid="21363" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1331" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="1332" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21318" />
                    <RANKING order="2" place="2" resultid="21336" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1333" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21379" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1334" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1335" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1336" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1337" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1338" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1339" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1340" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24366" daytime="11:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24367" daytime="11:05" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1222" daytime="09:25" gender="F" number="12" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1223" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22297" />
                    <RANKING order="2" place="2" resultid="23066" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1224" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20776" />
                    <RANKING order="2" place="2" resultid="21202" />
                    <RANKING order="3" place="3" resultid="22638" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1225" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22987" />
                    <RANKING order="2" place="2" resultid="21740" />
                    <RANKING order="3" place="3" resultid="21994" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1226" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20748" />
                    <RANKING order="2" place="2" resultid="22912" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1227" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20245" />
                    <RANKING order="2" place="2" resultid="19789" />
                    <RANKING order="3" place="3" resultid="21754" />
                    <RANKING order="4" place="4" resultid="21272" />
                    <RANKING order="5" place="5" resultid="21535" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1228" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19900" />
                    <RANKING order="2" place="2" resultid="21685" />
                    <RANKING order="3" place="3" resultid="24067" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1229" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20204" />
                    <RANKING order="2" place="2" resultid="22901" />
                    <RANKING order="3" place="3" resultid="23081" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1230" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22482" />
                    <RANKING order="2" place="2" resultid="23371" />
                    <RANKING order="3" place="3" resultid="21864" />
                    <RANKING order="4" place="-1" resultid="23404" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1231" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22283" />
                    <RANKING order="2" place="2" resultid="21616" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1232" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22276" />
                    <RANKING order="2" place="2" resultid="20448" />
                    <RANKING order="3" place="3" resultid="19854" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1233" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21229" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1234" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19893" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1235" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20428" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1236" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1237" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1238" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24337" daytime="09:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24338" daytime="09:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24339" daytime="09:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24340" daytime="09:40" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1341" daytime="11:10" gender="M" number="17" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1342" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22963" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1343" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21282" />
                    <RANKING order="2" place="2" resultid="20432" />
                    <RANKING order="3" place="3" resultid="22050" />
                    <RANKING order="4" place="4" resultid="20187" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1344" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21724" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1345" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="23006" />
                    <RANKING order="2" place="2" resultid="22357" />
                    <RANKING order="3" place="-1" resultid="22077" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1346" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20684" />
                    <RANKING order="2" place="2" resultid="19764" />
                    <RANKING order="3" place="-1" resultid="21579" />
                    <RANKING order="4" place="-1" resultid="22937" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1347" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21872" />
                    <RANKING order="2" place="2" resultid="20290" />
                    <RANKING order="3" place="3" resultid="21402" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1348" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21982" />
                    <RANKING order="2" place="2" resultid="20925" />
                    <RANKING order="3" place="3" resultid="20254" />
                    <RANKING order="4" place="4" resultid="19816" />
                    <RANKING order="5" place="5" resultid="20227" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1349" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20180" />
                    <RANKING order="2" place="2" resultid="22269" />
                    <RANKING order="3" place="3" resultid="20918" />
                    <RANKING order="4" place="-1" resultid="19804" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1350" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22003" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1351" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21973" />
                    <RANKING order="2" place="2" resultid="20143" />
                    <RANKING order="3" place="3" resultid="23430" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1352" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22673" />
                    <RANKING order="2" place="2" resultid="21327" />
                    <RANKING order="3" place="3" resultid="20387" />
                    <RANKING order="4" place="4" resultid="20516" />
                    <RANKING order="5" place="-1" resultid="20134" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1353" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19939" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1354" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1355" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1356" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1357" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24368" daytime="11:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24369" daytime="11:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24370" daytime="11:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24371" daytime="11:25" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1239" daytime="09:45" gender="M" number="13" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1240" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19953" />
                    <RANKING order="2" place="2" resultid="21426" />
                    <RANKING order="3" place="3" resultid="20969" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1241" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21885" />
                    <RANKING order="2" place="2" resultid="23075" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1242" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21703" />
                    <RANKING order="2" place="2" resultid="21723" />
                    <RANKING order="3" place="3" resultid="20499" />
                    <RANKING order="4" place="4" resultid="22245" />
                    <RANKING order="5" place="5" resultid="22263" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1243" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22331" />
                    <RANKING order="2" place="2" resultid="22084" />
                    <RANKING order="3" place="-1" resultid="22076" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1244" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20683" />
                    <RANKING order="2" place="2" resultid="21166" />
                    <RANKING order="3" place="3" resultid="23413" />
                    <RANKING order="4" place="4" resultid="22473" />
                    <RANKING order="5" place="5" resultid="21849" />
                    <RANKING order="6" place="6" resultid="20196" />
                    <RANKING order="7" place="7" resultid="22390" />
                    <RANKING order="8" place="8" resultid="23415" />
                    <RANKING order="9" place="-1" resultid="21452" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1245" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20901" />
                    <RANKING order="2" place="2" resultid="21416" />
                    <RANKING order="3" place="3" resultid="19974" />
                    <RANKING order="4" place="4" resultid="21305" />
                    <RANKING order="5" place="5" resultid="22402" />
                    <RANKING order="6" place="-1" resultid="20268" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1246" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21573" />
                    <RANKING order="2" place="2" resultid="21235" />
                    <RANKING order="3" place="3" resultid="21354" />
                    <RANKING order="4" place="4" resultid="20924" />
                    <RANKING order="5" place="5" resultid="20253" />
                    <RANKING order="6" place="6" resultid="22382" />
                    <RANKING order="7" place="-1" resultid="22896" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1247" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22314" />
                    <RANKING order="2" place="2" resultid="21345" />
                    <RANKING order="3" place="-1" resultid="19803" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1248" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21998" />
                    <RANKING order="2" place="2" resultid="21152" />
                    <RANKING order="3" place="3" resultid="22446" />
                    <RANKING order="4" place="4" resultid="23410" />
                    <RANKING order="5" place="5" resultid="19797" />
                    <RANKING order="6" place="6" resultid="22307" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1249" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22433" />
                    <RANKING order="2" place="2" resultid="20884" />
                    <RANKING order="3" place="3" resultid="20422" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1250" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21106" />
                    <RANKING order="2" place="2" resultid="20386" />
                    <RANKING order="3" place="3" resultid="20133" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1251" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19888" />
                    <RANKING order="2" place="2" resultid="19938" />
                    <RANKING order="3" place="3" resultid="20940" />
                    <RANKING order="4" place="4" resultid="20439" />
                    <RANKING order="5" place="-1" resultid="20151" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1252" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20891" />
                    <RANKING order="2" place="2" resultid="22417" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1253" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21495" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1254" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1255" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24341" daytime="09:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24342" daytime="09:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24343" daytime="10:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24344" daytime="10:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="24345" daytime="10:05" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="24346" daytime="10:10" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1381" daytime="11:35" gender="M" number="19" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="16653" agemax="99" agemin="80" calculate="TOTAL" />
                <AGEGROUP agegroupid="16654" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21964" />
                    <RANKING order="2" place="2" resultid="22687" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16655" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22510" />
                    <RANKING order="2" place="2" resultid="22095" />
                    <RANKING order="3" place="3" resultid="22982" />
                    <RANKING order="4" place="-1" resultid="22512" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16656" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22367" />
                    <RANKING order="2" place="2" resultid="22981" />
                    <RANKING order="3" place="3" resultid="21422" />
                    <RANKING order="4" place="4" resultid="21716" />
                    <RANKING order="5" place="-1" resultid="21892" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16657" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="21206" />
                    <RANKING order="2" place="-1" resultid="22368" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16658" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21208" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16659" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19923" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24373" daytime="11:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24374" daytime="11:40" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1256" daytime="10:15" gender="F" number="14" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1257" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21291" />
                    <RANKING order="2" place="2" resultid="22664" />
                    <RANKING order="3" place="3" resultid="20753" />
                    <RANKING order="4" place="4" resultid="20768" />
                    <RANKING order="5" place="5" resultid="20744" />
                    <RANKING order="6" place="6" resultid="22298" />
                    <RANKING order="7" place="7" resultid="21443" />
                    <RANKING order="8" place="8" resultid="23393" />
                    <RANKING order="9" place="9" resultid="23067" />
                    <RANKING order="10" place="10" resultid="20760" />
                    <RANKING order="11" place="11" resultid="21953" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1258" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21586" />
                    <RANKING order="2" place="2" resultid="22019" />
                    <RANKING order="3" place="3" resultid="23421" />
                    <RANKING order="4" place="4" resultid="21188" />
                    <RANKING order="5" place="5" resultid="21897" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1259" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22988" />
                    <RANKING order="2" place="2" resultid="20735" />
                    <RANKING order="3" place="3" resultid="21937" />
                    <RANKING order="4" place="4" resultid="22457" />
                    <RANKING order="5" place="5" resultid="20640" />
                    <RANKING order="6" place="6" resultid="21907" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1260" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20647" />
                    <RANKING order="2" place="2" resultid="20956" />
                    <RANKING order="3" place="3" resultid="22924" />
                    <RANKING order="4" place="-1" resultid="20167" />
                    <RANKING order="5" place="-1" resultid="22913" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1261" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20259" />
                    <RANKING order="2" place="2" resultid="23061" />
                    <RANKING order="3" place="3" resultid="21822" />
                    <RANKING order="4" place="4" resultid="22026" />
                    <RANKING order="5" place="5" resultid="21755" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1262" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21750" />
                    <RANKING order="2" place="2" resultid="20218" />
                    <RANKING order="3" place="3" resultid="23353" />
                    <RANKING order="4" place="4" resultid="21686" />
                    <RANKING order="5" place="-1" resultid="21903" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1263" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20395" />
                    <RANKING order="2" place="2" resultid="21299" />
                    <RANKING order="3" place="3" resultid="22890" />
                    <RANKING order="4" place="4" resultid="22289" />
                    <RANKING order="5" place="5" resultid="23082" />
                    <RANKING order="6" place="6" resultid="22902" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1264" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21317" />
                    <RANKING order="2" place="2" resultid="21114" />
                    <RANKING order="3" place="3" resultid="23372" />
                    <RANKING order="4" place="4" resultid="20446" />
                    <RANKING order="5" place="-1" resultid="23405" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1265" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20409" />
                    <RANKING order="2" place="2" resultid="21378" />
                    <RANKING order="3" place="3" resultid="21608" />
                    <RANKING order="4" place="4" resultid="19910" />
                    <RANKING order="5" place="5" resultid="20484" />
                    <RANKING order="6" place="6" resultid="20709" />
                    <RANKING order="7" place="7" resultid="23855" />
                    <RANKING order="8" place="-1" resultid="20718" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1266" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21486" />
                    <RANKING order="2" place="2" resultid="22277" />
                    <RANKING order="3" place="3" resultid="19839" />
                    <RANKING order="4" place="4" resultid="21631" />
                    <RANKING order="5" place="5" resultid="22694" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1267" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20118" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1268" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19885" />
                    <RANKING order="2" place="2" resultid="21225" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1269" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1270" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1271" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1272" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24347" daytime="10:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24348" daytime="10:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24349" daytime="10:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24350" daytime="10:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="24351" daytime="10:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="24352" daytime="10:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="24353" daytime="10:30" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1358" daytime="11:30" gender="F" number="18" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="16646" agemax="99" agemin="80" calculate="TOTAL" />
                <AGEGROUP agegroupid="16647" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21961" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16648" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22089" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16649" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21210" />
                    <RANKING order="2" place="2" resultid="21767" />
                    <RANKING order="3" place="3" resultid="22928" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16650" agemax="239" agemin="200" calculate="TOTAL" />
                <AGEGROUP agegroupid="16651" agemax="279" agemin="240" calculate="TOTAL" />
                <AGEGROUP agegroupid="16652" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19922" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24372" daytime="11:30" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1205" daytime="09:10" gender="M" number="11" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1206" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21955" />
                    <RANKING order="2" place="2" resultid="23398" />
                    <RANKING order="3" place="3" resultid="21561" />
                    <RANKING order="4" place="4" resultid="23380" />
                    <RANKING order="5" place="5" resultid="23386" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1207" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21542" />
                    <RANKING order="2" place="2" resultid="21547" />
                    <RANKING order="3" place="3" resultid="22049" />
                    <RANKING order="4" place="4" resultid="22668" />
                    <RANKING order="5" place="5" resultid="22974" />
                    <RANKING order="6" place="6" resultid="21281" />
                    <RANKING order="7" place="7" resultid="21663" />
                    <RANKING order="8" place="8" resultid="22681" />
                    <RANKING order="9" place="9" resultid="21509" />
                    <RANKING order="10" place="10" resultid="19785" />
                    <RANKING order="11" place="11" resultid="20947" />
                    <RANKING order="12" place="12" resultid="23074" />
                    <RANKING order="13" place="13" resultid="20632" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1208" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19847" />
                    <RANKING order="2" place="2" resultid="22996" />
                    <RANKING order="3" place="3" resultid="21250" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1209" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="23005" />
                    <RANKING order="2" place="2" resultid="22506" />
                    <RANKING order="3" place="3" resultid="21158" />
                    <RANKING order="4" place="4" resultid="20506" />
                    <RANKING order="5" place="5" resultid="20654" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1210" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22933" />
                    <RANKING order="2" place="2" resultid="22340" />
                    <RANKING order="3" place="3" resultid="21858" />
                    <RANKING order="4" place="4" resultid="21451" />
                    <RANKING order="5" place="5" resultid="20195" />
                    <RANKING order="6" place="6" resultid="20110" />
                    <RANKING order="7" place="7" resultid="22942" />
                    <RANKING order="8" place="8" resultid="22252" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1211" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20727" />
                    <RANKING order="2" place="2" resultid="19966" />
                    <RANKING order="3" place="3" resultid="22957" />
                    <RANKING order="4" place="4" resultid="21828" />
                    <RANKING order="5" place="5" resultid="23092" />
                    <RANKING order="6" place="6" resultid="21592" />
                    <RANKING order="7" place="7" resultid="21477" />
                    <RANKING order="8" place="8" resultid="22040" />
                    <RANKING order="9" place="9" resultid="21183" />
                    <RANKING order="10" place="10" resultid="23368" />
                    <RANKING order="11" place="-1" resultid="21304" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1212" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20240" />
                    <RANKING order="2" place="2" resultid="21234" />
                    <RANKING order="3" place="3" resultid="21353" />
                    <RANKING order="4" place="4" resultid="20226" />
                    <RANKING order="5" place="5" resultid="22895" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1213" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21257" />
                    <RANKING order="2" place="2" resultid="21344" />
                    <RANKING order="3" place="3" resultid="20277" />
                    <RANKING order="4" place="4" resultid="20470" />
                    <RANKING order="5" place="-1" resultid="20402" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1214" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21121" />
                    <RANKING order="2" place="2" resultid="21151" />
                    <RANKING order="3" place="3" resultid="19859" />
                    <RANKING order="4" place="4" resultid="21623" />
                    <RANKING order="5" place="5" resultid="21469" />
                    <RANKING order="6" place="6" resultid="20455" />
                    <RANKING order="7" place="7" resultid="20462" />
                    <RANKING order="8" place="8" resultid="21241" />
                    <RANKING order="9" place="9" resultid="22306" />
                    <RANKING order="10" place="-1" resultid="19796" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1215" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21844" />
                    <RANKING order="2" place="2" resultid="23429" />
                    <RANKING order="3" place="3" resultid="20142" />
                    <RANKING order="4" place="4" resultid="19774" />
                    <RANKING order="5" place="5" resultid="21972" />
                    <RANKING order="6" place="-1" resultid="20961" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1216" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21105" />
                    <RANKING order="2" place="2" resultid="19878" />
                    <RANKING order="3" place="3" resultid="20263" />
                    <RANKING order="4" place="4" resultid="20515" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1217" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21460" />
                    <RANKING order="2" place="2" resultid="22425" />
                    <RANKING order="3" place="3" resultid="22625" />
                    <RANKING order="4" place="4" resultid="20438" />
                    <RANKING order="5" place="5" resultid="20124" />
                    <RANKING order="6" place="-1" resultid="20150" />
                    <RANKING order="7" place="-1" resultid="20939" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1218" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22651" />
                    <RANKING order="2" place="2" resultid="20890" />
                    <RANKING order="3" place="3" resultid="21989" />
                    <RANKING order="4" place="4" resultid="22416" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1219" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20701" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1220" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1221" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24328" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24329" daytime="09:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24330" daytime="09:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24331" daytime="09:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="24332" daytime="09:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="24333" daytime="09:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="24334" daytime="09:20" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="24335" daytime="09:20" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="24336" daytime="09:20" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1273" daytime="10:35" gender="M" number="15" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1274" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="23399" />
                    <RANKING order="2" place="2" resultid="20308" />
                    <RANKING order="3" place="3" resultid="21428" />
                    <RANKING order="4" place="4" resultid="23381" />
                    <RANKING order="5" place="5" resultid="21562" />
                    <RANKING order="6" place="6" resultid="21437" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1275" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22669" />
                    <RANKING order="2" place="2" resultid="22442" />
                    <RANKING order="3" place="3" resultid="21664" />
                    <RANKING order="4" place="4" resultid="22968" />
                    <RANKING order="5" place="5" resultid="22975" />
                    <RANKING order="6" place="6" resultid="21096" />
                    <RANKING order="7" place="7" resultid="21931" />
                    <RANKING order="8" place="8" resultid="20303" />
                    <RANKING order="9" place="9" resultid="21510" />
                    <RANKING order="10" place="10" resultid="23358" />
                    <RANKING order="11" place="11" resultid="21941" />
                    <RANKING order="12" place="12" resultid="21945" />
                    <RANKING order="13" place="13" resultid="22659" />
                    <RANKING order="14" place="14" resultid="19786" />
                    <RANKING order="15" place="15" resultid="20633" />
                    <RANKING order="16" place="16" resultid="22643" />
                    <RANKING order="17" place="17" resultid="21913" />
                    <RANKING order="18" place="-1" resultid="21949" />
                    <RANKING order="19" place="-1" resultid="22682" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1276" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22409" />
                    <RANKING order="2" place="2" resultid="21920" />
                    <RANKING order="3" place="3" resultid="21251" />
                    <RANKING order="4" place="4" resultid="21707" />
                    <RANKING order="5" place="5" resultid="22462" />
                    <RANKING order="6" place="6" resultid="19848" />
                    <RANKING order="7" place="7" resultid="22997" />
                    <RANKING order="8" place="8" resultid="21693" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1277" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22332" />
                    <RANKING order="2" place="2" resultid="20234" />
                    <RANKING order="3" place="3" resultid="19758" />
                    <RANKING order="4" place="4" resultid="20507" />
                    <RANKING order="5" place="5" resultid="21696" />
                    <RANKING order="6" place="6" resultid="20625" />
                    <RANKING order="7" place="7" resultid="21916" />
                    <RANKING order="8" place="-1" resultid="22507" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1278" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22341" />
                    <RANKING order="2" place="2" resultid="22617" />
                    <RANKING order="3" place="3" resultid="22323" />
                    <RANKING order="4" place="4" resultid="22070" />
                    <RANKING order="5" place="5" resultid="21167" />
                    <RANKING order="6" place="6" resultid="22478" />
                    <RANKING order="7" place="7" resultid="21679" />
                    <RANKING order="8" place="8" resultid="22489" />
                    <RANKING order="9" place="9" resultid="21850" />
                    <RANKING order="10" place="10" resultid="22241" />
                    <RANKING order="11" place="11" resultid="22379" />
                    <RANKING order="12" place="12" resultid="21600" />
                    <RANKING order="13" place="-1" resultid="20111" />
                    <RANKING order="14" place="-1" resultid="22943" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1279" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20173" />
                    <RANKING order="2" place="2" resultid="22032" />
                    <RANKING order="3" place="3" resultid="20728" />
                    <RANKING order="4" place="4" resultid="19967" />
                    <RANKING order="5" place="5" resultid="20286" />
                    <RANKING order="6" place="6" resultid="21829" />
                    <RANKING order="7" place="7" resultid="21478" />
                    <RANKING order="8" place="8" resultid="21879" />
                    <RANKING order="9" place="9" resultid="21593" />
                    <RANKING order="10" place="10" resultid="21401" />
                    <RANKING order="11" place="11" resultid="23093" />
                    <RANKING order="12" place="12" resultid="19975" />
                    <RANKING order="13" place="13" resultid="23369" />
                    <RANKING order="14" place="14" resultid="22041" />
                    <RANKING order="15" place="15" resultid="21184" />
                    <RANKING order="16" place="16" resultid="21711" />
                    <RANKING order="17" place="17" resultid="22403" />
                    <RANKING order="18" place="-1" resultid="20269" />
                    <RANKING order="19" place="-1" resultid="20415" />
                    <RANKING order="20" place="-1" resultid="21219" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1280" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22877" />
                    <RANKING order="2" place="2" resultid="20910" />
                    <RANKING order="3" place="3" resultid="21100" />
                    <RANKING order="4" place="4" resultid="21981" />
                    <RANKING order="5" place="5" resultid="20932" />
                    <RANKING order="6" place="6" resultid="19811" />
                    <RANKING order="7" place="7" resultid="21672" />
                    <RANKING order="8" place="-1" resultid="21140" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1281" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22467" />
                    <RANKING order="2" place="2" resultid="20278" />
                    <RANKING order="3" place="3" resultid="20471" />
                    <RANKING order="4" place="4" resultid="20403" />
                    <RANKING order="5" place="5" resultid="22064" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1282" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21122" />
                    <RANKING order="2" place="2" resultid="21265" />
                    <RANKING order="3" place="3" resultid="19860" />
                    <RANKING order="4" place="4" resultid="21529" />
                    <RANKING order="5" place="5" resultid="20693" />
                    <RANKING order="6" place="6" resultid="21624" />
                    <RANKING order="7" place="7" resultid="22395" />
                    <RANKING order="8" place="8" resultid="20463" />
                    <RANKING order="9" place="9" resultid="21242" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1283" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22452" />
                    <RANKING order="2" place="2" resultid="19775" />
                    <RANKING order="3" place="3" resultid="20492" />
                    <RANKING order="4" place="4" resultid="19947" />
                    <RANKING order="5" place="-1" resultid="20962" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1284" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21326" />
                    <RANKING order="2" place="2" resultid="21135" />
                    <RANKING order="3" place="3" resultid="19875" />
                    <RANKING order="4" place="4" resultid="19931" />
                    <RANKING order="5" place="-1" resultid="20160" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1285" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21461" />
                    <RANKING order="2" place="2" resultid="21637" />
                    <RANKING order="3" place="3" resultid="22426" />
                    <RANKING order="4" place="4" resultid="22626" />
                    <RANKING order="5" place="5" resultid="21371" />
                    <RANKING order="6" place="6" resultid="20125" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1286" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1287" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20702" />
                    <RANKING order="2" place="2" resultid="21496" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1288" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1289" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24354" daytime="10:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24355" daytime="10:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24356" daytime="10:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24357" daytime="10:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="24358" daytime="10:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="24359" daytime="10:45" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="24360" daytime="10:50" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="24361" daytime="10:50" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="24362" daytime="10:50" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="24363" daytime="10:55" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="24364" daytime="10:55" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="24365" daytime="11:00" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2019-06-01" daytime="16:00" endtime="20:21" name="BLOK III" number="3" warmupfrom="15:00">
          <EVENTS>
            <EVENT eventid="1508" daytime="17:45" gender="M" number="27" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1509" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20309" />
                    <RANKING order="2" place="-1" resultid="19954" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1510" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21284" />
                    <RANKING order="2" place="2" resultid="22051" />
                    <RANKING order="3" place="3" resultid="22976" />
                    <RANKING order="4" place="4" resultid="22969" />
                    <RANKING order="5" place="5" resultid="21666" />
                    <RANKING order="6" place="6" resultid="20188" />
                    <RANKING order="7" place="7" resultid="20304" />
                    <RANKING order="8" place="8" resultid="21512" />
                    <RANKING order="9" place="9" resultid="19787" />
                    <RANKING order="10" place="10" resultid="20635" />
                    <RANKING order="11" place="11" resultid="21914" />
                    <RANKING order="12" place="-1" resultid="21887" />
                    <RANKING order="13" place="-1" resultid="22645" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1511" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19849" />
                    <RANKING order="2" place="2" resultid="22463" />
                    <RANKING order="3" place="3" resultid="21503" />
                    <RANKING order="4" place="4" resultid="21708" />
                    <RANKING order="5" place="5" resultid="22411" />
                    <RANKING order="6" place="6" resultid="21922" />
                    <RANKING order="7" place="7" resultid="21253" />
                    <RANKING order="8" place="-1" resultid="20501" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1512" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19759" />
                    <RANKING order="2" place="2" resultid="22358" />
                    <RANKING order="3" place="3" resultid="19782" />
                    <RANKING order="4" place="4" resultid="20627" />
                    <RANKING order="5" place="5" resultid="21917" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1513" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20685" />
                    <RANKING order="2" place="2" resultid="22071" />
                    <RANKING order="3" place="3" resultid="22479" />
                    <RANKING order="4" place="4" resultid="22325" />
                    <RANKING order="5" place="5" resultid="22343" />
                    <RANKING order="6" place="6" resultid="22491" />
                    <RANKING order="7" place="7" resultid="20952" />
                    <RANKING order="8" place="8" resultid="21852" />
                    <RANKING order="9" place="9" resultid="22475" />
                    <RANKING order="10" place="10" resultid="21601" />
                    <RANKING order="11" place="11" resultid="22242" />
                    <RANKING order="12" place="12" resultid="22391" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1514" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20175" />
                    <RANKING order="2" place="2" resultid="22033" />
                    <RANKING order="3" place="3" resultid="20417" />
                    <RANKING order="4" place="4" resultid="21831" />
                    <RANKING order="5" place="5" resultid="21595" />
                    <RANKING order="6" place="6" resultid="21404" />
                    <RANKING order="7" place="7" resultid="21480" />
                    <RANKING order="8" place="8" resultid="22043" />
                    <RANKING order="9" place="9" resultid="19977" />
                    <RANKING order="10" place="10" resultid="21713" />
                    <RANKING order="11" place="11" resultid="22405" />
                    <RANKING order="12" place="-1" resultid="20271" />
                    <RANKING order="13" place="-1" resultid="21220" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1515" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22879" />
                    <RANKING order="2" place="2" resultid="20912" />
                    <RANKING order="3" place="3" resultid="21984" />
                    <RANKING order="4" place="4" resultid="20934" />
                    <RANKING order="5" place="5" resultid="21674" />
                    <RANKING order="6" place="6" resultid="22384" />
                    <RANKING order="7" place="7" resultid="22898" />
                    <RANKING order="8" place="-1" resultid="19984" />
                    <RANKING order="9" place="-1" resultid="21142" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1516" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22468" />
                    <RANKING order="2" place="2" resultid="20473" />
                    <RANKING order="3" place="3" resultid="20405" />
                    <RANKING order="4" place="4" resultid="22065" />
                    <RANKING order="5" place="5" resultid="20181" />
                    <RANKING order="6" place="6" resultid="22271" />
                    <RANKING order="7" place="-1" resultid="19805" />
                    <RANKING order="8" place="-1" resultid="20919" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1517" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21124" />
                    <RANKING order="2" place="2" resultid="21530" />
                    <RANKING order="3" place="3" resultid="20694" />
                    <RANKING order="4" place="4" resultid="21626" />
                    <RANKING order="5" place="5" resultid="22397" />
                    <RANKING order="6" place="6" resultid="22309" />
                    <RANKING order="7" place="-1" resultid="21524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1518" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20494" />
                    <RANKING order="2" place="2" resultid="20964" />
                    <RANKING order="3" place="3" resultid="19949" />
                    <RANKING order="4" place="-1" resultid="19776" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1519" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21328" />
                    <RANKING order="2" place="2" resultid="20161" />
                    <RANKING order="3" place="3" resultid="20517" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1520" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22628" />
                    <RANKING order="2" place="2" resultid="21639" />
                    <RANKING order="3" place="3" resultid="22428" />
                    <RANKING order="4" place="4" resultid="21372" />
                    <RANKING order="5" place="5" resultid="20127" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1521" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22654" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1522" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20704" />
                    <RANKING order="2" place="2" resultid="21498" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1523" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1524" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24415" daytime="17:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24416" daytime="17:55" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24417" daytime="18:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24418" daytime="18:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="24419" daytime="18:05" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="24420" daytime="18:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="24421" daytime="18:15" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="24422" daytime="18:20" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="24423" daytime="18:20" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="24424" daytime="18:25" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1474" daytime="17:05" gender="M" number="25" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1475" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21956" />
                    <RANKING order="2" place="2" resultid="23387" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1476" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21544" />
                    <RANKING order="2" place="2" resultid="21548" />
                    <RANKING order="3" place="3" resultid="22684" />
                    <RANKING order="4" place="4" resultid="21386" />
                    <RANKING order="5" place="5" resultid="20948" />
                    <RANKING order="6" place="-1" resultid="23077" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1477" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22612" />
                    <RANKING order="2" place="2" resultid="22999" />
                    <RANKING order="3" place="3" resultid="21252" />
                    <RANKING order="4" place="4" resultid="22247" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1478" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22509" />
                    <RANKING order="2" place="2" resultid="23008" />
                    <RANKING order="3" place="3" resultid="21160" />
                    <RANKING order="4" place="4" resultid="20508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1479" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22342" />
                    <RANKING order="2" place="2" resultid="21580" />
                    <RANKING order="3" place="3" resultid="21859" />
                    <RANKING order="4" place="4" resultid="20198" />
                    <RANKING order="5" place="5" resultid="22253" />
                    <RANKING order="6" place="-1" resultid="20113" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1480" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20730" />
                    <RANKING order="2" place="2" resultid="19968" />
                    <RANKING order="3" place="3" resultid="21830" />
                    <RANKING order="4" place="4" resultid="23094" />
                    <RANKING order="5" place="5" resultid="21307" />
                    <RANKING order="6" place="6" resultid="21403" />
                    <RANKING order="7" place="7" resultid="22042" />
                    <RANKING order="8" place="-1" resultid="20416" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1481" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20241" />
                    <RANKING order="2" place="2" resultid="21983" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1482" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21258" />
                    <RANKING order="2" place="2" resultid="21347" />
                    <RANKING order="3" place="-1" resultid="20280" />
                    <RANKING order="4" place="-1" resultid="20404" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1483" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21154" />
                    <RANKING order="2" place="2" resultid="19862" />
                    <RANKING order="3" place="3" resultid="21470" />
                    <RANKING order="4" place="4" resultid="20456" />
                    <RANKING order="5" place="5" resultid="21244" />
                    <RANKING order="6" place="-1" resultid="21123" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1484" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22453" />
                    <RANKING order="2" place="2" resultid="23431" />
                    <RANKING order="3" place="3" resultid="20144" />
                    <RANKING order="4" place="4" resultid="21975" />
                    <RANKING order="5" place="-1" resultid="20963" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1485" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21108" />
                    <RANKING order="2" place="2" resultid="19879" />
                    <RANKING order="3" place="3" resultid="20264" />
                    <RANKING order="4" place="4" resultid="20388" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1486" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21463" />
                    <RANKING order="2" place="2" resultid="22427" />
                    <RANKING order="3" place="3" resultid="20941" />
                    <RANKING order="4" place="4" resultid="20441" />
                    <RANKING order="5" place="5" resultid="20126" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1487" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20893" />
                    <RANKING order="2" place="2" resultid="21990" />
                    <RANKING order="3" place="3" resultid="22419" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1488" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1489" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1490" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24403" daytime="17:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24404" daytime="17:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24405" daytime="17:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24406" daytime="17:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="24407" daytime="17:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="24408" daytime="17:15" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1548" daytime="18:30" gender="M" number="29" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="16667" agemax="99" agemin="80" calculate="TOTAL" />
                <AGEGROUP agegroupid="16668" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22688" />
                    <RANKING order="2" place="2" resultid="21966" />
                    <RANKING order="3" place="-1" resultid="21967" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16669" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22513" />
                    <RANKING order="2" place="2" resultid="22091" />
                    <RANKING order="3" place="3" resultid="21717" />
                    <RANKING order="4" place="4" resultid="22979" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16670" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22980" />
                    <RANKING order="2" place="2" resultid="22369" />
                    <RANKING order="3" place="3" resultid="21423" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16671" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21890" />
                    <RANKING order="2" place="-1" resultid="21207" />
                    <RANKING order="3" place="-1" resultid="22370" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16672" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22006" />
                    <RANKING order="2" place="2" resultid="21209" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16673" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19925" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24426" daytime="18:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24427" daytime="18:35" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1457" daytime="16:50" gender="F" number="24" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1458" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21199" />
                    <RANKING order="2" place="2" resultid="21557" />
                    <RANKING order="3" place="3" resultid="22920" />
                    <RANKING order="4" place="4" resultid="20754" />
                    <RANKING order="5" place="5" resultid="22364" />
                    <RANKING order="6" place="6" resultid="23394" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1459" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21553" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1460" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="1461" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20648" />
                    <RANKING order="2" place="2" resultid="22884" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1462" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21179" />
                    <RANKING order="2" place="2" resultid="22027" />
                    <RANKING order="3" place="2" resultid="22258" />
                    <RANKING order="4" place="4" resultid="21823" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1463" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21173" />
                    <RANKING order="2" place="2" resultid="21733" />
                    <RANKING order="3" place="3" resultid="20219" />
                    <RANKING order="4" place="4" resultid="23355" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1464" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22891" />
                    <RANKING order="2" place="2" resultid="21301" />
                    <RANKING order="3" place="3" resultid="22290" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1465" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21116" />
                    <RANKING order="2" place="2" resultid="21865" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1466" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21517" />
                    <RANKING order="2" place="2" resultid="20410" />
                    <RANKING order="3" place="3" resultid="19911" />
                    <RANKING order="4" place="4" resultid="20485" />
                    <RANKING order="5" place="5" resultid="22908" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1467" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19871" />
                    <RANKING order="2" place="2" resultid="21632" />
                    <RANKING order="3" place="3" resultid="22695" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1468" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20119" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1469" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1470" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1471" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1472" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1473" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24399" daytime="16:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24400" daytime="16:55" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24401" daytime="17:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24402" daytime="17:00" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1406" daytime="16:15" gender="M" number="21" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1407" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="23400" />
                    <RANKING order="2" place="2" resultid="21438" />
                    <RANKING order="3" place="3" resultid="21429" />
                    <RANKING order="4" place="4" resultid="20970" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1408" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22619" />
                    <RANKING order="2" place="2" resultid="21568" />
                    <RANKING order="3" place="3" resultid="23076" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1409" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21704" />
                    <RANKING order="2" place="2" resultid="20500" />
                    <RANKING order="3" place="3" resultid="21725" />
                    <RANKING order="4" place="4" resultid="22246" />
                    <RANKING order="5" place="5" resultid="23088" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1410" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22333" />
                    <RANKING order="2" place="2" resultid="22085" />
                    <RANKING order="3" place="-1" resultid="22078" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1411" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21168" />
                    <RANKING order="2" place="2" resultid="22474" />
                    <RANKING order="3" place="3" resultid="21453" />
                    <RANKING order="4" place="4" resultid="21851" />
                    <RANKING order="5" place="5" resultid="20197" />
                    <RANKING order="6" place="6" resultid="23416" />
                    <RANKING order="7" place="7" resultid="22380" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1412" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20902" />
                    <RANKING order="2" place="2" resultid="21417" />
                    <RANKING order="3" place="3" resultid="22958" />
                    <RANKING order="4" place="4" resultid="21306" />
                    <RANKING order="5" place="5" resultid="22404" />
                    <RANKING order="6" place="6" resultid="21712" />
                    <RANKING order="7" place="-1" resultid="20270" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1413" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21574" />
                    <RANKING order="2" place="2" resultid="21236" />
                    <RANKING order="3" place="3" resultid="21193" />
                    <RANKING order="4" place="4" resultid="21355" />
                    <RANKING order="5" place="5" resultid="21673" />
                    <RANKING order="6" place="6" resultid="22383" />
                    <RANKING order="7" place="7" resultid="22897" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1414" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22315" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1415" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21999" />
                    <RANKING order="2" place="2" resultid="22447" />
                    <RANKING order="3" place="3" resultid="23411" />
                    <RANKING order="4" place="4" resultid="21243" />
                    <RANKING order="5" place="-1" resultid="19798" />
                    <RANKING order="6" place="-1" resultid="21153" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1416" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22434" />
                    <RANKING order="2" place="2" resultid="20885" />
                    <RANKING order="3" place="3" resultid="20423" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1417" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21107" />
                    <RANKING order="2" place="2" resultid="19932" />
                    <RANKING order="3" place="3" resultid="20135" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1418" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19889" />
                    <RANKING order="2" place="2" resultid="19940" />
                    <RANKING order="3" place="3" resultid="20440" />
                    <RANKING order="4" place="-1" resultid="20152" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1419" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20892" />
                    <RANKING order="2" place="2" resultid="22418" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1420" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20703" />
                    <RANKING order="2" place="2" resultid="21497" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1421" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1422" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24380" daytime="16:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24381" daytime="16:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24382" daytime="16:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24383" daytime="16:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="24384" daytime="16:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="24385" daytime="16:30" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1491" daytime="17:20" gender="F" number="26" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1492" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21293" />
                    <RANKING order="2" place="2" resultid="22665" />
                    <RANKING order="3" place="3" resultid="20755" />
                    <RANKING order="4" place="4" resultid="20761" />
                    <RANKING order="5" place="-1" resultid="21558" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1493" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21587" />
                    <RANKING order="2" place="2" resultid="22020" />
                    <RANKING order="3" place="3" resultid="22059" />
                    <RANKING order="4" place="4" resultid="23423" />
                    <RANKING order="5" place="5" resultid="21189" />
                    <RANKING order="6" place="6" resultid="22639" />
                    <RANKING order="7" place="7" resultid="21898" />
                    <RANKING order="8" place="-1" resultid="21204" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1494" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22990" />
                    <RANKING order="2" place="2" resultid="21938" />
                    <RANKING order="3" place="3" resultid="22459" />
                    <RANKING order="4" place="4" resultid="20641" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1495" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20649" />
                    <RANKING order="2" place="2" resultid="22496" />
                    <RANKING order="3" place="3" resultid="22915" />
                    <RANKING order="4" place="4" resultid="22925" />
                    <RANKING order="5" place="-1" resultid="21764" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1496" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20260" />
                    <RANKING order="2" place="2" resultid="21410" />
                    <RANKING order="3" place="3" resultid="19791" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1497" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19902" />
                    <RANKING order="2" place="2" resultid="21751" />
                    <RANKING order="3" place="3" resultid="20220" />
                    <RANKING order="4" place="4" resultid="21841" />
                    <RANKING order="5" place="5" resultid="23364" />
                    <RANKING order="6" place="6" resultid="21688" />
                    <RANKING order="7" place="7" resultid="21365" />
                    <RANKING order="8" place="-1" resultid="21904" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1498" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20396" />
                    <RANKING order="2" place="2" resultid="22291" />
                    <RANKING order="3" place="3" resultid="23084" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1499" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21320" />
                    <RANKING order="2" place="2" resultid="22484" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1500" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20411" />
                    <RANKING order="2" place="2" resultid="21610" />
                    <RANKING order="3" place="3" resultid="19912" />
                    <RANKING order="4" place="4" resultid="21618" />
                    <RANKING order="5" place="5" resultid="20711" />
                    <RANKING order="6" place="-1" resultid="20486" />
                    <RANKING order="7" place="-1" resultid="20720" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1501" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21488" />
                    <RANKING order="2" place="2" resultid="22279" />
                    <RANKING order="3" place="3" resultid="19841" />
                    <RANKING order="4" place="4" resultid="21633" />
                    <RANKING order="5" place="5" resultid="22696" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1502" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20120" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1503" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19886" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1504" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1505" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1506" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1507" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24409" daytime="17:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24410" daytime="17:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24411" daytime="17:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24412" daytime="17:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="24413" daytime="17:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="24414" daytime="17:45" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1525" daytime="18:25" gender="F" number="28" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="16660" agemax="99" agemin="80" calculate="TOTAL" />
                <AGEGROUP agegroupid="16661" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21962" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16662" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22090" />
                    <RANKING order="2" place="2" resultid="22927" />
                    <RANKING order="3" place="3" resultid="21963" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16663" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21211" />
                    <RANKING order="2" place="2" resultid="21768" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16664" agemax="239" agemin="200" calculate="TOTAL" />
                <AGEGROUP agegroupid="16665" agemax="279" agemin="240" calculate="TOTAL" />
                <AGEGROUP agegroupid="16666" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19924" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24425" daytime="18:25" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1578" daytime="18:55" gender="M" number="31" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1579" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22319" />
                    <RANKING order="2" place="2" resultid="23388" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1580" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22052" />
                    <RANKING order="2" place="2" resultid="22970" />
                    <RANKING order="3" place="3" resultid="20189" />
                    <RANKING order="4" place="4" resultid="21933" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1581" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19850" />
                    <RANKING order="2" place="2" resultid="21726" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1582" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20509" />
                    <RANKING order="2" place="2" resultid="22086" />
                    <RANKING order="3" place="3" resultid="22359" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1583" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20686" />
                    <RANKING order="2" place="2" resultid="22072" />
                    <RANKING order="3" place="3" resultid="19765" />
                    <RANKING order="4" place="4" resultid="21581" />
                    <RANKING order="5" place="5" resultid="19769" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1584" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22034" />
                    <RANKING order="2" place="2" resultid="20903" />
                    <RANKING order="3" place="3" resultid="19969" />
                    <RANKING order="4" place="4" resultid="21418" />
                    <RANKING order="5" place="-1" resultid="21874" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1585" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20255" />
                    <RANKING order="2" place="2" resultid="19817" />
                    <RANKING order="3" place="3" resultid="20229" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1586" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20182" />
                    <RANKING order="2" place="-1" resultid="19806" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1587" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21471" />
                    <RANKING order="2" place="2" resultid="22448" />
                    <RANKING order="3" place="3" resultid="20457" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1588" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22435" />
                    <RANKING order="2" place="2" resultid="20145" />
                    <RANKING order="3" place="3" resultid="23432" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1589" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21329" />
                    <RANKING order="2" place="2" resultid="22674" />
                    <RANKING order="3" place="3" resultid="20389" />
                    <RANKING order="4" place="4" resultid="20518" />
                    <RANKING order="5" place="-1" resultid="20136" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1590" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19941" />
                    <RANKING order="2" place="2" resultid="20942" />
                    <RANKING order="3" place="-1" resultid="20153" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1591" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1592" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1593" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1594" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24430" daytime="18:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24431" daytime="19:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24432" daytime="19:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24433" daytime="19:25" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1388" daytime="16:00" gender="F" number="20" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1390" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22299" />
                    <RANKING order="2" place="2" resultid="21444" />
                    <RANKING order="3" place="3" resultid="20745" />
                    <RANKING order="4" place="4" resultid="23068" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1391" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20777" />
                    <RANKING order="2" place="2" resultid="21203" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1392" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22989" />
                    <RANKING order="2" place="2" resultid="21926" />
                    <RANKING order="3" place="3" resultid="21742" />
                    <RANKING order="4" place="4" resultid="21995" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1393" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22914" />
                    <RANKING order="2" place="-1" resultid="21763" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1394" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20246" />
                    <RANKING order="2" place="2" resultid="21178" />
                    <RANKING order="3" place="3" resultid="19790" />
                    <RANKING order="4" place="4" resultid="22953" />
                    <RANKING order="5" place="5" resultid="21756" />
                    <RANKING order="6" place="6" resultid="21274" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1395" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19901" />
                    <RANKING order="2" place="2" resultid="21687" />
                    <RANKING order="3" place="3" resultid="21840" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1396" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20205" />
                    <RANKING order="2" place="2" resultid="22903" />
                    <RANKING order="3" place="3" resultid="23083" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1397" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22483" />
                    <RANKING order="2" place="2" resultid="23373" />
                    <RANKING order="3" place="-1" resultid="23406" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1398" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22284" />
                    <RANKING order="2" place="2" resultid="22633" />
                    <RANKING order="3" place="3" resultid="21609" />
                    <RANKING order="4" place="4" resultid="21617" />
                    <RANKING order="5" place="5" resultid="22907" />
                    <RANKING order="6" place="6" resultid="23854" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1399" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22278" />
                    <RANKING order="2" place="2" resultid="19840" />
                    <RANKING order="3" place="3" resultid="19855" />
                    <RANKING order="4" place="4" resultid="20449" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1400" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19919" />
                    <RANKING order="2" place="2" resultid="21230" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1401" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19894" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1402" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1403" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1404" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1405" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24375" daytime="16:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24376" daytime="16:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24377" daytime="16:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24378" daytime="16:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="24379" daytime="16:10" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1555" daytime="18:40" gender="F" number="30" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1562" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22300" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1563" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="1564" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22014" />
                    <RANKING order="2" place="2" resultid="22502" />
                    <RANKING order="3" place="3" resultid="21743" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1565" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22949" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1566" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21411" />
                    <RANKING order="2" place="2" resultid="21538" />
                    <RANKING order="3" place="3" resultid="23435" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1567" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21734" />
                    <RANKING order="2" place="2" resultid="21312" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1568" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="1569" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21866" />
                    <RANKING order="2" place="2" resultid="21338" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1570" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21518" />
                    <RANKING order="2" place="2" resultid="21381" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1571" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1572" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1573" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1574" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1575" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1576" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1577" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24428" daytime="18:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24429" daytime="18:50" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1423" daytime="16:30" gender="F" number="22" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1424" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20769" />
                    <RANKING order="2" place="2" resultid="21292" />
                    <RANKING order="3" place="3" resultid="20746" />
                    <RANKING order="4" place="4" resultid="22363" />
                    <RANKING order="5" place="5" resultid="21445" />
                    <RANKING order="6" place="-1" resultid="23069" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1425" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22058" />
                    <RANKING order="2" place="2" resultid="23422" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1426" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20736" />
                    <RANKING order="2" place="2" resultid="22013" />
                    <RANKING order="3" place="3" resultid="22458" />
                    <RANKING order="4" place="4" resultid="22501" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1427" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22495" />
                    <RANKING order="2" place="-1" resultid="20168" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1428" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20247" />
                    <RANKING order="2" place="2" resultid="21146" />
                    <RANKING order="3" place="3" resultid="21757" />
                    <RANKING order="4" place="4" resultid="21537" />
                    <RANKING order="5" place="-1" resultid="19907" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1429" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21130" />
                    <RANKING order="2" place="2" resultid="21311" />
                    <RANKING order="3" place="3" resultid="23354" />
                    <RANKING order="4" place="4" resultid="21364" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1430" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21300" />
                    <RANKING order="2" place="2" resultid="20206" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1431" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21115" />
                    <RANKING order="2" place="2" resultid="21319" />
                    <RANKING order="3" place="3" resultid="23374" />
                    <RANKING order="4" place="4" resultid="21337" />
                    <RANKING order="5" place="-1" resultid="23407" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1432" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22634" />
                    <RANKING order="2" place="2" resultid="21380" />
                    <RANKING order="3" place="3" resultid="20719" />
                    <RANKING order="4" place="4" resultid="20710" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1433" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19870" />
                    <RANKING order="2" place="2" resultid="21487" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1434" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1435" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19895" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1436" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1437" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1438" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1439" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24386" daytime="16:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24387" daytime="16:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24388" daytime="16:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24389" daytime="16:35" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1440" daytime="16:35" gender="M" number="23" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1441" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="23401" />
                    <RANKING order="2" place="2" resultid="21430" />
                    <RANKING order="3" place="3" resultid="22964" />
                    <RANKING order="4" place="4" resultid="23382" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1442" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22670" />
                    <RANKING order="2" place="2" resultid="22620" />
                    <RANKING order="3" place="3" resultid="21665" />
                    <RANKING order="4" place="4" resultid="20433" />
                    <RANKING order="5" place="5" resultid="21886" />
                    <RANKING order="6" place="6" resultid="21932" />
                    <RANKING order="7" place="7" resultid="22443" />
                    <RANKING order="8" place="8" resultid="21569" />
                    <RANKING order="9" place="9" resultid="21283" />
                    <RANKING order="10" place="10" resultid="23359" />
                    <RANKING order="11" place="11" resultid="22683" />
                    <RANKING order="12" place="12" resultid="22660" />
                    <RANKING order="13" place="13" resultid="21511" />
                    <RANKING order="14" place="14" resultid="20634" />
                    <RANKING order="15" place="-1" resultid="21385" />
                    <RANKING order="16" place="-1" resultid="21543" />
                    <RANKING order="17" place="-1" resultid="21942" />
                    <RANKING order="18" place="-1" resultid="21946" />
                    <RANKING order="19" place="-1" resultid="21950" />
                    <RANKING order="20" place="-1" resultid="22644" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1443" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22410" />
                    <RANKING order="2" place="2" resultid="21921" />
                    <RANKING order="3" place="3" resultid="22998" />
                    <RANKING order="4" place="4" resultid="22264" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1444" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22508" />
                    <RANKING order="2" place="2" resultid="23007" />
                    <RANKING order="3" place="3" resultid="21159" />
                    <RANKING order="4" place="4" resultid="22334" />
                    <RANKING order="5" place="5" resultid="20235" />
                    <RANKING order="6" place="6" resultid="20626" />
                    <RANKING order="7" place="-1" resultid="22079" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1445" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22934" />
                    <RANKING order="2" place="2" resultid="22938" />
                    <RANKING order="3" place="3" resultid="21454" />
                    <RANKING order="4" place="4" resultid="22324" />
                    <RANKING order="5" place="5" resultid="22490" />
                    <RANKING order="6" place="6" resultid="21169" />
                    <RANKING order="7" place="7" resultid="21680" />
                    <RANKING order="8" place="8" resultid="20951" />
                    <RANKING order="9" place="-1" resultid="20112" />
                    <RANKING order="10" place="-1" resultid="22946" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1446" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20174" />
                    <RANKING order="2" place="2" resultid="20729" />
                    <RANKING order="3" place="3" resultid="20287" />
                    <RANKING order="4" place="4" resultid="21873" />
                    <RANKING order="5" place="5" resultid="20291" />
                    <RANKING order="6" place="6" resultid="21594" />
                    <RANKING order="7" place="7" resultid="21880" />
                    <RANKING order="8" place="8" resultid="19976" />
                    <RANKING order="9" place="-1" resultid="21479" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1447" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21101" />
                    <RANKING order="2" place="2" resultid="20911" />
                    <RANKING order="3" place="3" resultid="21141" />
                    <RANKING order="4" place="4" resultid="21356" />
                    <RANKING order="5" place="5" resultid="20926" />
                    <RANKING order="6" place="6" resultid="19812" />
                    <RANKING order="7" place="7" resultid="20228" />
                    <RANKING order="8" place="-1" resultid="19983" />
                    <RANKING order="9" place="-1" resultid="20933" />
                    <RANKING order="10" place="-1" resultid="21194" />
                    <RANKING order="11" place="-1" resultid="21575" />
                    <RANKING order="12" place="-1" resultid="22878" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1448" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20279" />
                    <RANKING order="2" place="2" resultid="21346" />
                    <RANKING order="3" place="3" resultid="20472" />
                    <RANKING order="4" place="4" resultid="22270" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1449" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22004" />
                    <RANKING order="2" place="2" resultid="19861" />
                    <RANKING order="3" place="3" resultid="21266" />
                    <RANKING order="4" place="4" resultid="21625" />
                    <RANKING order="5" place="5" resultid="22396" />
                    <RANKING order="6" place="6" resultid="20464" />
                    <RANKING order="7" place="-1" resultid="22308" />
                    <RANKING order="8" place="-1" resultid="21523" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1450" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21845" />
                    <RANKING order="2" place="2" resultid="21974" />
                    <RANKING order="3" place="3" resultid="20493" />
                    <RANKING order="4" place="4" resultid="19948" />
                    <RANKING order="5" place="-1" resultid="20424" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1451" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19876" />
                    <RANKING order="2" place="2" resultid="19933" />
                    <RANKING order="3" place="3" resultid="21136" />
                    <RANKING order="4" place="-1" resultid="19917" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1452" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22627" />
                    <RANKING order="2" place="2" resultid="21638" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1453" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22653" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1454" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1455" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1456" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24390" daytime="16:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24391" daytime="16:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24392" daytime="16:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24393" daytime="16:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="24394" daytime="16:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="24395" daytime="16:45" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="24396" daytime="16:45" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="24397" daytime="16:50" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="24398" daytime="16:50" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2019-06-02" daytime="09:00" endtime="13:21" name="BLOK IV" number="4" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="1613" daytime="09:10" gender="M" number="33" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1614" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22965" />
                    <RANKING order="2" place="2" resultid="23383" />
                    <RANKING order="3" place="3" resultid="20310" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1615" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22053" />
                    <RANKING order="2" place="2" resultid="22671" />
                    <RANKING order="3" place="3" resultid="20434" />
                    <RANKING order="4" place="4" resultid="21888" />
                    <RANKING order="5" place="5" resultid="21285" />
                    <RANKING order="6" place="6" resultid="20477" />
                    <RANKING order="7" place="7" resultid="20305" />
                    <RANKING order="8" place="-1" resultid="21934" />
                    <RANKING order="9" place="-1" resultid="22661" />
                    <RANKING order="10" place="-1" resultid="23360" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1616" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21923" />
                    <RANKING order="2" place="2" resultid="21727" />
                    <RANKING order="3" place="3" resultid="23000" />
                    <RANKING order="4" place="-1" resultid="22412" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1617" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="23009" />
                    <RANKING order="2" place="2" resultid="21161" />
                    <RANKING order="3" place="3" resultid="22360" />
                    <RANKING order="4" place="-1" resultid="22080" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1618" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20687" />
                    <RANKING order="2" place="2" resultid="22326" />
                    <RANKING order="3" place="3" resultid="21582" />
                    <RANKING order="4" place="4" resultid="22939" />
                    <RANKING order="5" place="5" resultid="22073" />
                    <RANKING order="6" place="6" resultid="20953" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1619" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20176" />
                    <RANKING order="2" place="2" resultid="22035" />
                    <RANKING order="3" place="3" resultid="21875" />
                    <RANKING order="4" place="4" resultid="20292" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1620" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20913" />
                    <RANKING order="2" place="2" resultid="21985" />
                    <RANKING order="3" place="3" resultid="20927" />
                    <RANKING order="4" place="4" resultid="19985" />
                    <RANKING order="5" place="5" resultid="19818" />
                    <RANKING order="6" place="6" resultid="20230" />
                    <RANKING order="7" place="-1" resultid="19813" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1621" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20281" />
                    <RANKING order="2" place="2" resultid="22272" />
                    <RANKING order="3" place="-1" resultid="20920" />
                    <RANKING order="4" place="-1" resultid="21348" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1622" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22005" />
                    <RANKING order="2" place="2" resultid="21267" />
                    <RANKING order="3" place="3" resultid="20465" />
                    <RANKING order="4" place="-1" resultid="21525" />
                    <RANKING order="5" place="-1" resultid="21155" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1623" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21846" />
                    <RANKING order="2" place="2" resultid="20146" />
                    <RANKING order="3" place="3" resultid="21976" />
                    <RANKING order="4" place="-1" resultid="20495" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1624" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21137" />
                    <RANKING order="2" place="2" resultid="21330" />
                    <RANKING order="3" place="3" resultid="20390" />
                    <RANKING order="4" place="4" resultid="20137" />
                    <RANKING order="5" place="5" resultid="20519" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1625" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22629" />
                    <RANKING order="2" place="-1" resultid="20154" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1626" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="22655" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1627" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1628" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1629" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24437" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24438" daytime="09:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24439" daytime="09:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24440" daytime="09:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="24441" daytime="09:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="24442" daytime="09:20" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1647" daytime="09:40" gender="M" number="35" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1648" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21957" />
                    <RANKING order="2" place="2" resultid="21563" />
                    <RANKING order="3" place="3" resultid="23389" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1649" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21545" />
                    <RANKING order="2" place="2" resultid="22054" />
                    <RANKING order="3" place="3" resultid="22977" />
                    <RANKING order="4" place="4" resultid="20190" />
                    <RANKING order="5" place="5" resultid="21667" />
                    <RANKING order="6" place="-1" resultid="22685" />
                    <RANKING order="7" place="-1" resultid="23078" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1650" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22613" />
                    <RANKING order="2" place="2" resultid="22248" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1651" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="23010" />
                    <RANKING order="2" place="2" resultid="21162" />
                    <RANKING order="3" place="3" resultid="20510" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1652" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22344" />
                    <RANKING order="2" place="2" resultid="21583" />
                    <RANKING order="3" place="3" resultid="20199" />
                    <RANKING order="4" place="4" resultid="21860" />
                    <RANKING order="5" place="5" resultid="21394" />
                    <RANKING order="6" place="-1" resultid="20114" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1653" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20731" />
                    <RANKING order="2" place="2" resultid="20177" />
                    <RANKING order="3" place="3" resultid="19970" />
                    <RANKING order="4" place="4" resultid="21832" />
                    <RANKING order="5" place="5" resultid="21405" />
                    <RANKING order="6" place="6" resultid="21308" />
                    <RANKING order="7" place="7" resultid="22044" />
                    <RANKING order="8" place="8" resultid="21481" />
                    <RANKING order="9" place="-1" resultid="20418" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1654" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20242" />
                    <RANKING order="2" place="2" resultid="21237" />
                    <RANKING order="3" place="3" resultid="21986" />
                    <RANKING order="4" place="4" resultid="20256" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1655" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21259" />
                    <RANKING order="2" place="2" resultid="20183" />
                    <RANKING order="3" place="3" resultid="20406" />
                    <RANKING order="4" place="-1" resultid="19807" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1656" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21472" />
                    <RANKING order="2" place="2" resultid="20695" />
                    <RANKING order="3" place="3" resultid="20458" />
                    <RANKING order="4" place="4" resultid="21836" />
                    <RANKING order="5" place="-1" resultid="19863" />
                    <RANKING order="6" place="-1" resultid="21125" />
                    <RANKING order="7" place="-1" resultid="22310" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1657" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22454" />
                    <RANKING order="2" place="2" resultid="20147" />
                    <RANKING order="3" place="3" resultid="23433" />
                    <RANKING order="4" place="4" resultid="21977" />
                    <RANKING order="5" place="-1" resultid="20965" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1658" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21109" />
                    <RANKING order="2" place="2" resultid="19880" />
                    <RANKING order="3" place="3" resultid="20265" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1659" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21464" />
                    <RANKING order="2" place="2" resultid="22429" />
                    <RANKING order="3" place="3" resultid="20943" />
                    <RANKING order="4" place="4" resultid="19942" />
                    <RANKING order="5" place="5" resultid="20442" />
                    <RANKING order="6" place="6" resultid="20128" />
                    <RANKING order="7" place="-1" resultid="20155" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1660" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21991" />
                    <RANKING order="2" place="2" resultid="22420" />
                    <RANKING order="3" place="-1" resultid="20894" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1661" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1662" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1663" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24446" daytime="09:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24447" daytime="09:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24448" daytime="09:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24449" daytime="09:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="24450" daytime="10:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="24451" daytime="10:05" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="24452" daytime="10:10" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1595" daytime="09:00" gender="F" number="32" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1597" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21294" />
                    <RANKING order="2" place="2" resultid="20770" />
                    <RANKING order="3" place="3" resultid="22365" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1598" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22060" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1599" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22015" />
                    <RANKING order="2" place="2" resultid="21744" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1600" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="1601" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20248" />
                    <RANKING order="2" place="2" resultid="21412" />
                    <RANKING order="3" place="3" resultid="21147" />
                    <RANKING order="4" place="4" resultid="21275" />
                    <RANKING order="5" place="-1" resultid="21758" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1602" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21131" />
                    <RANKING order="2" place="2" resultid="21313" />
                    <RANKING order="3" place="3" resultid="21366" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1603" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20207" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1604" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21321" />
                    <RANKING order="2" place="2" resultid="21339" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1605" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21382" />
                    <RANKING order="2" place="2" resultid="21619" />
                    <RANKING order="3" place="3" resultid="20721" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1606" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1607" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1608" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19896" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1609" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1610" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1611" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1612" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24434" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24435" daytime="09:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24436" daytime="09:05" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="19754" daytime="11:30" gender="M" number="40" order="10" round="FHT" preveventid="1744">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="24482" daytime="11:30" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1630" daytime="09:25" gender="F" number="34" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1631" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21559" />
                    <RANKING order="2" place="2" resultid="22921" />
                    <RANKING order="3" place="3" resultid="22366" />
                    <RANKING order="4" place="4" resultid="23395" />
                    <RANKING order="5" place="-1" resultid="23070" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1632" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22021" />
                    <RANKING order="2" place="2" resultid="21554" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1633" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22503" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1634" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20650" />
                    <RANKING order="2" place="2" resultid="22885" />
                    <RANKING order="3" place="-1" resultid="21765" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1635" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22259" />
                    <RANKING order="2" place="2" resultid="21824" />
                    <RANKING order="3" place="3" resultid="22028" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1636" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21174" />
                    <RANKING order="2" place="2" resultid="21735" />
                    <RANKING order="3" place="3" resultid="20221" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1637" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20397" />
                    <RANKING order="2" place="2" resultid="22292" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1638" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21867" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1639" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21519" />
                    <RANKING order="2" place="2" resultid="20412" />
                    <RANKING order="3" place="3" resultid="20487" />
                    <RANKING order="4" place="-1" resultid="19913" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1640" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19872" />
                    <RANKING order="2" place="2" resultid="21489" />
                    <RANKING order="3" place="3" resultid="21634" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1641" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20121" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1642" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1643" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1644" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1645" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1646" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24443" daytime="09:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24444" daytime="09:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24445" daytime="09:35" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1744" daytime="11:35" gender="M" number="40" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="24563" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="23384" />
                    <RANKING order="2" place="2" resultid="21432" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24564" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21286" />
                    <RANKING order="2" place="2" resultid="20478" />
                    <RANKING order="3" place="3" resultid="22971" />
                    <RANKING order="4" place="4" resultid="21668" />
                    <RANKING order="5" place="5" resultid="20191" />
                    <RANKING order="6" place="6" resultid="20636" />
                    <RANKING order="7" place="-1" resultid="21889" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24565" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21504" />
                    <RANKING order="2" place="2" resultid="21709" />
                    <RANKING order="3" place="3" resultid="20503" />
                    <RANKING order="4" place="4" resultid="22464" />
                    <RANKING order="5" place="5" resultid="22413" />
                    <RANKING order="6" place="-1" resultid="21728" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24566" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22336" />
                    <RANKING order="2" place="2" resultid="20511" />
                    <RANKING order="3" place="3" resultid="22361" />
                    <RANKING order="4" place="4" resultid="19783" />
                    <RANKING order="5" place="5" resultid="20237" />
                    <RANKING order="6" place="6" resultid="20629" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24567" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20688" />
                    <RANKING order="2" place="2" resultid="22074" />
                    <RANKING order="3" place="3" resultid="22480" />
                    <RANKING order="4" place="4" resultid="22327" />
                    <RANKING order="5" place="5" resultid="21854" />
                    <RANKING order="6" place="6" resultid="21602" />
                    <RANKING order="7" place="-1" resultid="22492" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24568" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22036" />
                    <RANKING order="2" place="2" resultid="20905" />
                    <RANKING order="3" place="3" resultid="20419" />
                    <RANKING order="4" place="4" resultid="21596" />
                    <RANKING order="5" place="5" resultid="21833" />
                    <RANKING order="6" place="6" resultid="22045" />
                    <RANKING order="7" place="7" resultid="21482" />
                    <RANKING order="8" place="8" resultid="19979" />
                    <RANKING order="9" place="9" resultid="22407" />
                    <RANKING order="10" place="-1" resultid="20273" />
                    <RANKING order="11" place="-1" resultid="21221" />
                    <RANKING order="12" place="-1" resultid="21406" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24569" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22880" />
                    <RANKING order="2" place="2" resultid="22374" />
                    <RANKING order="3" place="3" resultid="20914" />
                    <RANKING order="4" place="4" resultid="21358" />
                    <RANKING order="5" place="5" resultid="20935" />
                    <RANKING order="6" place="6" resultid="19986" />
                    <RANKING order="7" place="7" resultid="20928" />
                    <RANKING order="8" place="8" resultid="22386" />
                    <RANKING order="9" place="9" resultid="21676" />
                    <RANKING order="10" place="10" resultid="23859" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24570" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20474" />
                    <RANKING order="2" place="2" resultid="22066" />
                    <RANKING order="3" place="3" resultid="20407" />
                    <RANKING order="4" place="4" resultid="20921" />
                    <RANKING order="5" place="-1" resultid="19808" />
                    <RANKING order="6" place="-1" resultid="20184" />
                    <RANKING order="7" place="-1" resultid="22273" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24571" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21126" />
                    <RANKING order="2" place="2" resultid="21531" />
                    <RANKING order="3" place="3" resultid="20696" />
                    <RANKING order="4" place="4" resultid="21627" />
                    <RANKING order="5" place="5" resultid="22398" />
                    <RANKING order="6" place="6" resultid="21837" />
                    <RANKING order="7" place="7" resultid="22311" />
                    <RANKING order="8" place="-1" resultid="21473" />
                    <RANKING order="9" place="-1" resultid="21526" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24572" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20496" />
                    <RANKING order="2" place="2" resultid="23434" />
                    <RANKING order="3" place="3" resultid="19778" />
                    <RANKING order="4" place="4" resultid="19950" />
                    <RANKING order="5" place="-1" resultid="20966" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24573" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21331" />
                    <RANKING order="2" place="2" resultid="20162" />
                    <RANKING order="3" place="3" resultid="20391" />
                    <RANKING order="4" place="4" resultid="20520" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24574" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22630" />
                    <RANKING order="2" place="2" resultid="22430" />
                    <RANKING order="3" place="3" resultid="19943" />
                    <RANKING order="4" place="4" resultid="21374" />
                    <RANKING order="5" place="-1" resultid="20129" />
                    <RANKING order="6" place="-1" resultid="20944" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24575" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="24576" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21500" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24577" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="24578" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24474" daytime="11:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24475" daytime="11:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24476" daytime="11:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24477" daytime="12:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="24478" daytime="12:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="24479" daytime="12:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="24480" daytime="12:25" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="24481" daytime="12:30" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1681" daytime="10:25" gender="M" number="37" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1682" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21431" />
                    <RANKING order="2" place="2" resultid="21439" />
                    <RANKING order="3" place="3" resultid="20971" />
                    <RANKING order="4" place="-1" resultid="23402" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1683" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21434" />
                    <RANKING order="2" place="2" resultid="22621" />
                    <RANKING order="3" place="3" resultid="21570" />
                    <RANKING order="4" place="4" resultid="22686" />
                    <RANKING order="5" place="-1" resultid="21549" />
                    <RANKING order="6" place="-1" resultid="23079" />
                    <RANKING order="7" place="-1" resultid="23361" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1684" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21705" />
                    <RANKING order="2" place="2" resultid="20502" />
                    <RANKING order="3" place="-1" resultid="22265" />
                    <RANKING order="4" place="-1" resultid="23001" />
                    <RANKING order="5" place="-1" resultid="23089" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1685" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22335" />
                    <RANKING order="2" place="2" resultid="22087" />
                    <RANKING order="3" place="3" resultid="20236" />
                    <RANKING order="4" place="4" resultid="20628" />
                    <RANKING order="5" place="-1" resultid="22081" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1686" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21455" />
                    <RANKING order="2" place="2" resultid="22476" />
                    <RANKING order="3" place="3" resultid="21853" />
                    <RANKING order="4" place="4" resultid="20200" />
                    <RANKING order="5" place="5" resultid="22345" />
                    <RANKING order="6" place="6" resultid="21681" />
                    <RANKING order="7" place="7" resultid="22254" />
                    <RANKING order="8" place="8" resultid="21391" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1687" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20904" />
                    <RANKING order="2" place="2" resultid="22959" />
                    <RANKING order="3" place="3" resultid="21419" />
                    <RANKING order="4" place="4" resultid="22406" />
                    <RANKING order="5" place="5" resultid="19978" />
                    <RANKING order="6" place="6" resultid="21714" />
                    <RANKING order="7" place="7" resultid="21881" />
                    <RANKING order="8" place="8" resultid="21185" />
                    <RANKING order="9" place="-1" resultid="20272" />
                    <RANKING order="10" place="-1" resultid="21309" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1688" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21576" />
                    <RANKING order="2" place="2" resultid="21102" />
                    <RANKING order="3" place="3" resultid="21238" />
                    <RANKING order="4" place="4" resultid="21195" />
                    <RANKING order="5" place="5" resultid="21357" />
                    <RANKING order="6" place="6" resultid="21675" />
                    <RANKING order="7" place="7" resultid="22385" />
                    <RANKING order="8" place="8" resultid="23858" />
                    <RANKING order="9" place="9" resultid="20231" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1689" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22469" />
                    <RANKING order="2" place="2" resultid="20282" />
                    <RANKING order="3" place="3" resultid="21349" />
                    <RANKING order="4" place="4" resultid="22316" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1690" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22000" />
                    <RANKING order="2" place="2" resultid="23412" />
                    <RANKING order="3" place="3" resultid="22449" />
                    <RANKING order="4" place="4" resultid="21269" />
                    <RANKING order="5" place="5" resultid="19799" />
                    <RANKING order="6" place="6" resultid="21245" />
                    <RANKING order="7" place="-1" resultid="21156" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1691" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22436" />
                    <RANKING order="2" place="2" resultid="20886" />
                    <RANKING order="3" place="3" resultid="20425" />
                    <RANKING order="4" place="4" resultid="19777" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1692" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21110" />
                    <RANKING order="2" place="2" resultid="19934" />
                    <RANKING order="3" place="3" resultid="20138" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1693" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19890" />
                    <RANKING order="2" place="2" resultid="20443" />
                    <RANKING order="3" place="3" resultid="21373" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1694" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20895" />
                    <RANKING order="2" place="2" resultid="21992" />
                    <RANKING order="3" place="3" resultid="22421" />
                    <RANKING order="4" place="-1" resultid="22656" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1695" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20705" />
                    <RANKING order="2" place="2" resultid="21499" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1696" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1697" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24459" daytime="10:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24460" daytime="10:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24461" daytime="10:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24462" daytime="10:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="24463" daytime="10:30" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="24464" daytime="10:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="24465" daytime="10:35" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="24466" daytime="10:35" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1664" daytime="10:10" gender="F" number="36" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1665" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22301" />
                    <RANKING order="2" place="2" resultid="20771" />
                    <RANKING order="3" place="3" resultid="21295" />
                    <RANKING order="4" place="4" resultid="21446" />
                    <RANKING order="5" place="5" resultid="20756" />
                    <RANKING order="6" place="-1" resultid="23071" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1666" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21205" />
                    <RANKING order="2" place="2" resultid="21901" />
                    <RANKING order="3" place="3" resultid="23424" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1667" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22991" />
                    <RANKING order="2" place="2" resultid="21927" />
                    <RANKING order="3" place="3" resultid="20642" />
                    <RANKING order="4" place="4" resultid="21911" />
                    <RANKING order="5" place="5" resultid="21996" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1668" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20957" />
                    <RANKING order="2" place="-1" resultid="21766" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1669" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20249" />
                    <RANKING order="2" place="2" resultid="21180" />
                    <RANKING order="3" place="3" resultid="19792" />
                    <RANKING order="4" place="4" resultid="22954" />
                    <RANKING order="5" place="5" resultid="21759" />
                    <RANKING order="6" place="6" resultid="21276" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1670" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19903" />
                    <RANKING order="2" place="2" resultid="22376" />
                    <RANKING order="3" place="3" resultid="21689" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1671" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21302" />
                    <RANKING order="2" place="2" resultid="20208" />
                    <RANKING order="3" place="3" resultid="23085" />
                    <RANKING order="4" place="4" resultid="22904" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1672" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22485" />
                    <RANKING order="2" place="2" resultid="21117" />
                    <RANKING order="3" place="-1" resultid="23375" />
                    <RANKING order="4" place="-1" resultid="23408" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1673" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22285" />
                    <RANKING order="2" place="2" resultid="22635" />
                    <RANKING order="3" place="3" resultid="21383" />
                    <RANKING order="4" place="4" resultid="21611" />
                    <RANKING order="5" place="5" resultid="21620" />
                    <RANKING order="6" place="6" resultid="20712" />
                    <RANKING order="7" place="7" resultid="22909" />
                    <RANKING order="8" place="8" resultid="23857" />
                    <RANKING order="9" place="-1" resultid="19866" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1674" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22280" />
                    <RANKING order="2" place="2" resultid="19842" />
                    <RANKING order="3" place="3" resultid="19856" />
                    <RANKING order="4" place="4" resultid="20450" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1675" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19920" />
                    <RANKING order="2" place="2" resultid="21231" />
                    <RANKING order="3" place="3" resultid="20122" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1676" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19897" />
                    <RANKING order="2" place="2" resultid="21226" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1677" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20430" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1678" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1679" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1680" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24453" daytime="10:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24454" daytime="10:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24455" daytime="10:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24456" daytime="10:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="24457" daytime="10:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="24458" daytime="10:20" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="19753" daytime="10:45" gender="F" number="39" order="8" round="FHT" preveventid="1721">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="24473" daytime="10:45" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1721" daytime="10:50" gender="F" number="39" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="24547" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22302" />
                    <RANKING order="2" place="2" resultid="20757" />
                    <RANKING order="3" place="3" resultid="20762" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24548" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21588" />
                    <RANKING order="2" place="2" resultid="22061" />
                    <RANKING order="3" place="3" resultid="22022" />
                    <RANKING order="4" place="4" resultid="23425" />
                    <RANKING order="5" place="5" resultid="22640" />
                    <RANKING order="6" place="-1" resultid="21190" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24549" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22992" />
                    <RANKING order="2" place="2" resultid="22016" />
                    <RANKING order="3" place="3" resultid="24645" />
                    <RANKING order="4" place="4" resultid="20643" />
                    <RANKING order="5" place="-1" resultid="21745" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24550" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22497" />
                    <RANKING order="2" place="2" resultid="20651" />
                    <RANKING order="3" place="3" resultid="24644" />
                    <RANKING order="4" place="4" resultid="22926" />
                    <RANKING order="5" place="-1" resultid="22886" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24551" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20261" />
                    <RANKING order="2" place="2" resultid="19793" />
                    <RANKING order="3" place="3" resultid="21413" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24552" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19904" />
                    <RANKING order="2" place="2" resultid="21752" />
                    <RANKING order="3" place="3" resultid="20222" />
                    <RANKING order="4" place="4" resultid="21736" />
                    <RANKING order="5" place="5" resultid="21690" />
                    <RANKING order="6" place="6" resultid="21367" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24553" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20398" />
                    <RANKING order="2" place="2" resultid="22293" />
                    <RANKING order="3" place="3" resultid="23086" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24554" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21322" />
                    <RANKING order="2" place="2" resultid="21868" />
                    <RANKING order="3" place="3" resultid="21340" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24555" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21520" />
                    <RANKING order="2" place="2" resultid="21612" />
                    <RANKING order="3" place="3" resultid="19914" />
                    <RANKING order="4" place="4" resultid="20488" />
                    <RANKING order="5" place="5" resultid="20713" />
                    <RANKING order="6" place="-1" resultid="20722" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24556" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21490" />
                    <RANKING order="2" place="2" resultid="19843" />
                    <RANKING order="3" place="-1" resultid="22697" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24557" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22439" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24558" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="24559" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="24560" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="24561" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="24562" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24469" daytime="10:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24470" daytime="11:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="24471" daytime="11:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="24472" daytime="11:20" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1698" daytime="10:35" gender="X" number="38" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="16674" agemax="99" agemin="80" calculate="TOTAL" />
                <AGEGROUP agegroupid="16675" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21565" />
                    <RANKING order="2" place="2" resultid="22092" />
                    <RANKING order="3" place="-1" resultid="21960" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16676" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="20656" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16677" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="22093" />
                    <RANKING order="2" place="2" resultid="21213" />
                    <RANKING order="3" place="3" resultid="22514" />
                    <RANKING order="4" place="4" resultid="21893" />
                    <RANKING order="5" place="5" resultid="22978" />
                    <RANKING order="6" place="-1" resultid="23376" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16678" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21215" />
                    <RANKING order="2" place="2" resultid="22372" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16679" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="21396" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16680" agemax="-1" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="19926" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24467" daytime="10:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="24468" daytime="10:40" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" nation="POL" clubid="23057" name="3Waters Akademia Sportów Wodnych">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1975-08-09" firstname="Sonia" gender="F" lastname="Borkowska" nation="POL" athleteid="23058">
              <RESULTS>
                <RESULT eventid="1062" points="367" reactiontime="+75" swimtime="00:00:33.05" resultid="23059" heatid="24279" lane="3" entrytime="00:00:32.80" />
                <RESULT eventid="1256" points="305" swimtime="00:01:16.81" resultid="23061" heatid="24351" lane="6" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="WAR" clubid="21597" name="5Styl Warszawa">
          <CONTACT name="Korzeniowski" />
          <ATHLETES>
            <ATHLETE birthdate="1977-06-16" firstname="Adrian" gender="M" lastname="Kulisz" nation="POL" athleteid="21598">
              <RESULTS>
                <RESULT eventid="1079" points="285" reactiontime="+110" swimtime="00:00:31.75" resultid="21599" heatid="24288" lane="2" entrytime="00:00:31.70" />
                <RESULT eventid="1273" points="286" swimtime="00:01:11.15" resultid="21600" heatid="24359" lane="9" entrytime="00:01:09.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="268" swimtime="00:02:38.20" resultid="21601" heatid="24420" lane="9" entrytime="00:02:37.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.29" />
                    <SPLIT distance="150" swimtime="00:01:57.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="259" reactiontime="+70" swimtime="00:05:44.99" resultid="21602" heatid="24478" lane="2" entrytime="00:05:56.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.33" />
                    <SPLIT distance="100" swimtime="00:01:21.29" />
                    <SPLIT distance="150" swimtime="00:02:04.94" />
                    <SPLIT distance="200" swimtime="00:02:50.20" />
                    <SPLIT distance="250" swimtime="00:03:34.66" />
                    <SPLIT distance="350" swimtime="00:05:03.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="23064" name="Akademia WSB">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1996-03-24" firstname="Kinga" gender="F" lastname="Pluta" nation="POL" athleteid="23065">
              <RESULTS>
                <RESULT eventid="1222" points="351" swimtime="00:03:17.06" resultid="23066" heatid="24340" lane="9" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.00" />
                    <SPLIT distance="100" swimtime="00:01:32.98" />
                    <SPLIT distance="150" swimtime="00:02:25.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="411" reactiontime="+85" swimtime="00:01:09.54" resultid="23067" heatid="24350" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="374" swimtime="00:01:28.98" resultid="23068" heatid="24378" lane="9" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" status="DNS" swimtime="00:00:00.00" resultid="23069" heatid="24387" lane="0" entrytime="00:00:45.00" />
                <RESULT eventid="1630" status="DNS" swimtime="00:00:00.00" resultid="23070" heatid="24444" lane="8" entrytime="00:03:20.00" />
                <RESULT eventid="1664" status="DNS" swimtime="00:00:00.00" resultid="23071" heatid="24456" lane="5" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="22610" name="Aqua Fit Środa Śląska">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1985-07-05" firstname="Sebastian" gender="M" lastname="Figarski" nation="POL" athleteid="22611">
              <RESULTS>
                <RESULT eventid="1474" points="503" reactiontime="+71" swimtime="00:01:05.19" resultid="22612" heatid="24408" lane="7" entrytime="00:01:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="464" reactiontime="+68" swimtime="00:02:24.53" resultid="22613" heatid="24452" lane="7" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                    <SPLIT distance="100" swimtime="00:01:09.81" />
                    <SPLIT distance="150" swimtime="00:01:47.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="22007" name="AQUASFERA Masters Olsztyn">
          <CONTACT name="Goździejewska Anna" />
          <ATHLETES>
            <ATHLETE birthdate="1993-06-11" firstname="Zuzanna" gender="F" lastname="Brzozowska" nation="POL" athleteid="22017">
              <RESULTS>
                <RESULT eventid="1147" points="443" reactiontime="+76" swimtime="00:10:35.94" resultid="22018" heatid="24312" lane="7" entrytime="00:10:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                    <SPLIT distance="100" swimtime="00:01:14.08" />
                    <SPLIT distance="150" swimtime="00:01:53.99" />
                    <SPLIT distance="200" swimtime="00:02:34.31" />
                    <SPLIT distance="250" swimtime="00:03:14.36" />
                    <SPLIT distance="300" swimtime="00:03:54.95" />
                    <SPLIT distance="350" swimtime="00:04:34.77" />
                    <SPLIT distance="400" swimtime="00:05:15.16" />
                    <SPLIT distance="450" swimtime="00:05:55.56" />
                    <SPLIT distance="500" swimtime="00:06:36.18" />
                    <SPLIT distance="550" swimtime="00:07:16.13" />
                    <SPLIT distance="600" swimtime="00:07:56.31" />
                    <SPLIT distance="650" swimtime="00:08:36.75" />
                    <SPLIT distance="700" swimtime="00:09:18.00" />
                    <SPLIT distance="750" swimtime="00:09:57.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="505" swimtime="00:01:04.90" resultid="22019" heatid="24352" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="487" reactiontime="+73" swimtime="00:02:23.55" resultid="22020" heatid="24414" lane="8" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="100" swimtime="00:01:08.57" />
                    <SPLIT distance="150" swimtime="00:01:46.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="428" reactiontime="+68" swimtime="00:02:44.52" resultid="22021" heatid="24445" lane="7" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.02" />
                    <SPLIT distance="100" swimtime="00:01:19.04" />
                    <SPLIT distance="150" swimtime="00:02:02.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="409" reactiontime="+49" swimtime="00:05:18.45" resultid="22022" heatid="24473" lane="6" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                    <SPLIT distance="100" swimtime="00:01:16.67" />
                    <SPLIT distance="150" swimtime="00:01:57.36" />
                    <SPLIT distance="200" swimtime="00:02:38.48" />
                    <SPLIT distance="250" swimtime="00:03:18.80" />
                    <SPLIT distance="300" swimtime="00:03:59.54" />
                    <SPLIT distance="350" swimtime="00:04:39.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-10-26" firstname="Joanna" gender="F" lastname="Drzewicka" nation="POL" athleteid="22023">
              <RESULTS>
                <RESULT eventid="1062" points="329" reactiontime="+82" swimtime="00:00:34.28" resultid="22024" heatid="24278" lane="7" entrytime="00:00:36.55" />
                <RESULT eventid="1187" points="399" swimtime="00:00:36.75" resultid="22025" heatid="24325" lane="4" entrytime="00:00:40.04" />
                <RESULT eventid="1256" points="275" reactiontime="+42" swimtime="00:01:19.46" resultid="22026" heatid="24350" lane="1" entrytime="00:01:25.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="329" reactiontime="+91" swimtime="00:01:23.95" resultid="22027" heatid="24401" lane="0" entrytime="00:01:30.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="242" reactiontime="+85" swimtime="00:03:18.95" resultid="22028" heatid="24443" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-30" firstname="Paweł" gender="M" lastname="Gregorowicz" nation="POL" athleteid="22029">
              <RESULTS>
                <RESULT eventid="1079" points="471" reactiontime="+70" swimtime="00:00:26.87" resultid="22030" heatid="24291" lane="9" entrytime="00:00:29.50" />
                <RESULT eventid="14189" points="481" reactiontime="+82" swimtime="00:09:36.96" resultid="22031" heatid="24317" lane="3" entrytime="00:09:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                    <SPLIT distance="100" swimtime="00:01:07.88" />
                    <SPLIT distance="150" swimtime="00:01:43.56" />
                    <SPLIT distance="200" swimtime="00:02:20.29" />
                    <SPLIT distance="250" swimtime="00:02:56.44" />
                    <SPLIT distance="300" swimtime="00:03:33.20" />
                    <SPLIT distance="350" swimtime="00:04:09.79" />
                    <SPLIT distance="400" swimtime="00:04:46.57" />
                    <SPLIT distance="450" swimtime="00:05:23.04" />
                    <SPLIT distance="500" swimtime="00:06:00.03" />
                    <SPLIT distance="550" swimtime="00:06:36.66" />
                    <SPLIT distance="600" swimtime="00:07:13.17" />
                    <SPLIT distance="650" swimtime="00:07:49.60" />
                    <SPLIT distance="700" swimtime="00:08:26.05" />
                    <SPLIT distance="750" swimtime="00:09:02.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="517" reactiontime="+69" swimtime="00:00:58.44" resultid="22032" heatid="24363" lane="4" entrytime="00:00:58.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="458" swimtime="00:02:12.29" resultid="22033" heatid="24424" lane="0" entrytime="00:02:07.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.64" />
                    <SPLIT distance="100" swimtime="00:01:03.98" />
                    <SPLIT distance="150" swimtime="00:01:38.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="429" swimtime="00:05:23.28" resultid="22034" heatid="24433" lane="9" entrytime="00:05:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                    <SPLIT distance="100" swimtime="00:01:09.97" />
                    <SPLIT distance="200" swimtime="00:02:39.26" />
                    <SPLIT distance="250" swimtime="00:03:25.43" />
                    <SPLIT distance="300" swimtime="00:04:11.27" />
                    <SPLIT distance="350" swimtime="00:04:47.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="479" reactiontime="+69" swimtime="00:01:03.67" resultid="22035" heatid="24441" lane="7" entrytime="00:01:05.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="501" reactiontime="+72" swimtime="00:04:37.08" resultid="22036" heatid="24482" lane="2" entrytime="00:04:38.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.78" />
                    <SPLIT distance="100" swimtime="00:01:06.46" />
                    <SPLIT distance="150" swimtime="00:01:41.50" />
                    <SPLIT distance="200" swimtime="00:02:17.07" />
                    <SPLIT distance="250" swimtime="00:02:52.48" />
                    <SPLIT distance="300" swimtime="00:03:28.42" />
                    <SPLIT distance="350" swimtime="00:04:03.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-06-13" firstname="Michał" gender="M" lastname="Kieres" nation="POL" athleteid="22075">
              <RESULTS>
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="22076" heatid="24345" lane="2" entrytime="00:02:59.00" />
                <RESULT eventid="1341" status="DNS" swimtime="00:00:00.00" resultid="22077" heatid="24370" lane="3" entrytime="00:02:50.00" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="22078" heatid="24384" lane="0" entrytime="00:01:21.00" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="22079" heatid="24393" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="22080" heatid="24440" lane="6" entrytime="00:01:10.00" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="22081" heatid="24464" lane="5" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-04-01" firstname="Piotr" gender="M" lastname="Konopacki" nation="POL" athleteid="22067">
              <RESULTS>
                <RESULT eventid="1079" points="416" reactiontime="+93" swimtime="00:00:28.01" resultid="22068" heatid="24292" lane="4" entrytime="00:00:27.99" />
                <RESULT eventid="14207" points="417" reactiontime="+71" swimtime="00:19:25.21" resultid="22069" heatid="24322" lane="7" entrytime="00:20:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.87" />
                    <SPLIT distance="100" swimtime="00:01:12.67" />
                    <SPLIT distance="150" swimtime="00:01:52.05" />
                    <SPLIT distance="200" swimtime="00:02:31.93" />
                    <SPLIT distance="250" swimtime="00:03:12.08" />
                    <SPLIT distance="300" swimtime="00:03:52.48" />
                    <SPLIT distance="350" swimtime="00:04:32.09" />
                    <SPLIT distance="400" swimtime="00:05:12.16" />
                    <SPLIT distance="450" swimtime="00:05:51.74" />
                    <SPLIT distance="500" swimtime="00:06:31.26" />
                    <SPLIT distance="550" swimtime="00:07:10.66" />
                    <SPLIT distance="600" swimtime="00:07:50.04" />
                    <SPLIT distance="650" swimtime="00:08:29.43" />
                    <SPLIT distance="700" swimtime="00:09:08.86" />
                    <SPLIT distance="750" swimtime="00:09:47.86" />
                    <SPLIT distance="800" swimtime="00:10:27.05" />
                    <SPLIT distance="850" swimtime="00:11:06.05" />
                    <SPLIT distance="900" swimtime="00:11:44.70" />
                    <SPLIT distance="950" swimtime="00:12:23.49" />
                    <SPLIT distance="1000" swimtime="00:13:02.39" />
                    <SPLIT distance="1050" swimtime="00:13:41.25" />
                    <SPLIT distance="1100" swimtime="00:14:20.43" />
                    <SPLIT distance="1150" swimtime="00:14:59.15" />
                    <SPLIT distance="1200" swimtime="00:15:38.38" />
                    <SPLIT distance="1250" swimtime="00:16:16.90" />
                    <SPLIT distance="1300" swimtime="00:16:56.16" />
                    <SPLIT distance="1350" swimtime="00:17:34.40" />
                    <SPLIT distance="1400" swimtime="00:18:12.18" />
                    <SPLIT distance="1450" swimtime="00:18:49.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="451" swimtime="00:01:01.15" resultid="22070" heatid="24362" lane="9" entrytime="00:01:02.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="433" reactiontime="+71" swimtime="00:02:14.81" resultid="22071" heatid="24422" lane="7" entrytime="00:02:18.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.42" />
                    <SPLIT distance="100" swimtime="00:01:05.03" />
                    <SPLIT distance="150" swimtime="00:01:40.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="383" swimtime="00:05:35.70" resultid="22072" heatid="24432" lane="6" entrytime="00:05:48.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                    <SPLIT distance="100" swimtime="00:01:19.72" />
                    <SPLIT distance="150" swimtime="00:02:05.68" />
                    <SPLIT distance="200" swimtime="00:02:48.82" />
                    <SPLIT distance="250" swimtime="00:03:37.99" />
                    <SPLIT distance="300" swimtime="00:04:26.17" />
                    <SPLIT distance="350" swimtime="00:05:02.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="322" swimtime="00:01:12.65" resultid="22073" heatid="24440" lane="9" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="440" swimtime="00:04:49.34" resultid="22074" heatid="24481" lane="6" entrytime="00:04:53.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.61" />
                    <SPLIT distance="100" swimtime="00:01:09.29" />
                    <SPLIT distance="150" swimtime="00:01:46.23" />
                    <SPLIT distance="200" swimtime="00:02:23.85" />
                    <SPLIT distance="250" swimtime="00:03:00.65" />
                    <SPLIT distance="300" swimtime="00:03:38.63" />
                    <SPLIT distance="350" swimtime="00:04:15.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-15" firstname="Michał" gender="M" lastname="Kozikowski" nation="POL" athleteid="22082">
              <RESULTS>
                <RESULT eventid="1079" points="430" reactiontime="+77" swimtime="00:00:27.70" resultid="22083" heatid="24292" lane="6" entrytime="00:00:28.00" />
                <RESULT eventid="1239" points="406" swimtime="00:02:50.96" resultid="22084" heatid="24346" lane="0" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.10" />
                    <SPLIT distance="100" swimtime="00:01:22.56" />
                    <SPLIT distance="150" swimtime="00:02:06.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="390" reactiontime="+72" swimtime="00:01:18.15" resultid="22085" heatid="24384" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="303" reactiontime="+71" swimtime="00:06:02.77" resultid="22086" heatid="24432" lane="2" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.89" />
                    <SPLIT distance="100" swimtime="00:01:27.57" />
                    <SPLIT distance="150" swimtime="00:02:14.46" />
                    <SPLIT distance="200" swimtime="00:02:59.85" />
                    <SPLIT distance="250" swimtime="00:03:47.75" />
                    <SPLIT distance="300" swimtime="00:04:35.14" />
                    <SPLIT distance="350" swimtime="00:05:19.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="449" reactiontime="+51" swimtime="00:00:33.87" resultid="22087" heatid="24465" lane="7" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-03-19" firstname="Oriana" gender="F" lastname="Lewandowska" nation="POL" athleteid="22055">
              <RESULTS>
                <RESULT eventid="1147" points="500" reactiontime="+95" swimtime="00:10:10.76" resultid="22056" heatid="24312" lane="4" entrytime="00:10:20.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                    <SPLIT distance="100" swimtime="00:01:14.42" />
                    <SPLIT distance="150" swimtime="00:01:54.08" />
                    <SPLIT distance="200" swimtime="00:02:33.21" />
                    <SPLIT distance="250" swimtime="00:03:12.00" />
                    <SPLIT distance="300" swimtime="00:03:50.81" />
                    <SPLIT distance="350" swimtime="00:04:29.19" />
                    <SPLIT distance="400" swimtime="00:05:07.78" />
                    <SPLIT distance="450" swimtime="00:05:45.69" />
                    <SPLIT distance="500" swimtime="00:06:24.07" />
                    <SPLIT distance="550" swimtime="00:07:02.35" />
                    <SPLIT distance="600" swimtime="00:07:41.26" />
                    <SPLIT distance="650" swimtime="00:08:19.36" />
                    <SPLIT distance="700" swimtime="00:08:57.33" />
                    <SPLIT distance="750" swimtime="00:09:34.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="529" reactiontime="+91" swimtime="00:02:30.53" resultid="22057" heatid="24367" lane="4" entrytime="00:02:40.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                    <SPLIT distance="100" swimtime="00:01:11.48" />
                    <SPLIT distance="150" swimtime="00:01:51.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="464" reactiontime="+81" swimtime="00:00:31.55" resultid="22058" heatid="24389" lane="6" entrytime="00:00:31.00" />
                <RESULT eventid="1491" points="473" reactiontime="+88" swimtime="00:02:24.92" resultid="22059" heatid="24414" lane="1" entrytime="00:02:24.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.60" />
                    <SPLIT distance="100" swimtime="00:01:10.51" />
                    <SPLIT distance="150" swimtime="00:01:48.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="492" reactiontime="+87" swimtime="00:01:10.24" resultid="22060" heatid="24436" lane="6" entrytime="00:01:11.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="463" reactiontime="+93" swimtime="00:05:05.51" resultid="22061" heatid="24473" lane="2" entrytime="00:05:01.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                    <SPLIT distance="100" swimtime="00:01:15.45" />
                    <SPLIT distance="150" swimtime="00:03:12.48" />
                    <SPLIT distance="200" swimtime="00:02:34.18" />
                    <SPLIT distance="300" swimtime="00:03:50.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-06-25" firstname="Adam" gender="M" lastname="Matusiak vel Matuszewski" nation="POL" athleteid="22037">
              <RESULTS>
                <RESULT eventid="1079" points="226" reactiontime="+81" swimtime="00:00:34.30" resultid="22038" heatid="24286" lane="8" entrytime="00:00:35.11" />
                <RESULT eventid="14189" points="260" reactiontime="+105" swimtime="00:11:47.93" resultid="22039" heatid="24316" lane="1" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.40" />
                    <SPLIT distance="200" swimtime="00:02:50.14" />
                    <SPLIT distance="250" swimtime="00:03:35.30" />
                    <SPLIT distance="300" swimtime="00:04:20.39" />
                    <SPLIT distance="350" swimtime="00:05:05.54" />
                    <SPLIT distance="400" swimtime="00:05:49.99" />
                    <SPLIT distance="450" swimtime="00:06:35.17" />
                    <SPLIT distance="500" swimtime="00:07:19.96" />
                    <SPLIT distance="550" swimtime="00:08:04.98" />
                    <SPLIT distance="600" swimtime="00:08:49.60" />
                    <SPLIT distance="700" swimtime="00:10:19.24" />
                    <SPLIT distance="750" swimtime="00:11:03.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="184" swimtime="00:00:42.13" resultid="22040" heatid="24331" lane="2" entrytime="00:00:43.49" />
                <RESULT eventid="1273" points="246" swimtime="00:01:14.83" resultid="22041" heatid="24357" lane="8" entrytime="00:01:18.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="182" swimtime="00:01:31.40" resultid="22042" heatid="24404" lane="5" entrytime="00:01:37.99" />
                <RESULT eventid="1508" points="249" reactiontime="+42" swimtime="00:02:41.97" resultid="22043" heatid="24419" lane="1" entrytime="00:02:48.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.67" />
                    <SPLIT distance="100" swimtime="00:01:19.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="183" reactiontime="+82" swimtime="00:03:17.12" resultid="22044" heatid="24448" lane="2" entrytime="00:03:40.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.95" />
                    <SPLIT distance="100" swimtime="00:01:37.50" />
                    <SPLIT distance="150" swimtime="00:02:30.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="256" swimtime="00:05:46.20" resultid="22045" heatid="24478" lane="1" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.67" />
                    <SPLIT distance="100" swimtime="00:01:22.05" />
                    <SPLIT distance="150" swimtime="00:02:06.31" />
                    <SPLIT distance="200" swimtime="00:02:50.69" />
                    <SPLIT distance="250" swimtime="00:03:35.23" />
                    <SPLIT distance="300" swimtime="00:04:19.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-09-15" firstname="Mieszko" gender="M" lastname="Palmi-Kukiełko" nation="POL" athleteid="22046">
              <RESULTS>
                <RESULT eventid="1113" points="625" reactiontime="+76" swimtime="00:02:13.30" resultid="22047" heatid="24307" lane="4" entrytime="00:02:14.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.96" />
                    <SPLIT distance="100" swimtime="00:01:00.89" />
                    <SPLIT distance="150" swimtime="00:01:40.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14207" points="539" reactiontime="+78" swimtime="00:17:50.24" resultid="22048" heatid="24322" lane="5" entrytime="00:18:03.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.97" />
                    <SPLIT distance="100" swimtime="00:01:03.50" />
                    <SPLIT distance="150" swimtime="00:01:38.19" />
                    <SPLIT distance="200" swimtime="00:02:13.45" />
                    <SPLIT distance="250" swimtime="00:02:49.05" />
                    <SPLIT distance="300" swimtime="00:03:25.32" />
                    <SPLIT distance="350" swimtime="00:04:01.88" />
                    <SPLIT distance="400" swimtime="00:04:38.22" />
                    <SPLIT distance="450" swimtime="00:05:14.78" />
                    <SPLIT distance="500" swimtime="00:05:51.84" />
                    <SPLIT distance="550" swimtime="00:06:28.48" />
                    <SPLIT distance="600" swimtime="00:07:04.92" />
                    <SPLIT distance="650" swimtime="00:07:40.87" />
                    <SPLIT distance="700" swimtime="00:08:17.23" />
                    <SPLIT distance="750" swimtime="00:08:53.29" />
                    <SPLIT distance="800" swimtime="00:09:29.71" />
                    <SPLIT distance="850" swimtime="00:10:05.99" />
                    <SPLIT distance="900" swimtime="00:10:42.44" />
                    <SPLIT distance="950" swimtime="00:11:18.38" />
                    <SPLIT distance="1000" swimtime="00:11:54.86" />
                    <SPLIT distance="1050" swimtime="00:12:30.82" />
                    <SPLIT distance="1100" swimtime="00:13:07.17" />
                    <SPLIT distance="1150" swimtime="00:13:43.05" />
                    <SPLIT distance="1200" swimtime="00:14:19.31" />
                    <SPLIT distance="1250" swimtime="00:14:55.15" />
                    <SPLIT distance="1300" swimtime="00:15:31.42" />
                    <SPLIT distance="1350" swimtime="00:16:06.60" />
                    <SPLIT distance="1400" swimtime="00:16:42.59" />
                    <SPLIT distance="1450" swimtime="00:17:16.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="594" swimtime="00:00:28.54" resultid="22049" heatid="24336" lane="3" entrytime="00:00:27.49" />
                <RESULT eventid="1341" points="548" reactiontime="+67" swimtime="00:02:16.20" resultid="22050" heatid="24371" lane="4" entrytime="00:02:14.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.53" />
                    <SPLIT distance="100" swimtime="00:01:02.19" />
                    <SPLIT distance="150" swimtime="00:01:37.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="585" swimtime="00:02:01.91" resultid="22051" heatid="24424" lane="5" entrytime="00:01:57.74">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.57" />
                    <SPLIT distance="150" swimtime="00:01:30.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="568" swimtime="00:04:54.27" resultid="22052" heatid="24433" lane="4" entrytime="00:04:51.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.93" />
                    <SPLIT distance="100" swimtime="00:01:03.21" />
                    <SPLIT distance="150" swimtime="00:01:43.14" />
                    <SPLIT distance="200" swimtime="00:02:22.74" />
                    <SPLIT distance="250" swimtime="00:03:05.73" />
                    <SPLIT distance="300" swimtime="00:03:48.35" />
                    <SPLIT distance="350" swimtime="00:04:21.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="656" swimtime="00:00:57.32" resultid="22053" heatid="24442" lane="4" entrytime="00:00:57.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="528" swimtime="00:02:18.42" resultid="22054" heatid="24452" lane="5" entrytime="00:02:14.89">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-09-15" firstname="Adam" gender="M" lastname="Szmit" nation="POL" athleteid="22062">
              <RESULTS>
                <RESULT eventid="14207" points="279" reactiontime="+100" swimtime="00:22:12.25" resultid="22063" heatid="24322" lane="9" entrytime="00:22:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                    <SPLIT distance="100" swimtime="00:01:19.96" />
                    <SPLIT distance="150" swimtime="00:03:31.78" />
                    <SPLIT distance="200" swimtime="00:05:44.81" />
                    <SPLIT distance="250" swimtime="00:09:26.05" />
                    <SPLIT distance="350" swimtime="00:10:54.81" />
                    <SPLIT distance="450" swimtime="00:12:24.74" />
                    <SPLIT distance="500" swimtime="00:11:40.85" />
                    <SPLIT distance="550" swimtime="00:16:57.43" />
                    <SPLIT distance="600" swimtime="00:16:11.36" />
                    <SPLIT distance="650" swimtime="00:21:29.68" />
                    <SPLIT distance="700" swimtime="00:20:42.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="270" reactiontime="+103" swimtime="00:01:12.56" resultid="22064" heatid="24358" lane="8" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="266" reactiontime="+64" swimtime="00:02:38.59" resultid="22065" heatid="24419" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.27" />
                    <SPLIT distance="100" swimtime="00:01:16.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="289" reactiontime="+91" swimtime="00:05:32.60" resultid="22066" heatid="24479" lane="8" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                    <SPLIT distance="150" swimtime="00:02:00.90" />
                    <SPLIT distance="300" swimtime="00:05:32.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-17" firstname="Anna" gender="F" lastname="Zaleska" nation="POL" athleteid="22008">
              <RESULTS>
                <RESULT eventid="1096" points="364" reactiontime="+93" swimtime="00:02:56.61" resultid="22009" heatid="24298" lane="7" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.92" />
                    <SPLIT distance="100" swimtime="00:01:21.85" />
                    <SPLIT distance="150" swimtime="00:02:15.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="331" reactiontime="+87" swimtime="00:11:40.80" resultid="22010" heatid="24312" lane="9" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.77" />
                    <SPLIT distance="100" swimtime="00:01:20.10" />
                    <SPLIT distance="150" swimtime="00:02:04.11" />
                    <SPLIT distance="200" swimtime="00:02:48.13" />
                    <SPLIT distance="250" swimtime="00:03:32.50" />
                    <SPLIT distance="300" swimtime="00:04:16.60" />
                    <SPLIT distance="350" swimtime="00:05:00.91" />
                    <SPLIT distance="400" swimtime="00:05:45.68" />
                    <SPLIT distance="450" swimtime="00:06:30.36" />
                    <SPLIT distance="500" swimtime="00:07:14.45" />
                    <SPLIT distance="550" swimtime="00:07:59.19" />
                    <SPLIT distance="600" swimtime="00:08:44.03" />
                    <SPLIT distance="650" swimtime="00:09:28.86" />
                    <SPLIT distance="700" swimtime="00:10:13.77" />
                    <SPLIT distance="750" swimtime="00:10:57.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="357" swimtime="00:00:38.12" resultid="22011" heatid="24326" lane="1" entrytime="00:00:39.00" />
                <RESULT eventid="1324" points="376" reactiontime="+87" swimtime="00:02:48.67" resultid="22012" heatid="24367" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                    <SPLIT distance="100" swimtime="00:01:20.90" />
                    <SPLIT distance="150" swimtime="00:02:04.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="355" reactiontime="+48" swimtime="00:00:34.50" resultid="22013" heatid="24388" lane="7" entrytime="00:00:35.50" />
                <RESULT eventid="1555" points="345" reactiontime="+63" swimtime="00:06:19.77" resultid="22014" heatid="24429" lane="5" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="200" swimtime="00:03:02.98" />
                    <SPLIT distance="300" swimtime="00:04:51.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="361" reactiontime="+80" swimtime="00:01:17.91" resultid="22015" heatid="24436" lane="7" entrytime="00:01:17.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="354" reactiontime="+84" swimtime="00:05:33.97" resultid="22016" heatid="24471" lane="6" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.50" />
                    <SPLIT distance="100" swimtime="00:01:20.73" />
                    <SPLIT distance="150" swimtime="00:02:03.92" />
                    <SPLIT distance="200" swimtime="00:02:47.72" />
                    <SPLIT distance="250" swimtime="00:03:29.81" />
                    <SPLIT distance="300" swimtime="00:04:12.74" />
                    <SPLIT distance="350" swimtime="00:04:53.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="GENTELMEN" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="481" reactiontime="+67" swimtime="00:01:59.22" resultid="22095" heatid="24374" lane="2" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.88" />
                    <SPLIT distance="100" swimtime="00:01:03.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22046" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="22082" number="2" />
                    <RELAYPOSITION athleteid="22029" number="3" reactiontime="+5" />
                    <RELAYPOSITION athleteid="22067" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" name="WŚCIEKŁY PIES" number="1">
              <RESULTS>
                <RESULT eventid="1548" points="497" swimtime="00:01:47.09" resultid="22091" heatid="24427" lane="2" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.48" />
                    <SPLIT distance="100" swimtime="00:00:54.87" />
                    <SPLIT distance="150" swimtime="00:01:21.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22029" number="1" />
                    <RELAYPOSITION athleteid="22082" number="2" />
                    <RELAYPOSITION athleteid="22067" number="3" />
                    <RELAYPOSITION athleteid="22046" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="LEJDIS" number="1">
              <RESULTS>
                <RESULT eventid="1358" points="427" reactiontime="+75" swimtime="00:02:21.18" resultid="22089" heatid="24372" lane="6" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.64" />
                    <SPLIT distance="100" swimtime="00:01:19.82" />
                    <SPLIT distance="150" swimtime="00:01:52.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22023" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="22008" number="2" />
                    <RELAYPOSITION athleteid="22055" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="22017" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" name="PINA COLADA" number="1">
              <RESULTS>
                <RESULT eventid="1525" points="427" reactiontime="+80" swimtime="00:02:08.07" resultid="22090" heatid="24425" lane="6" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                    <SPLIT distance="100" swimtime="00:01:00.97" />
                    <SPLIT distance="150" swimtime="00:01:34.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22055" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="22017" number="2" />
                    <RELAYPOSITION athleteid="22008" number="3" reactiontime="+4" />
                    <RELAYPOSITION athleteid="22023" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" name="KAMIKAZE" number="1">
              <RESULTS>
                <RESULT eventid="1698" reactiontime="+116" swimtime="00:02:04.34" resultid="22092" heatid="24468" lane="4" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.44" />
                    <SPLIT distance="100" swimtime="00:01:03.00" />
                    <SPLIT distance="150" swimtime="00:01:35.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22046" number="1" reactiontime="+116" />
                    <RELAYPOSITION athleteid="22082" number="2" />
                    <RELAYPOSITION athleteid="22055" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="22017" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="MOJITO" number="1">
              <RESULTS>
                <RESULT eventid="1698" reactiontime="+78" swimtime="00:02:12.56" resultid="22093" heatid="24468" lane="7" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.04" />
                    <SPLIT distance="100" swimtime="00:01:11.47" />
                    <SPLIT distance="150" swimtime="00:01:45.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22023" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="22029" number="2" />
                    <RELAYPOSITION athleteid="22008" number="3" reactiontime="+23" />
                    <RELAYPOSITION athleteid="22067" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="SŁODZIAKI" number="1">
              <RESULTS>
                <RESULT eventid="1130" reactiontime="+70" swimtime="00:02:01.13" resultid="22088" heatid="24309" lane="8" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.47" />
                    <SPLIT distance="100" swimtime="00:00:54.63" />
                    <SPLIT distance="150" swimtime="00:01:27.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22029" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="22067" number="2" />
                    <RELAYPOSITION athleteid="22008" number="3" reactiontime="+30" />
                    <RELAYPOSITION athleteid="22023" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" name="ŚWIERZAKI" number="1">
              <RESULTS>
                <RESULT eventid="1130" reactiontime="+78" swimtime="00:01:54.34" resultid="22094" heatid="24309" lane="5" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.01" />
                    <SPLIT distance="100" swimtime="00:00:54.88" />
                    <SPLIT distance="150" swimtime="00:01:25.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22046" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="22082" number="2" />
                    <RELAYPOSITION athleteid="22055" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="22017" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="POM" clubid="21447" name="AquaStars Gdynia">
          <CONTACT email="mariuszgolon5@wp.pl" name="GOLON" phone="609649755" />
          <ATHLETES>
            <ATHLETE birthdate="1978-11-20" firstname="Mariusz" gender="M" lastname="Golon" nation="POL" athleteid="21448">
              <RESULTS>
                <RESULT eventid="1079" points="403" reactiontime="+88" swimtime="00:00:28.30" resultid="21449" heatid="24290" lane="0" entrytime="00:00:30.00" />
                <RESULT eventid="1113" points="265" reactiontime="+89" swimtime="00:02:57.43" resultid="21450" heatid="24305" lane="9" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.20" />
                    <SPLIT distance="100" swimtime="00:01:19.57" />
                    <SPLIT distance="150" swimtime="00:02:15.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="351" swimtime="00:00:34.01" resultid="21451" heatid="24330" lane="5" entrytime="00:00:45.00" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="21452" heatid="24344" lane="8" entrytime="00:03:15.00" />
                <RESULT eventid="1406" points="339" reactiontime="+47" swimtime="00:01:21.84" resultid="21453" heatid="24381" lane="2" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="437" swimtime="00:00:29.33" resultid="21454" heatid="24395" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="1681" points="411" swimtime="00:00:34.90" resultid="21455" heatid="24464" lane="8" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00611" nation="POL" region="SLA" clubid="21491" name="AZS AWF Katowice">
          <CONTACT city="Katowice" email="m.skora@awf.katowice.pl" name="Michał Skóra" phone="501370222" state="ŚLĄSK" street="Mikołowska 72a" zip="40-065" />
          <ATHLETES>
            <ATHLETE birthdate="1986-10-19" firstname="Michał" gender="M" lastname="Skrodzki" nation="POL" athleteid="21501">
              <RESULTS>
                <RESULT eventid="14207" points="470" reactiontime="+86" swimtime="00:18:39.63" resultid="21502" heatid="24322" lane="6" entrytime="00:18:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                    <SPLIT distance="100" swimtime="00:01:08.26" />
                    <SPLIT distance="150" swimtime="00:01:44.89" />
                    <SPLIT distance="200" swimtime="00:02:22.00" />
                    <SPLIT distance="250" swimtime="00:02:59.25" />
                    <SPLIT distance="300" swimtime="00:03:36.46" />
                    <SPLIT distance="350" swimtime="00:04:14.25" />
                    <SPLIT distance="400" swimtime="00:04:51.31" />
                    <SPLIT distance="450" swimtime="00:05:28.93" />
                    <SPLIT distance="500" swimtime="00:06:06.12" />
                    <SPLIT distance="550" swimtime="00:06:43.91" />
                    <SPLIT distance="600" swimtime="00:07:21.44" />
                    <SPLIT distance="650" swimtime="00:07:59.58" />
                    <SPLIT distance="700" swimtime="00:08:36.87" />
                    <SPLIT distance="750" swimtime="00:09:14.78" />
                    <SPLIT distance="800" swimtime="00:09:53.10" />
                    <SPLIT distance="850" swimtime="00:10:31.16" />
                    <SPLIT distance="900" swimtime="00:11:08.79" />
                    <SPLIT distance="950" swimtime="00:11:46.76" />
                    <SPLIT distance="1000" swimtime="00:12:24.21" />
                    <SPLIT distance="1050" swimtime="00:13:02.23" />
                    <SPLIT distance="1100" swimtime="00:13:39.86" />
                    <SPLIT distance="1150" swimtime="00:14:17.97" />
                    <SPLIT distance="1200" swimtime="00:14:55.30" />
                    <SPLIT distance="1250" swimtime="00:15:33.24" />
                    <SPLIT distance="1300" swimtime="00:16:11.27" />
                    <SPLIT distance="1350" swimtime="00:16:49.43" />
                    <SPLIT distance="1400" swimtime="00:17:27.11" />
                    <SPLIT distance="1450" swimtime="00:18:04.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="488" swimtime="00:02:09.48" resultid="21503" heatid="24423" lane="1" entrytime="00:02:12.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.20" />
                    <SPLIT distance="100" swimtime="00:01:03.07" />
                    <SPLIT distance="150" swimtime="00:01:36.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="479" reactiontime="+77" swimtime="00:04:41.11" resultid="21504" heatid="24482" lane="7" entrytime="00:04:40.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.92" />
                    <SPLIT distance="100" swimtime="00:01:05.91" />
                    <SPLIT distance="150" swimtime="00:01:41.31" />
                    <SPLIT distance="200" swimtime="00:02:17.57" />
                    <SPLIT distance="250" swimtime="00:02:53.58" />
                    <SPLIT distance="300" swimtime="00:03:29.99" />
                    <SPLIT distance="350" swimtime="00:04:05.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1931-04-27" firstname="Jan" gender="M" lastname="Ślężyński" nation="POL" license="100611700315" athleteid="21492">
              <RESULTS>
                <RESULT eventid="1079" points="38" reactiontime="+96" swimtime="00:01:02.11" resultid="21493" heatid="24283" lane="2" entrytime="00:00:58.48" />
                <RESULT eventid="14207" points="28" reactiontime="+118" swimtime="00:47:15.25" resultid="21494" heatid="24320" lane="0" entrytime="00:44:33.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.79" />
                    <SPLIT distance="100" swimtime="00:02:50.49" />
                    <SPLIT distance="150" swimtime="00:04:23.38" />
                    <SPLIT distance="200" swimtime="00:05:55.19" />
                    <SPLIT distance="250" swimtime="00:07:29.99" />
                    <SPLIT distance="300" swimtime="00:09:03.30" />
                    <SPLIT distance="350" swimtime="00:10:36.86" />
                    <SPLIT distance="400" swimtime="00:12:11.71" />
                    <SPLIT distance="450" swimtime="00:13:47.10" />
                    <SPLIT distance="500" swimtime="00:15:20.83" />
                    <SPLIT distance="550" swimtime="00:16:56.94" />
                    <SPLIT distance="600" swimtime="00:18:29.72" />
                    <SPLIT distance="650" swimtime="00:20:05.29" />
                    <SPLIT distance="700" swimtime="00:21:39.89" />
                    <SPLIT distance="750" swimtime="00:23:16.22" />
                    <SPLIT distance="800" swimtime="00:24:52.96" />
                    <SPLIT distance="850" swimtime="00:26:29.09" />
                    <SPLIT distance="900" swimtime="00:28:06.98" />
                    <SPLIT distance="950" swimtime="00:29:41.27" />
                    <SPLIT distance="1000" swimtime="00:31:18.57" />
                    <SPLIT distance="1050" swimtime="00:32:51.99" />
                    <SPLIT distance="1100" swimtime="00:34:28.66" />
                    <SPLIT distance="1150" swimtime="00:36:07.88" />
                    <SPLIT distance="1200" swimtime="00:36:59.93" />
                    <SPLIT distance="1250" swimtime="00:39:20.21" />
                    <SPLIT distance="1300" swimtime="00:37:43.71" />
                    <SPLIT distance="1350" swimtime="00:42:33.47" />
                    <SPLIT distance="1400" swimtime="00:44:08.39" />
                    <SPLIT distance="1450" swimtime="00:45:40.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="37" reactiontime="+47" swimtime="00:06:17.12" resultid="21495" heatid="24341" lane="3" entrytime="00:05:52.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.70" />
                    <SPLIT distance="100" swimtime="00:03:04.64" />
                    <SPLIT distance="150" swimtime="00:04:43.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="29" reactiontime="+95" swimtime="00:02:31.59" resultid="21496" heatid="24355" lane="8" entrytime="00:02:32.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="31" reactiontime="+78" swimtime="00:03:01.74" resultid="21497" heatid="24380" lane="6" entrytime="00:02:43.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="29" reactiontime="+44" swimtime="00:05:31.58" resultid="21498" heatid="24416" lane="7" entrytime="00:05:15.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.55" />
                    <SPLIT distance="100" swimtime="00:02:44.47" />
                    <SPLIT distance="150" swimtime="00:04:14.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="34" reactiontime="+49" swimtime="00:01:19.93" resultid="21499" heatid="24460" lane="0" entrytime="00:01:08.57" />
                <RESULT eventid="1744" points="30" reactiontime="+57" swimtime="00:11:46.03" resultid="21500" heatid="24475" lane="0" entrytime="00:10:21.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.06" />
                    <SPLIT distance="100" swimtime="00:02:56.11" />
                    <SPLIT distance="150" swimtime="00:04:28.31" />
                    <SPLIT distance="200" swimtime="00:05:58.26" />
                    <SPLIT distance="250" swimtime="00:07:28.90" />
                    <SPLIT distance="300" swimtime="00:08:58.50" />
                    <SPLIT distance="350" swimtime="00:10:27.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="SLA" clubid="21539" name="BAZA PŁYWANIA Mysłowice">
          <CONTACT city="Mysłowice" email="adrian,kisiel93@gmail.com" name="Kisiel" phone="502593038" state="ŚLĄSK" zip="41-400" />
          <ATHLETES>
            <ATHLETE birthdate="1994-06-16" firstname="Paulina" gender="F" lastname="Dąbrowska" nation="POL" athleteid="21550">
              <RESULTS>
                <RESULT eventid="1062" points="443" reactiontime="+86" swimtime="00:00:31.05" resultid="21551" heatid="24281" lane="8" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT eventid="1187" points="431" swimtime="00:00:35.80" resultid="21552" heatid="24327" lane="2" entrytime="00:00:34.00" entrycourse="LCM" />
                <RESULT eventid="1457" points="410" reactiontime="+76" swimtime="00:01:18.05" resultid="21553" heatid="24402" lane="3" entrytime="00:01:12.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="393" reactiontime="+83" swimtime="00:02:49.36" resultid="21554" heatid="24445" lane="3" entrytime="00:02:38.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.41" />
                    <SPLIT distance="100" swimtime="00:01:22.29" />
                    <SPLIT distance="150" swimtime="00:02:06.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-05-20" firstname="Rafał" gender="M" lastname="Handzlik" nation="POL" athleteid="21560">
              <RESULTS>
                <RESULT eventid="1205" points="539" reactiontime="+59" swimtime="00:00:29.49" resultid="21561" heatid="24336" lane="7" entrytime="00:00:28.00" entrycourse="LCM" />
                <RESULT eventid="1273" points="492" swimtime="00:00:59.41" resultid="21562" heatid="24364" lane="0" entrytime="00:00:58.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="462" reactiontime="+56" swimtime="00:02:24.76" resultid="21563" heatid="24452" lane="3" entrytime="00:02:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                    <SPLIT distance="100" swimtime="00:01:09.91" />
                    <SPLIT distance="150" swimtime="00:01:48.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-03-26" firstname="Adrian" gender="M" lastname="Kisiel" nation="POL" athleteid="21540">
              <RESULTS>
                <RESULT eventid="1079" points="616" reactiontime="+73" swimtime="00:00:24.57" resultid="21541" heatid="24296" lane="2" entrytime="00:00:24.50" entrycourse="LCM" />
                <RESULT eventid="1205" points="620" reactiontime="+74" swimtime="00:00:28.14" resultid="21542" heatid="24336" lane="2" entrytime="00:00:27.50" entrycourse="LCM" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="21543" heatid="24398" lane="1" entrytime="00:00:26.00" entrycourse="LCM" />
                <RESULT eventid="1474" points="592" reactiontime="+69" swimtime="00:01:01.74" resultid="21544" heatid="24408" lane="3" entrytime="00:00:59.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="544" swimtime="00:02:17.10" resultid="21545" heatid="24452" lane="6" entrytime="00:02:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                    <SPLIT distance="100" swimtime="00:01:07.45" />
                    <SPLIT distance="150" swimtime="00:01:43.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-05-27" firstname="Monika" gender="F" lastname="Kisiel" nation="POL" athleteid="21555">
              <RESULTS>
                <RESULT eventid="1187" points="493" swimtime="00:00:34.24" resultid="21556" heatid="24327" lane="3" entrytime="00:00:33.50" entrycourse="LCM" />
                <RESULT eventid="1457" points="472" swimtime="00:01:14.45" resultid="21557" heatid="24402" lane="5" entrytime="00:01:12.00" entrycourse="LCM" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="21558" heatid="24413" lane="5" entrytime="00:02:32.00" entrycourse="LCM" />
                <RESULT eventid="1630" points="405" swimtime="00:02:47.63" resultid="21559" heatid="24445" lane="5" entrytime="00:02:38.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.70" />
                    <SPLIT distance="100" swimtime="00:01:22.60" />
                    <SPLIT distance="150" swimtime="00:02:05.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-06-29" firstname="Paweł" gender="M" lastname="Trenda" nation="POL" athleteid="21546">
              <RESULTS>
                <RESULT eventid="1205" points="596" reactiontime="+108" swimtime="00:00:28.51" resultid="21547" heatid="24336" lane="4" entrytime="00:00:27.00" entrycourse="LCM" />
                <RESULT eventid="1474" points="547" reactiontime="+64" swimtime="00:01:03.39" resultid="21548" heatid="24408" lane="5" entrytime="00:00:59.00" entrycourse="LCM" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="21549" heatid="24466" lane="8" entrytime="00:00:31.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" reactiontime="+120" swimtime="00:01:51.19" resultid="21564" heatid="24309" lane="2" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.82" />
                    <SPLIT distance="100" swimtime="00:00:56.41" />
                    <SPLIT distance="150" swimtime="00:01:27.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21546" number="1" reactiontime="+120" />
                    <RELAYPOSITION athleteid="21555" number="2" />
                    <RELAYPOSITION athleteid="21550" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="21540" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" reactiontime="+68" swimtime="00:02:00.80" resultid="21565" heatid="24468" lane="3" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                    <SPLIT distance="100" swimtime="00:01:04.41" />
                    <SPLIT distance="150" swimtime="00:01:30.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21555" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="21546" number="2" />
                    <RELAYPOSITION athleteid="21540" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="21550" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="CMUJKR" nation="POL" region="MAL" clubid="21097" name="Collegium Medicum UJ Masters Kraków">
          <CONTACT city="Kraków" email="mariuszbaranik@gmail.com" name="Mariusz Baranik" phone="69812822" state="MAL" street="Białopradnicka 32c/3" zip="31-221" />
          <ATHLETES>
            <ATHLETE birthdate="1969-06-29" firstname="Mariusz" gender="M" lastname="Baranik" nation="POL" athleteid="21098">
              <RESULTS>
                <RESULT eventid="1079" points="434" reactiontime="+79" swimtime="00:00:27.60" resultid="21099" heatid="24293" lane="7" entrytime="00:00:27.40" />
                <RESULT eventid="1273" points="424" swimtime="00:01:02.42" resultid="21100" heatid="24362" lane="1" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="427" reactiontime="+70" swimtime="00:00:29.57" resultid="21101" heatid="24396" lane="8" entrytime="00:00:29.40" />
                <RESULT eventid="1681" points="382" reactiontime="+78" swimtime="00:00:35.75" resultid="21102" heatid="24464" lane="3" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-03-25" firstname="Jacek" gender="M" lastname="Kwiatkowski" nation="POL" athleteid="22675">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="22676" heatid="24287" lane="4" entrytime="00:00:32.30" />
                <RESULT eventid="14207" points="195" swimtime="00:25:00.47" resultid="22677" heatid="24321" lane="8" entrytime="00:25:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.44" />
                    <SPLIT distance="100" swimtime="00:01:32.04" />
                    <SPLIT distance="150" swimtime="00:02:20.80" />
                    <SPLIT distance="200" swimtime="00:03:10.69" />
                    <SPLIT distance="250" swimtime="00:04:00.35" />
                    <SPLIT distance="300" swimtime="00:04:50.65" />
                    <SPLIT distance="350" swimtime="00:05:41.19" />
                    <SPLIT distance="400" swimtime="00:06:32.49" />
                    <SPLIT distance="450" swimtime="00:07:22.86" />
                    <SPLIT distance="500" swimtime="00:08:13.33" />
                    <SPLIT distance="550" swimtime="00:09:04.29" />
                    <SPLIT distance="600" swimtime="00:11:35.52" />
                    <SPLIT distance="650" swimtime="00:10:44.99" />
                    <SPLIT distance="700" swimtime="00:13:16.64" />
                    <SPLIT distance="750" swimtime="00:12:25.91" />
                    <SPLIT distance="800" swimtime="00:14:57.25" />
                    <SPLIT distance="850" swimtime="00:14:07.19" />
                    <SPLIT distance="900" swimtime="00:18:18.94" />
                    <SPLIT distance="950" swimtime="00:17:27.88" />
                    <SPLIT distance="1050" swimtime="00:19:08.84" />
                    <SPLIT distance="1150" swimtime="00:20:49.40" />
                    <SPLIT distance="1200" swimtime="00:19:58.82" />
                    <SPLIT distance="1250" swimtime="00:22:31.85" />
                    <SPLIT distance="1300" swimtime="00:21:40.87" />
                    <SPLIT distance="1400" swimtime="00:23:22.82" />
                    <SPLIT distance="1450" swimtime="00:24:13.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02711" nation="POL" region="SLA" clubid="21641" name="CSiR Dąbrowa Górnicza">
          <CONTACT name="Waliczek" />
          <ATHLETES>
            <ATHLETE birthdate="1997-01-01" firstname="Bernard" gender="M" lastname="Filek" nation="POL" athleteid="23385">
              <RESULTS>
                <RESULT eventid="1205" points="381" reactiontime="+70" swimtime="00:00:33.08" resultid="23386" heatid="24336" lane="0" entrytime="00:00:29.00" />
                <RESULT eventid="1474" points="308" reactiontime="+120" swimtime="00:01:16.73" resultid="23387" heatid="24407" lane="4" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="225" swimtime="00:06:40.86" resultid="23388" heatid="24430" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                    <SPLIT distance="100" swimtime="00:01:20.48" />
                    <SPLIT distance="150" swimtime="00:02:11.76" />
                    <SPLIT distance="200" swimtime="00:03:05.78" />
                    <SPLIT distance="250" swimtime="00:04:06.12" />
                    <SPLIT distance="300" swimtime="00:05:08.00" />
                    <SPLIT distance="350" swimtime="00:05:54.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="273" swimtime="00:02:52.51" resultid="23389" heatid="24451" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                    <SPLIT distance="100" swimtime="00:01:23.31" />
                    <SPLIT distance="150" swimtime="00:02:08.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Bartosz" gender="M" lastname="Katolik" nation="POL" athleteid="23378">
              <RESULTS>
                <RESULT eventid="1079" points="521" reactiontime="+66" swimtime="00:00:25.98" resultid="23379" heatid="24295" lane="6" entrytime="00:00:26.00" />
                <RESULT eventid="1205" points="415" reactiontime="+69" swimtime="00:00:32.17" resultid="23380" heatid="24336" lane="9" entrytime="00:00:29.00" />
                <RESULT eventid="1273" points="505" swimtime="00:00:58.89" resultid="23381" heatid="24363" lane="3" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="518" swimtime="00:00:27.72" resultid="23382" heatid="24397" lane="0" entrytime="00:00:28.50" />
                <RESULT eventid="1613" points="434" swimtime="00:01:05.76" resultid="23383" heatid="24441" lane="1" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="353" swimtime="00:05:11.29" resultid="23384" heatid="24480" lane="6" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                    <SPLIT distance="100" swimtime="00:01:15.13" />
                    <SPLIT distance="150" swimtime="00:01:55.25" />
                    <SPLIT distance="200" swimtime="00:02:34.61" />
                    <SPLIT distance="250" swimtime="00:03:13.09" />
                    <SPLIT distance="300" swimtime="00:03:53.38" />
                    <SPLIT distance="350" swimtime="00:04:33.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-06-01" firstname="Dawid" gender="M" lastname="Nowodworski" nation="POL" athleteid="23396">
              <RESULTS>
                <RESULT eventid="1079" points="628" reactiontime="+71" swimtime="00:00:24.41" resultid="23397" heatid="24296" lane="5" entrytime="00:00:24.00" />
                <RESULT eventid="1205" points="606" swimtime="00:00:28.36" resultid="23398" heatid="24336" lane="6" entrytime="00:00:27.50" />
                <RESULT eventid="1273" points="671" reactiontime="+65" swimtime="00:00:53.58" resultid="23399" heatid="24365" lane="4" entrytime="00:00:53.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="607" swimtime="00:01:07.43" resultid="23400" heatid="24385" lane="7" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="672" reactiontime="+57" swimtime="00:00:25.42" resultid="23401" heatid="24398" lane="4" entrytime="00:00:24.90" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="23402" heatid="24466" lane="5" entrytime="00:00:29.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Wiktoria" gender="F" lastname="Szlachcic" nation="POL" athleteid="23390">
              <RESULTS>
                <RESULT eventid="1062" status="DNS" swimtime="00:00:00.00" resultid="23391" heatid="24280" lane="1" entrytime="00:00:31.50" />
                <RESULT eventid="1187" points="473" swimtime="00:00:34.73" resultid="23392" heatid="24327" lane="1" entrytime="00:00:34.50" />
                <RESULT eventid="1256" points="417" swimtime="00:01:09.19" resultid="23393" heatid="24353" lane="9" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="413" reactiontime="+74" swimtime="00:01:17.86" resultid="23394" heatid="24402" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="363" reactiontime="+118" swimtime="00:02:53.84" resultid="23395" heatid="24445" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.57" />
                    <SPLIT distance="100" swimtime="00:01:22.86" />
                    <SPLIT distance="150" swimtime="00:02:08.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="20435" name="DELFIN92 Gliwice">
          <CONTACT email="cupialsport@op.pl" name="Cupiał" phone="605065587" />
          <ATHLETES>
            <ATHLETE birthdate="1951-01-01" firstname="Teodozja" gender="F" lastname="Gdula" nation="POL" athleteid="20447">
              <RESULTS>
                <RESULT eventid="1222" points="91" reactiontime="+87" swimtime="00:05:08.92" resultid="20448" heatid="24337" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.70" />
                    <SPLIT distance="100" swimtime="00:02:29.26" />
                    <SPLIT distance="150" swimtime="00:03:48.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="78" reactiontime="+92" swimtime="00:02:29.97" resultid="20449" heatid="24375" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="84" reactiontime="+117" swimtime="00:01:07.06" resultid="20450" heatid="24454" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-02-10" firstname="Barbara" gender="F" lastname="Lipowska" nation="POL" athleteid="20444">
              <RESULTS>
                <RESULT eventid="1062" points="89" reactiontime="+94" swimtime="00:00:52.88" resultid="20445" heatid="24276" lane="0" />
                <RESULT eventid="1256" points="59" reactiontime="+100" swimtime="00:02:12.24" resultid="20446" heatid="24348" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-11-23" firstname="Jerzy" gender="M" lastname="Marciniszko" nation="POL" athleteid="20436">
              <RESULTS>
                <RESULT eventid="1079" points="30" reactiontime="+85" swimtime="00:01:07.11" resultid="20437" heatid="24283" lane="7" entrytime="00:01:06.98" />
                <RESULT eventid="1205" points="35" swimtime="00:01:13.09" resultid="20438" heatid="24329" lane="0" entrytime="00:01:04.12" />
                <RESULT eventid="1239" points="58" reactiontime="+75" swimtime="00:05:25.85" resultid="20439" heatid="24341" lane="5" entrytime="00:05:30.81">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:41.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="50" reactiontime="+113" swimtime="00:02:34.95" resultid="20440" heatid="24380" lane="3" entrytime="00:02:26.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="38" reactiontime="+111" swimtime="00:02:32.92" resultid="20441" heatid="24403" lane="2" entrytime="00:02:22.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="30" reactiontime="+104" swimtime="00:05:58.35" resultid="20442" heatid="24447" lane="9" entrytime="00:05:33.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:25.46" />
                    <SPLIT distance="100" swimtime="00:03:01.88" />
                    <SPLIT distance="150" swimtime="00:04:32.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="72" reactiontime="+99" swimtime="00:01:02.25" resultid="20443" heatid="24460" lane="7" entrytime="00:01:00.65" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="23072" name="Dąbrowska Szkoła Pływania">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1993-02-05" firstname="Kacper" gender="M" lastname="Kaproń" nation="POL" athleteid="23073">
              <RESULTS>
                <RESULT eventid="1205" points="241" swimtime="00:00:38.52" resultid="23074" heatid="24331" lane="9" entrytime="00:00:45.00" />
                <RESULT eventid="1239" points="282" reactiontime="+78" swimtime="00:03:13.09" resultid="23075" heatid="24344" lane="3" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.60" />
                    <SPLIT distance="100" swimtime="00:01:29.00" />
                    <SPLIT distance="150" swimtime="00:02:19.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="296" reactiontime="+54" swimtime="00:01:25.62" resultid="23076" heatid="24381" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="23077" heatid="24404" lane="7" entrytime="00:01:45.00" />
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="23078" heatid="24449" lane="9" entrytime="00:03:20.00" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="23079" heatid="24461" lane="8" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="20881" name="Gdynia Masters">
          <CONTACT email="kasiiamysiak@gmail.com" name="Mysiak" />
          <ATHLETES>
            <ATHLETE birthdate="1953-01-01" firstname="Andrzej" gender="M" lastname="Jacaszek" nation="POL" athleteid="20882">
              <RESULTS>
                <RESULT eventid="1079" points="185" reactiontime="+108" swimtime="00:00:36.64" resultid="20883" heatid="24285" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="1239" points="204" reactiontime="+64" swimtime="00:03:35.14" resultid="20884" heatid="24343" lane="6" entrytime="00:03:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.77" />
                    <SPLIT distance="100" swimtime="00:01:41.19" />
                    <SPLIT distance="150" swimtime="00:02:40.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="220" reactiontime="+96" swimtime="00:01:34.48" resultid="20885" heatid="24382" lane="7" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="247" reactiontime="+75" swimtime="00:00:41.32" resultid="20886" heatid="24461" lane="4" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-01-01" firstname="Andrzej" gender="M" lastname="Skwarło" nation="POL" athleteid="20887">
              <RESULTS>
                <RESULT eventid="1079" points="110" reactiontime="+119" swimtime="00:00:43.51" resultid="20888" heatid="24284" lane="1" entrytime="00:00:42.50" />
                <RESULT eventid="1113" points="75" reactiontime="+113" swimtime="00:04:29.71" resultid="20889" heatid="24302" lane="0" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.14" />
                    <SPLIT distance="100" swimtime="00:02:21.58" />
                    <SPLIT distance="150" swimtime="00:03:32.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="91" swimtime="00:00:53.23" resultid="20890" heatid="24330" lane="6" entrytime="00:00:50.00" />
                <RESULT eventid="1239" points="98" reactiontime="+95" swimtime="00:04:34.12" resultid="20891" heatid="24342" lane="2" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.61" />
                    <SPLIT distance="100" swimtime="00:02:12.84" />
                    <SPLIT distance="150" swimtime="00:03:26.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="101" reactiontime="+91" swimtime="00:02:02.52" resultid="20892" heatid="24381" lane="1" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="62" reactiontime="+146" swimtime="00:02:10.72" resultid="20893" heatid="24403" lane="4" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.82" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O2 - Pływak nie miał kontaktu ze ścianą podczas nawrotu. (Time: 10:00)" eventid="1647" status="DSQ" swimtime="00:04:42.71" resultid="20894" heatid="24447" lane="6" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.43" />
                    <SPLIT distance="100" swimtime="00:02:07.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="131" reactiontime="+64" swimtime="00:00:51.01" resultid="20895" heatid="24461" lane="9" entrytime="00:00:48.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="22614" name="GVT Wrocław">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1979-09-26" firstname="Łukasz" gender="M" lastname="Malaczewski" nation="POL" athleteid="22615">
              <RESULTS>
                <RESULT eventid="1079" points="481" reactiontime="+80" swimtime="00:00:26.68" resultid="22616" heatid="24294" lane="2" entrytime="00:00:26.60" />
                <RESULT eventid="1273" points="468" swimtime="00:01:00.38" resultid="22617" heatid="24363" lane="9" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="20906" name="IKS Konstancin">
          <CONTACT email="golyswim@interia.pl" name="golon" phone="601385695" />
          <ATHLETES>
            <ATHLETE birthdate="1969-04-11" firstname="Paweł" gender="M" lastname="Obiedziński" nation="POL" athleteid="20907">
              <RESULTS>
                <RESULT eventid="1079" points="424" reactiontime="+72" swimtime="00:00:27.83" resultid="20908" heatid="24292" lane="8" entrytime="00:00:28.50" entrycourse="LCM" />
                <RESULT eventid="1113" points="321" reactiontime="+82" swimtime="00:02:46.40" resultid="20909" heatid="24305" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.89" />
                    <SPLIT distance="100" swimtime="00:01:19.63" />
                    <SPLIT distance="150" swimtime="00:02:09.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="440" swimtime="00:01:01.67" resultid="20910" heatid="24362" lane="8" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="354" swimtime="00:00:31.47" resultid="20911" heatid="24394" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="1508" points="394" swimtime="00:02:19.02" resultid="20912" heatid="24422" lane="5" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                    <SPLIT distance="100" swimtime="00:01:06.75" />
                    <SPLIT distance="150" swimtime="00:01:43.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="299" reactiontime="+59" swimtime="00:01:14.48" resultid="20913" heatid="24440" lane="8" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="364" swimtime="00:05:08.11" resultid="20914" heatid="24480" lane="1" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                    <SPLIT distance="100" swimtime="00:01:11.68" />
                    <SPLIT distance="150" swimtime="00:01:51.02" />
                    <SPLIT distance="200" swimtime="00:02:30.71" />
                    <SPLIT distance="250" swimtime="00:03:10.87" />
                    <SPLIT distance="300" swimtime="00:03:50.86" />
                    <SPLIT distance="350" swimtime="00:04:30.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-02-23" firstname="Maciej" gender="M" lastname="Piłatowicz" nation="POL" license="103714700120" athleteid="21216">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="21217" heatid="24288" lane="4" entrytime="00:00:31.01" />
                <RESULT eventid="14207" points="248" reactiontime="+96" swimtime="00:23:05.77" resultid="21218" heatid="24321" lane="4" entrytime="00:22:44.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.94" />
                    <SPLIT distance="100" swimtime="00:01:26.25" />
                    <SPLIT distance="150" swimtime="00:02:12.71" />
                    <SPLIT distance="200" swimtime="00:02:59.43" />
                    <SPLIT distance="250" swimtime="00:03:45.31" />
                    <SPLIT distance="300" swimtime="00:04:30.83" />
                    <SPLIT distance="350" swimtime="00:05:16.39" />
                    <SPLIT distance="400" swimtime="00:06:02.28" />
                    <SPLIT distance="450" swimtime="00:06:48.30" />
                    <SPLIT distance="500" swimtime="00:07:34.64" />
                    <SPLIT distance="550" swimtime="00:08:20.81" />
                    <SPLIT distance="600" swimtime="00:09:07.14" />
                    <SPLIT distance="650" swimtime="00:09:53.59" />
                    <SPLIT distance="700" swimtime="00:10:40.04" />
                    <SPLIT distance="750" swimtime="00:11:26.90" />
                    <SPLIT distance="800" swimtime="00:12:13.34" />
                    <SPLIT distance="850" swimtime="00:12:59.94" />
                    <SPLIT distance="900" swimtime="00:13:46.59" />
                    <SPLIT distance="950" swimtime="00:14:33.07" />
                    <SPLIT distance="1000" swimtime="00:15:20.28" />
                    <SPLIT distance="1050" swimtime="00:16:07.11" />
                    <SPLIT distance="1100" swimtime="00:16:54.34" />
                    <SPLIT distance="1150" swimtime="00:17:41.05" />
                    <SPLIT distance="1200" swimtime="00:18:28.01" />
                    <SPLIT distance="1250" swimtime="00:19:14.95" />
                    <SPLIT distance="1300" swimtime="00:20:01.35" />
                    <SPLIT distance="1350" swimtime="00:20:48.42" />
                    <SPLIT distance="1400" swimtime="00:21:34.66" />
                    <SPLIT distance="1450" swimtime="00:22:21.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="21219" heatid="24358" lane="4" entrytime="00:01:09.99" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="21220" heatid="24421" lane="2" entrytime="00:02:29.98" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="21221" heatid="24479" lane="6" entrytime="00:05:34.97" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="PDL" clubid="22929" name="Iswim Białystok">
          <CONTACT email="biuro@isiwm.bialystok.pl" internet="www.iswim.bialystok.pl" name="SEBSTAIN HUMBLA" phone="782997050" street="WIERZBOWA 3" street2="Białystok" />
          <ATHLETES>
            <ATHLETE birthdate="1979-11-12" firstname="Piotr" gender="M" lastname="Buczko" nation="POL" athleteid="22944">
              <RESULTS>
                <RESULT eventid="1079" points="442" reactiontime="+75" swimtime="00:00:27.45" resultid="22945" heatid="24294" lane="8" entrytime="00:00:26.80" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="22946" heatid="24396" lane="0" entrytime="00:00:29.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-12" firstname="Maciej" gender="M" lastname="Daszuta" nation="POL" athleteid="22955">
              <RESULTS>
                <RESULT eventid="1079" points="409" reactiontime="+80" swimtime="00:00:28.16" resultid="22956" heatid="24293" lane="1" entrytime="00:00:27.50" />
                <RESULT eventid="1205" points="383" reactiontime="+68" swimtime="00:00:33.02" resultid="22957" heatid="24334" lane="5" entrytime="00:00:31.90" />
                <RESULT eventid="1406" points="337" swimtime="00:01:22.01" resultid="22958" heatid="24384" lane="5" entrytime="00:01:17.00" />
                <RESULT eventid="1681" points="425" reactiontime="+46" swimtime="00:00:34.49" resultid="22959" heatid="24465" lane="4" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-01" firstname="Justyna" gender="F" lastname="Hermanowicz" nation="POL" athleteid="24643">
              <RESULTS>
                <RESULT eventid="1721" points="230" reactiontime="+85" swimtime="00:06:25.68" resultid="24644" heatid="24469" lane="6" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.45" />
                    <SPLIT distance="100" swimtime="00:01:29.05" />
                    <SPLIT distance="150" swimtime="00:02:16.72" />
                    <SPLIT distance="200" swimtime="00:03:07.07" />
                    <SPLIT distance="250" swimtime="00:03:56.89" />
                    <SPLIT distance="300" swimtime="00:04:47.73" />
                    <SPLIT distance="350" swimtime="00:05:37.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-07-17" firstname="Magda" gender="F" lastname="Iwaniuk Mróż" nation="POL" athleteid="22950">
              <RESULTS>
                <RESULT eventid="1062" points="409" reactiontime="+94" swimtime="00:00:31.87" resultid="22951" heatid="24279" lane="2" entrytime="00:00:32.90" />
                <RESULT eventid="1187" points="313" swimtime="00:00:39.84" resultid="22952" heatid="24326" lane="5" entrytime="00:00:37.20" />
                <RESULT eventid="1388" points="335" reactiontime="+84" swimtime="00:01:32.25" resultid="22953" heatid="24379" lane="2" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="328" reactiontime="+74" swimtime="00:00:42.63" resultid="22954" heatid="24457" lane="3" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-02-09" firstname="Piotr" gender="M" lastname="Iłendo" nation="POL" athleteid="22972">
              <RESULTS>
                <RESULT eventid="1079" points="561" reactiontime="+72" swimtime="00:00:25.34" resultid="22973" heatid="24295" lane="2" entrytime="00:00:26.00" />
                <RESULT eventid="1205" points="530" swimtime="00:00:29.64" resultid="22974" heatid="24335" lane="3" entrytime="00:00:29.90" />
                <RESULT eventid="1273" points="572" swimtime="00:00:56.50" resultid="22975" heatid="24364" lane="4" entrytime="00:00:57.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="512" reactiontime="+53" swimtime="00:02:07.42" resultid="22976" heatid="24424" lane="7" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                    <SPLIT distance="100" swimtime="00:01:01.79" />
                    <SPLIT distance="150" swimtime="00:01:35.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="439" reactiontime="+66" swimtime="00:02:27.17" resultid="22977" heatid="24452" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                    <SPLIT distance="100" swimtime="00:01:10.85" />
                    <SPLIT distance="150" swimtime="00:01:49.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-03-03" firstname="Mateusz" gender="M" lastname="Kliza" nation="POL" athleteid="22966">
              <RESULTS>
                <RESULT eventid="1113" points="501" reactiontime="+76" swimtime="00:02:23.46" resultid="22967" heatid="24307" lane="3" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.95" />
                    <SPLIT distance="100" swimtime="00:01:06.37" />
                    <SPLIT distance="150" swimtime="00:01:48.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="575" swimtime="00:00:56.41" resultid="22968" heatid="24364" lane="3" entrytime="00:00:57.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="510" swimtime="00:02:07.66" resultid="22969" heatid="24424" lane="2" entrytime="00:02:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.09" />
                    <SPLIT distance="100" swimtime="00:01:02.03" />
                    <SPLIT distance="150" swimtime="00:01:35.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="482" swimtime="00:05:10.86" resultid="22970" heatid="24433" lane="5" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                    <SPLIT distance="100" swimtime="00:01:06.63" />
                    <SPLIT distance="150" swimtime="00:01:48.98" />
                    <SPLIT distance="200" swimtime="00:02:32.29" />
                    <SPLIT distance="300" swimtime="00:03:57.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="500" swimtime="00:04:37.16" resultid="22971" heatid="24482" lane="3" entrytime="00:04:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:40.78" />
                    <SPLIT distance="100" swimtime="00:01:05.18" />
                    <SPLIT distance="150" swimtime="00:02:52.31" />
                    <SPLIT distance="200" swimtime="00:02:16.32" />
                    <SPLIT distance="250" swimtime="00:04:03.70" />
                    <SPLIT distance="300" swimtime="00:03:27.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-03-21" firstname="Ewa" gender="F" lastname="Markowska" nation="POL" athleteid="22947">
              <RESULTS>
                <RESULT comment="Przekroczenie limitu czasu" eventid="1165" reactiontime="+109" status="OTL" swimtime="00:00:00.00" resultid="22948" heatid="24319" lane="1" entrytime="00:25:50.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.98" />
                    <SPLIT distance="100" swimtime="00:01:38.35" />
                    <SPLIT distance="150" swimtime="00:02:33.89" />
                    <SPLIT distance="200" swimtime="00:03:30.52" />
                    <SPLIT distance="250" swimtime="00:04:28.72" />
                    <SPLIT distance="300" swimtime="00:05:26.32" />
                    <SPLIT distance="350" swimtime="00:06:24.18" />
                    <SPLIT distance="400" swimtime="00:07:22.21" />
                    <SPLIT distance="450" swimtime="00:08:20.77" />
                    <SPLIT distance="500" swimtime="00:09:19.16" />
                    <SPLIT distance="550" swimtime="00:10:17.14" />
                    <SPLIT distance="600" swimtime="00:11:16.59" />
                    <SPLIT distance="650" swimtime="00:12:15.53" />
                    <SPLIT distance="700" swimtime="00:13:14.55" />
                    <SPLIT distance="750" swimtime="00:14:14.22" />
                    <SPLIT distance="800" swimtime="00:15:13.76" />
                    <SPLIT distance="850" swimtime="00:16:14.15" />
                    <SPLIT distance="900" swimtime="00:17:13.56" />
                    <SPLIT distance="950" swimtime="00:18:13.45" />
                    <SPLIT distance="1000" swimtime="00:19:12.87" />
                    <SPLIT distance="1050" swimtime="00:20:12.09" />
                    <SPLIT distance="1100" swimtime="00:21:13.93" />
                    <SPLIT distance="1150" swimtime="00:22:12.97" />
                    <SPLIT distance="1200" swimtime="00:23:13.85" />
                    <SPLIT distance="1250" swimtime="00:24:14.36" />
                    <SPLIT distance="1300" swimtime="00:25:13.38" />
                    <SPLIT distance="1350" swimtime="00:26:00.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="150" reactiontime="+106" swimtime="00:08:20.74" resultid="22949" heatid="24429" lane="9" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.63" />
                    <SPLIT distance="100" swimtime="00:02:14.98" />
                    <SPLIT distance="150" swimtime="00:03:23.25" />
                    <SPLIT distance="200" swimtime="00:04:29.21" />
                    <SPLIT distance="250" swimtime="00:05:28.28" />
                    <SPLIT distance="300" swimtime="00:06:29.08" />
                    <SPLIT distance="350" swimtime="00:07:26.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-06-10" firstname="Dawid" gender="M" lastname="Perkowski" nation="POL" athleteid="22961">
              <RESULTS>
                <RESULT eventid="1079" points="524" reactiontime="+64" swimtime="00:00:25.93" resultid="22962" heatid="24295" lane="8" entrytime="00:00:26.10" />
                <RESULT eventid="1341" points="402" swimtime="00:02:30.99" resultid="22963" heatid="24371" lane="6" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                    <SPLIT distance="100" swimtime="00:01:08.69" />
                    <SPLIT distance="150" swimtime="00:01:47.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="528" swimtime="00:00:27.54" resultid="22964" heatid="24397" lane="5" entrytime="00:00:27.30" />
                <RESULT eventid="1613" points="514" swimtime="00:01:02.18" resultid="22965" heatid="24442" lane="9" entrytime="00:01:02.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-09-27" firstname="Józef" gender="M" lastname="Sawicki" nation="POL" athleteid="22960" />
            <ATHLETE birthdate="1979-01-24" firstname="Humbla" gender="M" lastname="Sebastian" nation="POL" athleteid="22930">
              <RESULTS>
                <RESULT eventid="1079" points="489" reactiontime="+79" swimtime="00:00:26.54" resultid="22931" heatid="24294" lane="1" entrytime="00:00:26.79" />
                <RESULT eventid="1113" points="419" reactiontime="+84" swimtime="00:02:32.25" resultid="22932" heatid="24306" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.46" />
                    <SPLIT distance="100" swimtime="00:01:09.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="435" reactiontime="+65" swimtime="00:00:31.67" resultid="22933" heatid="24335" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="1440" points="473" swimtime="00:00:28.58" resultid="22934" heatid="24396" lane="5" entrytime="00:00:28.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-08-16" firstname="Karol" gender="M" lastname="Traciecki" nation="POL" athleteid="23414">
              <RESULTS>
                <RESULT eventid="1239" points="287" reactiontime="+85" swimtime="00:03:11.87" resultid="23415" heatid="24341" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                    <SPLIT distance="100" swimtime="00:01:27.68" />
                    <SPLIT distance="150" swimtime="00:02:19.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="263" reactiontime="+73" swimtime="00:01:29.07" resultid="23416" heatid="24380" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="23417" heatid="24300" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-17" firstname="Filip" gender="M" lastname="Walczuk" nation="POL" athleteid="22940">
              <RESULTS>
                <RESULT eventid="1079" points="399" reactiontime="+103" swimtime="00:00:28.38" resultid="22941" heatid="24293" lane="0" entrytime="00:00:27.80" />
                <RESULT eventid="1205" points="302" swimtime="00:00:35.75" resultid="22942" heatid="24334" lane="9" entrytime="00:00:33.90" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="22943" heatid="24361" lane="8" entrytime="00:01:04.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-13" firstname="Dawid" gender="M" lastname="Świderski" nation="POL" athleteid="22935">
              <RESULTS>
                <RESULT eventid="1079" points="471" reactiontime="+85" swimtime="00:00:26.86" resultid="22936" heatid="24294" lane="7" entrytime="00:00:26.78" />
                <RESULT eventid="1341" status="DNS" swimtime="00:00:00.00" resultid="22937" heatid="24371" lane="8" entrytime="00:02:30.00" />
                <RESULT eventid="1440" points="465" reactiontime="+77" swimtime="00:00:28.74" resultid="22938" heatid="24397" lane="7" entrytime="00:00:28.39" />
                <RESULT eventid="1613" points="393" swimtime="00:01:07.96" resultid="22939" heatid="24441" lane="6" entrytime="00:01:04.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" points="515" swimtime="00:01:45.81" resultid="22980" heatid="24427" lane="6" entrytime="00:01:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.62" />
                    <SPLIT distance="100" swimtime="00:00:53.72" />
                    <SPLIT distance="150" swimtime="00:01:19.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22935" number="1" />
                    <RELAYPOSITION athleteid="22940" number="2" />
                    <RELAYPOSITION athleteid="22930" number="3" reactiontime="+7" />
                    <RELAYPOSITION athleteid="22944" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" points="429" reactiontime="+60" swimtime="00:02:03.80" resultid="22981" heatid="24374" lane="6" entrytime="00:01:57.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                    <SPLIT distance="100" swimtime="00:01:08.18" />
                    <SPLIT distance="150" swimtime="00:01:36.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22940" number="1" reactiontime="+60" />
                    <RELAYPOSITION athleteid="22935" number="2" />
                    <RELAYPOSITION athleteid="22930" number="3" reactiontime="+14" />
                    <RELAYPOSITION athleteid="22944" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1548" points="444" reactiontime="+76" swimtime="00:01:51.20" resultid="22979" heatid="24427" lane="3" entrytime="00:01:46.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.83" />
                    <SPLIT distance="100" swimtime="00:00:59.13" />
                    <SPLIT distance="150" swimtime="00:01:25.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22966" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="23414" number="2" />
                    <RELAYPOSITION athleteid="22955" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="22972" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" points="432" reactiontime="+68" swimtime="00:02:03.59" resultid="22982" heatid="24374" lane="5" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22972" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="22966" number="2" />
                    <RELAYPOSITION athleteid="22955" number="3" reactiontime="+12" />
                    <RELAYPOSITION athleteid="23414" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1698" reactiontime="+75" swimtime="00:02:48.70" resultid="22978" heatid="24468" lane="5" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.64" />
                    <SPLIT distance="100" swimtime="00:01:27.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22940" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="22947" number="2" />
                    <RELAYPOSITION athleteid="22955" number="3" reactiontime="+67" />
                    <RELAYPOSITION athleteid="22950" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1130" reactiontime="+71" swimtime="00:02:04.14" resultid="22983" heatid="24309" lane="7" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.89" />
                    <SPLIT distance="100" swimtime="00:00:59.06" />
                    <SPLIT distance="150" swimtime="00:01:37.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22955" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="22950" number="2" />
                    <RELAYPOSITION athleteid="22947" number="3" />
                    <RELAYPOSITION athleteid="22944" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="KORONA KRA" nation="POL" region="KR" clubid="20781" name="Korona Kraków Masters">
          <CONTACT city="Kraków" name="Mariola Kuliś" phone="500677133" state="MAŁ" />
          <ATHLETES>
            <ATHLETE birthdate="1988-10-27" firstname="Karolina" gender="F" lastname="Caba" nation="POL" athleteid="21387">
              <RESULTS>
                <RESULT eventid="1062" points="359" reactiontime="+100" swimtime="00:00:33.30" resultid="21388" heatid="24278" lane="3" entrytime="00:00:34.00" />
                <RESULT eventid="1147" points="336" reactiontime="+105" swimtime="00:11:37.16" resultid="21389" heatid="24312" lane="1" entrytime="00:11:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                    <SPLIT distance="100" swimtime="00:01:17.49" />
                    <SPLIT distance="150" swimtime="00:02:00.05" />
                    <SPLIT distance="200" swimtime="00:02:43.30" />
                    <SPLIT distance="250" swimtime="00:03:27.09" />
                    <SPLIT distance="300" swimtime="00:04:11.51" />
                    <SPLIT distance="350" swimtime="00:04:56.25" />
                    <SPLIT distance="400" swimtime="00:05:40.95" />
                    <SPLIT distance="450" swimtime="00:06:26.79" />
                    <SPLIT distance="500" swimtime="00:07:11.94" />
                    <SPLIT distance="550" swimtime="00:07:56.77" />
                    <SPLIT distance="600" swimtime="00:08:41.71" />
                    <SPLIT distance="650" swimtime="00:09:26.39" />
                    <SPLIT distance="700" swimtime="00:10:11.32" />
                    <SPLIT distance="750" swimtime="00:10:54.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-07-18" firstname="Kamil" gender="M" lastname="Dubicki" nation="POL" athleteid="21384">
              <RESULTS>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="21385" heatid="24395" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1474" points="276" reactiontime="+63" swimtime="00:01:19.58" resultid="21386" heatid="24406" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-12-23" firstname="Anna" gender="F" lastname="Janeczko" nation="POL" athleteid="21310">
              <RESULTS>
                <RESULT eventid="1423" points="299" reactiontime="+81" swimtime="00:00:36.52" resultid="21311" heatid="24387" lane="3" entrytime="00:00:39.90" />
                <RESULT eventid="1555" points="224" reactiontime="+59" swimtime="00:07:18.03" resultid="21312" heatid="24429" lane="0" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.20" />
                    <SPLIT distance="100" swimtime="00:01:44.77" />
                    <SPLIT distance="150" swimtime="00:02:41.99" />
                    <SPLIT distance="200" swimtime="00:03:40.26" />
                    <SPLIT distance="250" swimtime="00:04:41.10" />
                    <SPLIT distance="300" swimtime="00:05:41.56" />
                    <SPLIT distance="350" swimtime="00:06:31.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="176" reactiontime="+62" swimtime="00:01:38.97" resultid="21313" heatid="24435" lane="6" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-07-27" firstname="Mariola" gender="F" lastname="Kuliś" nation="POL" athleteid="21296">
              <RESULTS>
                <RESULT eventid="1062" points="450" reactiontime="+76" swimtime="00:00:30.87" resultid="21297" heatid="24280" lane="6" entrytime="00:00:30.50" />
                <RESULT eventid="1187" points="390" swimtime="00:00:37.03" resultid="21298" heatid="24326" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="1256" points="369" reactiontime="+68" swimtime="00:01:12.08" resultid="21299" heatid="24352" lane="7" entrytime="00:01:10.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="373" swimtime="00:00:33.91" resultid="21300" heatid="24389" lane="1" entrytime="00:00:33.70" />
                <RESULT eventid="1457" points="330" swimtime="00:01:23.93" resultid="21301" heatid="24401" lane="3" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="429" reactiontime="+67" swimtime="00:00:38.98" resultid="21302" heatid="24458" lane="7" entrytime="00:00:37.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-09-15" firstname="Mirosława" gender="F" lastname="Legutko" nation="POL" athleteid="21375">
              <RESULTS>
                <RESULT eventid="1062" points="296" reactiontime="+111" swimtime="00:00:35.48" resultid="21376" heatid="24278" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="1096" points="179" reactiontime="+107" swimtime="00:03:43.40" resultid="21377" heatid="24297" lane="5" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.41" />
                    <SPLIT distance="100" swimtime="00:01:49.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="218" reactiontime="+83" swimtime="00:01:25.85" resultid="21378" heatid="24347" lane="5" />
                <RESULT eventid="1324" points="124" reactiontime="+111" swimtime="00:04:03.75" resultid="21379" heatid="24367" lane="8" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.52" />
                    <SPLIT distance="100" swimtime="00:01:54.71" />
                    <SPLIT distance="150" swimtime="00:02:59.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="183" reactiontime="+87" swimtime="00:00:42.98" resultid="21380" heatid="24387" lane="1" entrytime="00:00:45.00" />
                <RESULT eventid="1555" points="169" reactiontime="+101" swimtime="00:08:00.94" resultid="21381" heatid="24428" lane="4" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.68" />
                    <SPLIT distance="100" swimtime="00:01:56.56" />
                    <SPLIT distance="150" swimtime="00:02:58.75" />
                    <SPLIT distance="200" swimtime="00:04:02.68" />
                    <SPLIT distance="250" swimtime="00:05:09.39" />
                    <SPLIT distance="300" swimtime="00:06:17.01" />
                    <SPLIT distance="350" swimtime="00:07:09.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="125" reactiontime="+102" swimtime="00:01:50.69" resultid="21382" heatid="24434" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="188" reactiontime="+78" swimtime="00:00:51.26" resultid="21383" heatid="24454" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-04-20" firstname="Agnieszka" gender="F" lastname="Macierzewska" nation="POL" athleteid="21314">
              <RESULTS>
                <RESULT eventid="1062" points="323" reactiontime="+100" swimtime="00:00:34.48" resultid="21315" heatid="24278" lane="4" entrytime="00:00:33.50" />
                <RESULT eventid="1147" points="268" reactiontime="+104" swimtime="00:12:31.18" resultid="21316" heatid="24311" lane="3" entrytime="00:12:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.82" />
                    <SPLIT distance="100" swimtime="00:01:24.47" />
                    <SPLIT distance="150" swimtime="00:02:10.94" />
                    <SPLIT distance="200" swimtime="00:02:58.26" />
                    <SPLIT distance="250" swimtime="00:03:46.16" />
                    <SPLIT distance="300" swimtime="00:04:34.28" />
                    <SPLIT distance="350" swimtime="00:05:22.83" />
                    <SPLIT distance="400" swimtime="00:06:11.87" />
                    <SPLIT distance="450" swimtime="00:07:00.03" />
                    <SPLIT distance="500" swimtime="00:07:48.22" />
                    <SPLIT distance="550" swimtime="00:08:36.35" />
                    <SPLIT distance="600" swimtime="00:09:24.90" />
                    <SPLIT distance="650" swimtime="00:10:12.82" />
                    <SPLIT distance="700" swimtime="00:11:00.91" />
                    <SPLIT distance="750" swimtime="00:11:47.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="311" reactiontime="+97" swimtime="00:01:16.32" resultid="21317" heatid="24351" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="206" reactiontime="+89" swimtime="00:03:25.92" resultid="21318" heatid="24367" lane="1" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.15" />
                    <SPLIT distance="100" swimtime="00:01:36.31" />
                    <SPLIT distance="150" swimtime="00:02:32.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="254" reactiontime="+90" swimtime="00:00:38.54" resultid="21319" heatid="24387" lane="4" entrytime="00:00:39.00" />
                <RESULT eventid="1491" points="298" reactiontime="+96" swimtime="00:02:49.07" resultid="21320" heatid="24412" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.80" />
                    <SPLIT distance="100" swimtime="00:01:22.03" />
                    <SPLIT distance="150" swimtime="00:02:06.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="220" reactiontime="+68" swimtime="00:01:31.88" resultid="21321" heatid="24436" lane="0" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="276" reactiontime="+84" swimtime="00:06:02.79" resultid="21322" heatid="24472" lane="1" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.58" />
                    <SPLIT distance="100" swimtime="00:01:24.31" />
                    <SPLIT distance="150" swimtime="00:02:10.46" />
                    <SPLIT distance="200" swimtime="00:02:57.77" />
                    <SPLIT distance="250" swimtime="00:03:45.80" />
                    <SPLIT distance="300" swimtime="00:04:33.65" />
                    <SPLIT distance="350" swimtime="00:05:20.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-08-26" firstname="Andrzej" gender="M" lastname="Mleczko" nation="POL" athleteid="21323">
              <RESULTS>
                <RESULT eventid="1113" points="120" reactiontime="+146" swimtime="00:03:51.00" resultid="21324" heatid="24302" lane="4" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.76" />
                    <SPLIT distance="100" swimtime="00:01:58.11" />
                    <SPLIT distance="150" swimtime="00:03:02.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14189" points="122" reactiontime="+137" swimtime="00:15:10.99" resultid="21325" heatid="24314" lane="5" entrytime="00:14:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.70" />
                    <SPLIT distance="100" swimtime="00:01:49.85" />
                    <SPLIT distance="150" swimtime="00:02:48.19" />
                    <SPLIT distance="200" swimtime="00:03:45.97" />
                    <SPLIT distance="250" swimtime="00:04:44.66" />
                    <SPLIT distance="300" swimtime="00:05:42.55" />
                    <SPLIT distance="350" swimtime="00:06:41.64" />
                    <SPLIT distance="400" swimtime="00:07:38.64" />
                    <SPLIT distance="450" swimtime="00:08:36.47" />
                    <SPLIT distance="500" swimtime="00:09:33.53" />
                    <SPLIT distance="550" swimtime="00:10:30.74" />
                    <SPLIT distance="600" swimtime="00:11:27.82" />
                    <SPLIT distance="650" swimtime="00:12:23.85" />
                    <SPLIT distance="700" swimtime="00:13:22.06" />
                    <SPLIT distance="750" swimtime="00:14:20.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="221" reactiontime="+98" swimtime="00:01:17.52" resultid="21326" heatid="24357" lane="2" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="52" reactiontime="+116" swimtime="00:04:57.26" resultid="21327" heatid="24369" lane="0" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.52" />
                    <SPLIT distance="100" swimtime="00:00:33.90" />
                    <SPLIT distance="150" swimtime="00:03:34.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="138" reactiontime="+111" swimtime="00:03:17.16" resultid="21328" heatid="24418" lane="6" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.19" />
                    <SPLIT distance="100" swimtime="00:01:37.20" />
                    <SPLIT distance="150" swimtime="00:02:27.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="97" reactiontime="+107" swimtime="00:08:50.56" resultid="21329" heatid="24431" lane="9" entrytime="00:08:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.44" />
                    <SPLIT distance="100" swimtime="00:02:09.97" />
                    <SPLIT distance="150" swimtime="00:03:23.88" />
                    <SPLIT distance="200" swimtime="00:04:31.97" />
                    <SPLIT distance="250" swimtime="00:05:42.75" />
                    <SPLIT distance="300" swimtime="00:06:57.56" />
                    <SPLIT distance="350" swimtime="00:07:55.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="75" reactiontime="+96" swimtime="00:01:57.95" resultid="21330" heatid="24438" lane="8" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="132" reactiontime="+102" swimtime="00:07:11.41" resultid="21331" heatid="24476" lane="5" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.43" />
                    <SPLIT distance="200" swimtime="00:03:34.04" />
                    <SPLIT distance="300" swimtime="00:05:27.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-05-06" firstname="Matteo" gender="M" lastname="Morlupi" nation="POL" athleteid="21390">
              <RESULTS>
                <RESULT eventid="1681" points="247" reactiontime="+82" swimtime="00:00:41.31" resultid="21391" heatid="24462" lane="7" entrytime="00:00:41.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-05-29" firstname="Małgorzata" gender="F" lastname="Orlewicz-Musiał" nation="POL" athleteid="21332">
              <RESULTS>
                <RESULT eventid="1096" points="85" reactiontime="+99" swimtime="00:04:46.14" resultid="21333" heatid="24297" lane="7" entrytime="00:04:34.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.50" />
                    <SPLIT distance="100" swimtime="00:02:15.18" />
                    <SPLIT distance="150" swimtime="00:03:43.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" reactiontime="+107" status="OTL" swimtime="00:33:16.55" resultid="21334" heatid="24318" lane="4" entrytime="00:31:33.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.91" />
                    <SPLIT distance="100" swimtime="00:01:55.16" />
                    <SPLIT distance="150" swimtime="00:02:59.75" />
                    <SPLIT distance="200" swimtime="00:04:04.29" />
                    <SPLIT distance="250" swimtime="00:05:10.18" />
                    <SPLIT distance="300" swimtime="00:06:15.24" />
                    <SPLIT distance="350" swimtime="00:07:20.47" />
                    <SPLIT distance="400" swimtime="00:08:27.01" />
                    <SPLIT distance="450" swimtime="00:09:33.85" />
                    <SPLIT distance="500" swimtime="00:10:41.65" />
                    <SPLIT distance="550" swimtime="00:11:48.74" />
                    <SPLIT distance="600" swimtime="00:12:54.74" />
                    <SPLIT distance="650" swimtime="00:14:01.61" />
                    <SPLIT distance="700" swimtime="00:15:09.10" />
                    <SPLIT distance="750" swimtime="00:16:18.16" />
                    <SPLIT distance="800" swimtime="00:17:25.44" />
                    <SPLIT distance="850" swimtime="00:18:32.58" />
                    <SPLIT distance="900" swimtime="00:19:39.16" />
                    <SPLIT distance="950" swimtime="00:20:47.03" />
                    <SPLIT distance="1000" swimtime="00:21:54.74" />
                    <SPLIT distance="1050" swimtime="00:23:02.78" />
                    <SPLIT distance="1100" swimtime="00:24:09.59" />
                    <SPLIT distance="1150" swimtime="00:25:18.00" />
                    <SPLIT distance="1200" swimtime="00:26:26.10" />
                    <SPLIT distance="1250" swimtime="00:27:35.29" />
                    <SPLIT distance="1300" swimtime="00:28:43.69" />
                    <SPLIT distance="1350" swimtime="00:29:52.12" />
                    <SPLIT distance="1400" swimtime="00:31:02.26" />
                    <SPLIT distance="1450" swimtime="00:32:10.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="87" swimtime="00:01:01.04" resultid="21335" heatid="24324" lane="1" entrytime="00:01:01.52" />
                <RESULT eventid="1324" points="52" reactiontime="+90" swimtime="00:05:25.60" resultid="21336" heatid="24366" lane="3" entrytime="00:04:48.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.00" />
                    <SPLIT distance="100" swimtime="00:02:28.15" />
                    <SPLIT distance="150" swimtime="00:03:59.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="65" reactiontime="+73" swimtime="00:01:00.63" resultid="21337" heatid="24386" lane="1" />
                <RESULT eventid="1555" points="80" reactiontime="+89" swimtime="00:10:17.06" resultid="21338" heatid="24428" lane="3" entrytime="00:09:55.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.76" />
                    <SPLIT distance="100" swimtime="00:02:24.76" />
                    <SPLIT distance="150" swimtime="00:03:45.20" />
                    <SPLIT distance="200" swimtime="00:05:03.70" />
                    <SPLIT distance="250" swimtime="00:06:34.12" />
                    <SPLIT distance="300" swimtime="00:08:03.75" />
                    <SPLIT distance="350" swimtime="00:09:11.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="59" reactiontime="+76" swimtime="00:02:21.81" resultid="21339" heatid="24435" lane="8" entrytime="00:02:10.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="91" reactiontime="+106" swimtime="00:08:43.86" resultid="21340" heatid="24470" lane="2" entrytime="00:08:39.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.00" />
                    <SPLIT distance="100" swimtime="00:01:58.12" />
                    <SPLIT distance="150" swimtime="00:03:04.95" />
                    <SPLIT distance="200" swimtime="00:04:12.60" />
                    <SPLIT distance="250" swimtime="00:05:19.85" />
                    <SPLIT distance="300" swimtime="00:06:28.11" />
                    <SPLIT distance="350" swimtime="00:07:36.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-11-10" firstname="Waldemar" gender="M" lastname="Piszczek" nation="POL" athleteid="21341">
              <RESULTS>
                <RESULT eventid="1079" points="325" reactiontime="+86" swimtime="00:00:30.41" resultid="21342" heatid="24289" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="21343" heatid="24304" lane="7" entrytime="00:03:00.00" />
                <RESULT eventid="1205" points="311" swimtime="00:00:35.40" resultid="21344" heatid="24333" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="1239" points="251" reactiontime="+43" swimtime="00:03:20.61" resultid="21345" heatid="24344" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.14" />
                    <SPLIT distance="100" swimtime="00:01:37.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="372" reactiontime="+63" swimtime="00:00:30.95" resultid="21346" heatid="24394" lane="4" entrytime="00:00:31.50" />
                <RESULT eventid="1474" points="293" swimtime="00:01:18.00" resultid="21347" heatid="24406" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="21348" heatid="24440" lane="1" entrytime="00:01:16.00" />
                <RESULT eventid="1681" points="328" reactiontime="+50" swimtime="00:00:37.59" resultid="21349" heatid="24463" lane="5" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-02-18" firstname="Bartosz" gender="M" lastname="Próchniewicz" nation="POL" athleteid="21392">
              <RESULTS>
                <RESULT eventid="1079" points="171" reactiontime="+88" swimtime="00:00:37.61" resultid="21393" heatid="24284" lane="0" entrytime="00:00:45.00" />
                <RESULT eventid="1647" points="79" reactiontime="+140" swimtime="00:04:20.17" resultid="21394" heatid="24447" lane="4" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.99" />
                    <SPLIT distance="150" swimtime="00:03:14.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-21" firstname="Adam" gender="M" lastname="Pycia" nation="POL" athleteid="21350">
              <RESULTS>
                <RESULT eventid="1079" points="287" reactiontime="+94" swimtime="00:00:31.70" resultid="21351" heatid="24287" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="14189" points="220" reactiontime="+93" swimtime="00:12:28.82" resultid="21352" heatid="24316" lane="7" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.66" />
                    <SPLIT distance="100" swimtime="00:01:19.39" />
                    <SPLIT distance="150" swimtime="00:02:04.79" />
                    <SPLIT distance="200" swimtime="00:02:51.42" />
                    <SPLIT distance="250" swimtime="00:03:40.38" />
                    <SPLIT distance="300" swimtime="00:04:28.19" />
                    <SPLIT distance="350" swimtime="00:05:16.24" />
                    <SPLIT distance="400" swimtime="00:06:04.20" />
                    <SPLIT distance="450" swimtime="00:06:52.27" />
                    <SPLIT distance="500" swimtime="00:07:40.19" />
                    <SPLIT distance="550" swimtime="00:08:28.22" />
                    <SPLIT distance="600" swimtime="00:09:16.91" />
                    <SPLIT distance="650" swimtime="00:10:06.00" />
                    <SPLIT distance="700" swimtime="00:10:54.47" />
                    <SPLIT distance="750" swimtime="00:11:43.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="154" swimtime="00:00:44.77" resultid="21353" heatid="24332" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1239" points="239" reactiontime="+99" swimtime="00:03:24.11" resultid="21354" heatid="24343" lane="4" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.80" />
                    <SPLIT distance="100" swimtime="00:01:38.39" />
                    <SPLIT distance="150" swimtime="00:02:33.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="256" reactiontime="+93" swimtime="00:01:29.88" resultid="21355" heatid="24383" lane="8" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="200" reactiontime="+45" swimtime="00:00:38.05" resultid="21356" heatid="24392" lane="0" entrytime="00:00:38.60" />
                <RESULT eventid="1681" points="268" swimtime="00:00:40.20" resultid="21357" heatid="24463" lane="9" entrytime="00:00:39.80" />
                <RESULT eventid="1744" points="233" reactiontime="+93" swimtime="00:05:57.47" resultid="21358" heatid="24478" lane="7" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.79" />
                    <SPLIT distance="100" swimtime="00:01:21.30" />
                    <SPLIT distance="150" swimtime="00:02:06.89" />
                    <SPLIT distance="200" swimtime="00:02:53.63" />
                    <SPLIT distance="250" swimtime="00:03:40.97" />
                    <SPLIT distance="300" swimtime="00:04:28.58" />
                    <SPLIT distance="350" swimtime="00:05:16.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-07-29" firstname="Jolanta" gender="F" lastname="Uczarczyk" nation="POL" athleteid="21359">
              <RESULTS>
                <RESULT eventid="1062" points="210" reactiontime="+106" swimtime="00:00:39.80" resultid="21360" heatid="24278" lane="0" entrytime="00:00:37.43" />
                <RESULT eventid="1096" points="149" reactiontime="+107" swimtime="00:03:57.37" resultid="21361" heatid="24297" lane="4" entrytime="00:03:39.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.45" />
                    <SPLIT distance="100" swimtime="00:01:52.25" />
                    <SPLIT distance="150" swimtime="00:03:00.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="119" swimtime="00:00:54.90" resultid="21362" heatid="24325" lane="9" entrytime="00:00:49.67" />
                <RESULT eventid="1324" points="110" reactiontime="+81" swimtime="00:04:13.99" resultid="21363" heatid="24367" lane="0" entrytime="00:03:53.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.15" />
                    <SPLIT distance="100" swimtime="00:02:00.87" />
                    <SPLIT distance="150" swimtime="00:03:07.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="136" reactiontime="+76" swimtime="00:00:47.50" resultid="21364" heatid="24387" lane="7" entrytime="00:00:43.63" />
                <RESULT eventid="1491" points="137" reactiontime="+95" swimtime="00:03:39.12" resultid="21365" heatid="24411" lane="2" entrytime="00:03:29.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.49" />
                    <SPLIT distance="100" swimtime="00:01:42.65" />
                    <SPLIT distance="150" swimtime="00:02:42.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="114" reactiontime="+88" swimtime="00:01:54.27" resultid="21366" heatid="24435" lane="2" entrytime="00:01:43.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="121" reactiontime="+70" swimtime="00:07:56.94" resultid="21367" heatid="24469" lane="5">
                  <SPLITS>
                    <SPLIT distance="300" swimtime="00:05:57.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-07-04" firstname="Stanisław" gender="M" lastname="Waga" nation="POL" athleteid="21368">
              <RESULTS>
                <RESULT eventid="1079" points="81" reactiontime="+123" swimtime="00:00:48.22" resultid="21369" heatid="24284" lane="9" entrytime="00:00:48.00" />
                <RESULT eventid="14207" reactiontime="+135" status="OTL" swimtime="00:36:19.70" resultid="21370" heatid="24320" lane="7" entrytime="00:33:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.57" />
                    <SPLIT distance="100" swimtime="00:02:10.77" />
                    <SPLIT distance="150" swimtime="00:03:22.10" />
                    <SPLIT distance="200" swimtime="00:04:33.66" />
                    <SPLIT distance="250" swimtime="00:05:44.67" />
                    <SPLIT distance="300" swimtime="00:06:54.65" />
                    <SPLIT distance="350" swimtime="00:08:06.23" />
                    <SPLIT distance="400" swimtime="00:09:15.74" />
                    <SPLIT distance="450" swimtime="00:10:27.82" />
                    <SPLIT distance="500" swimtime="00:11:39.74" />
                    <SPLIT distance="550" swimtime="00:12:50.42" />
                    <SPLIT distance="600" swimtime="00:14:02.54" />
                    <SPLIT distance="650" swimtime="00:15:16.45" />
                    <SPLIT distance="700" swimtime="00:16:30.98" />
                    <SPLIT distance="750" swimtime="00:20:13.95" />
                    <SPLIT distance="800" swimtime="00:18:59.86" />
                    <SPLIT distance="850" swimtime="00:22:40.62" />
                    <SPLIT distance="900" swimtime="00:21:27.14" />
                    <SPLIT distance="950" swimtime="00:25:10.29" />
                    <SPLIT distance="1000" swimtime="00:23:56.61" />
                    <SPLIT distance="1050" swimtime="00:27:39.80" />
                    <SPLIT distance="1100" swimtime="00:26:26.81" />
                    <SPLIT distance="1150" swimtime="00:30:08.98" />
                    <SPLIT distance="1200" swimtime="00:28:56.96" />
                    <SPLIT distance="1250" swimtime="00:32:41.58" />
                    <SPLIT distance="1300" swimtime="00:31:24.99" />
                    <SPLIT distance="1350" swimtime="00:35:08.87" />
                    <SPLIT distance="1400" swimtime="00:33:56.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="70" reactiontime="+98" swimtime="00:01:53.46" resultid="21371" heatid="24355" lane="2" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="61" reactiontime="+89" swimtime="00:04:18.99" resultid="21372" heatid="24416" lane="2" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.78" />
                    <SPLIT distance="100" swimtime="00:01:59.53" />
                    <SPLIT distance="150" swimtime="00:03:10.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="53" reactiontime="+77" swimtime="00:01:09.08" resultid="21373" heatid="24460" lane="9" entrytime="00:01:10.00" />
                <RESULT eventid="1744" points="60" reactiontime="+108" swimtime="00:09:20.16" resultid="21374" heatid="24475" lane="1" entrytime="00:08:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.79" />
                    <SPLIT distance="100" swimtime="00:02:14.08" />
                    <SPLIT distance="150" swimtime="00:03:28.34" />
                    <SPLIT distance="200" swimtime="00:04:41.80" />
                    <SPLIT distance="250" swimtime="00:05:54.12" />
                    <SPLIT distance="300" swimtime="00:07:07.60" />
                    <SPLIT distance="350" swimtime="00:08:16.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-30" firstname="Piotr" gender="M" lastname="Łysiak" nation="POL" athleteid="21303">
              <RESULTS>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="21304" heatid="24333" lane="7" entrytime="00:00:36.00" />
                <RESULT eventid="1239" points="303" reactiontime="+52" swimtime="00:03:08.57" resultid="21305" heatid="24345" lane="6" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.87" />
                    <SPLIT distance="100" swimtime="00:01:30.42" />
                    <SPLIT distance="150" swimtime="00:02:18.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="272" swimtime="00:01:28.05" resultid="21306" heatid="24384" lane="9" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="215" reactiontime="+72" swimtime="00:01:26.44" resultid="21307" heatid="24406" lane="2" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="210" reactiontime="+63" swimtime="00:03:08.17" resultid="21308" heatid="24450" lane="9" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.09" />
                    <SPLIT distance="100" swimtime="00:01:31.92" />
                    <SPLIT distance="150" swimtime="00:02:21.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="21309" heatid="24462" lane="4" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" name="Korona Kraków Masters E" number="1">
              <RESULTS>
                <RESULT eventid="1130" reactiontime="+79" swimtime="00:02:09.66" resultid="21395" heatid="24308" lane="5" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                    <SPLIT distance="100" swimtime="00:01:05.15" />
                    <SPLIT distance="150" swimtime="00:01:40.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21296" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="21314" number="2" />
                    <RELAYPOSITION athleteid="21323" number="3" reactiontime="+67" />
                    <RELAYPOSITION athleteid="21341" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" reactiontime="+86" swimtime="00:02:27.70" resultid="21396" heatid="24468" lane="0" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.93" />
                    <SPLIT distance="100" swimtime="00:01:21.40" />
                    <SPLIT distance="150" swimtime="00:01:52.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21314" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="21296" number="2" />
                    <RELAYPOSITION athleteid="21341" number="3" />
                    <RELAYPOSITION athleteid="21323" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00816" nation="POL" region="ZAC" clubid="20723" name="KP Neptun Stargard">
          <CONTACT city="Stargard" email="prezes@mksneptun.pl" internet="www.mksneptun.pl" name="Klub Pływacki &quot;Neptun&quot;" phone="602731410" state="ZACHO" street="Os. Zachód B 15" zip="73-110" />
          <ATHLETES>
            <ATHLETE birthdate="1973-02-20" firstname="Mariusz" gender="M" lastname="Chrzan" nation="POL" athleteid="20724">
              <RESULTS>
                <RESULT eventid="1079" points="458" reactiontime="+71" swimtime="00:00:27.11" resultid="20725" heatid="24295" lane="9" entrytime="00:00:26.20" />
                <RESULT eventid="1113" points="427" reactiontime="+78" swimtime="00:02:31.34" resultid="20726" heatid="24306" lane="5" entrytime="00:02:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                    <SPLIT distance="100" swimtime="00:01:10.72" />
                    <SPLIT distance="150" swimtime="00:01:56.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="454" reactiontime="+76" swimtime="00:00:31.21" resultid="20727" heatid="24335" lane="7" entrytime="00:00:30.60" />
                <RESULT eventid="1273" points="472" swimtime="00:01:00.21" resultid="20728" heatid="24363" lane="0" entrytime="00:00:59.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="451" swimtime="00:00:29.02" resultid="20729" heatid="24397" lane="9" entrytime="00:00:28.50" />
                <RESULT eventid="1474" points="453" reactiontime="+69" swimtime="00:01:07.50" resultid="20730" heatid="24408" lane="8" entrytime="00:01:06.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="432" reactiontime="+96" swimtime="00:02:28.00" resultid="20731" heatid="24451" lane="4" entrytime="00:02:29.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                    <SPLIT distance="100" swimtime="00:01:11.63" />
                    <SPLIT distance="150" swimtime="00:01:50.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02203" nation="POL" region="LU" clubid="21660" name="KS AZS AWF Biała Podlaska">
          <CONTACT city="Biała Podlaska" email="mielnik_pawel@wp.pl" name="Mielnik" phone="697552772" state="LUB" street="Akademicka" zip="21-500" />
          <ATHLETES>
            <ATHLETE birthdate="1992-08-30" firstname="Wojciech" gender="M" lastname="Suszek" nation="POL" license="102203700023" athleteid="21661">
              <RESULTS>
                <RESULT eventid="1079" points="562" reactiontime="+62" swimtime="00:00:25.33" resultid="21662" heatid="24296" lane="8" entrytime="00:00:25.00" entrycourse="LCM" />
                <RESULT eventid="1205" points="505" reactiontime="+63" swimtime="00:00:30.13" resultid="21663" heatid="24335" lane="2" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT eventid="1273" points="613" reactiontime="+62" swimtime="00:00:55.21" resultid="21664" heatid="24365" lane="3" entrytime="00:00:54.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="582" swimtime="00:00:26.66" resultid="21665" heatid="24398" lane="8" entrytime="00:00:26.50" entrycourse="LCM" />
                <RESULT eventid="1508" points="498" swimtime="00:02:08.65" resultid="21666" heatid="24423" lane="5" entrytime="00:02:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.64" />
                    <SPLIT distance="100" swimtime="00:01:02.63" />
                    <SPLIT distance="150" swimtime="00:01:36.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="339" reactiontime="+75" swimtime="00:02:40.46" resultid="21667" heatid="24451" lane="2" entrytime="00:02:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.13" />
                    <SPLIT distance="100" swimtime="00:01:18.09" />
                    <SPLIT distance="150" swimtime="00:01:59.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="459" reactiontime="+61" swimtime="00:04:45.27" resultid="21668" heatid="24481" lane="3" entrytime="00:04:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.79" />
                    <SPLIT distance="100" swimtime="00:01:06.41" />
                    <SPLIT distance="150" swimtime="00:01:42.52" />
                    <SPLIT distance="200" swimtime="00:02:19.35" />
                    <SPLIT distance="250" swimtime="00:02:55.93" />
                    <SPLIT distance="300" swimtime="00:03:33.10" />
                    <SPLIT distance="350" swimtime="00:04:10.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="EXOBO" nation="POL" region="WIE" clubid="20156" name="KS Extreme Team Oborniki">
          <CONTACT city="OBORNIKI" email="JANWOL@POCZTA.ONET.PL" name="WOLNIEWICZ" state="WIE" street="CZARNKOWSKA 84" zip="64-600" />
          <ATHLETES>
            <ATHLETE birthdate="1948-12-22" firstname="Janusz" gender="M" lastname="Wolniewicz" nation="POL" athleteid="20157">
              <RESULTS>
                <RESULT eventid="1079" points="160" reactiontime="+99" swimtime="00:00:38.49" resultid="20158" heatid="24285" lane="4" entrytime="00:00:36.00" entrycourse="SCM" />
                <RESULT eventid="14207" reactiontime="+115" status="OTL" swimtime="00:32:23.12" resultid="20159" heatid="24320" lane="6" entrytime="00:29:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.89" />
                    <SPLIT distance="100" swimtime="00:01:51.77" />
                    <SPLIT distance="150" swimtime="00:02:56.91" />
                    <SPLIT distance="200" swimtime="00:04:02.85" />
                    <SPLIT distance="250" swimtime="00:05:08.21" />
                    <SPLIT distance="300" swimtime="00:06:14.05" />
                    <SPLIT distance="350" swimtime="00:07:18.66" />
                    <SPLIT distance="400" swimtime="00:08:24.96" />
                    <SPLIT distance="450" swimtime="00:09:28.86" />
                    <SPLIT distance="500" swimtime="00:10:33.79" />
                    <SPLIT distance="550" swimtime="00:11:38.08" />
                    <SPLIT distance="600" swimtime="00:12:42.92" />
                    <SPLIT distance="650" swimtime="00:13:48.08" />
                    <SPLIT distance="700" swimtime="00:14:53.18" />
                    <SPLIT distance="750" swimtime="00:15:58.90" />
                    <SPLIT distance="800" swimtime="00:17:03.50" />
                    <SPLIT distance="850" swimtime="00:18:09.48" />
                    <SPLIT distance="900" swimtime="00:19:14.97" />
                    <SPLIT distance="950" swimtime="00:20:21.51" />
                    <SPLIT distance="1000" swimtime="00:21:28.96" />
                    <SPLIT distance="1050" swimtime="00:22:33.22" />
                    <SPLIT distance="1100" swimtime="00:23:39.56" />
                    <SPLIT distance="1150" swimtime="00:24:45.50" />
                    <SPLIT distance="1200" swimtime="00:25:53.45" />
                    <SPLIT distance="1250" swimtime="00:26:57.44" />
                    <SPLIT distance="1300" swimtime="00:28:04.29" />
                    <SPLIT distance="1350" swimtime="00:29:09.46" />
                    <SPLIT distance="1400" swimtime="00:30:15.56" />
                    <SPLIT distance="1450" swimtime="00:31:20.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="20160" heatid="24356" lane="2" entrytime="00:01:26.00" entrycourse="SCM" />
                <RESULT eventid="1508" points="101" reactiontime="+80" swimtime="00:03:38.45" resultid="20161" heatid="24417" lane="6" entrytime="00:03:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.81" />
                    <SPLIT distance="150" swimtime="00:02:43.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="92" reactiontime="+67" swimtime="00:08:06.01" resultid="20162" heatid="24476" lane="9" entrytime="00:07:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.87" />
                    <SPLIT distance="100" swimtime="00:01:50.37" />
                    <SPLIT distance="150" swimtime="00:02:51.42" />
                    <SPLIT distance="200" swimtime="00:03:55.48" />
                    <SPLIT distance="250" swimtime="00:04:59.42" />
                    <SPLIT distance="300" swimtime="00:06:03.06" />
                    <SPLIT distance="350" swimtime="00:07:06.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00211" nation="POL" region="SLA" clubid="20732" name="KS Górnik Radlin">
          <ATHLETES>
            <ATHLETE birthdate="1985-11-07" firstname="Iwona" gender="F" lastname="Cymerman" nation="POL" athleteid="20733">
              <RESULTS>
                <RESULT eventid="1062" points="487" reactiontime="+92" swimtime="00:00:30.08" resultid="20734" heatid="24280" lane="4" entrytime="00:00:30.17" />
                <RESULT eventid="1256" points="435" reactiontime="+79" swimtime="00:01:08.20" resultid="20735" heatid="24352" lane="4" entrytime="00:01:07.20" />
                <RESULT eventid="1423" points="362" reactiontime="+87" swimtime="00:00:34.25" resultid="20736" heatid="24389" lane="8" entrytime="00:00:33.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-02-22" firstname="Ryszard" gender="M" lastname="Kubica" nation="POL" license="100211700343" athleteid="21589">
              <RESULTS>
                <RESULT eventid="1079" points="340" reactiontime="+80" swimtime="00:00:29.93" resultid="21590" heatid="24290" lane="9" entrytime="00:00:30.00" />
                <RESULT eventid="14207" points="265" reactiontime="+104" swimtime="00:22:34.72" resultid="21591" heatid="24321" lane="3" entrytime="00:23:12.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.85" />
                    <SPLIT distance="100" swimtime="00:01:23.09" />
                    <SPLIT distance="150" swimtime="00:02:07.64" />
                    <SPLIT distance="200" swimtime="00:02:53.20" />
                    <SPLIT distance="250" swimtime="00:03:38.41" />
                    <SPLIT distance="300" swimtime="00:04:24.56" />
                    <SPLIT distance="350" swimtime="00:05:10.12" />
                    <SPLIT distance="400" swimtime="00:05:56.72" />
                    <SPLIT distance="450" swimtime="00:06:41.97" />
                    <SPLIT distance="500" swimtime="00:07:28.44" />
                    <SPLIT distance="550" swimtime="00:08:13.86" />
                    <SPLIT distance="600" swimtime="00:09:00.38" />
                    <SPLIT distance="650" swimtime="00:09:45.93" />
                    <SPLIT distance="700" swimtime="00:10:32.85" />
                    <SPLIT distance="750" swimtime="00:11:18.03" />
                    <SPLIT distance="800" swimtime="00:12:04.09" />
                    <SPLIT distance="850" swimtime="00:12:48.96" />
                    <SPLIT distance="900" swimtime="00:13:35.18" />
                    <SPLIT distance="950" swimtime="00:14:20.32" />
                    <SPLIT distance="1000" swimtime="00:15:06.64" />
                    <SPLIT distance="1050" swimtime="00:15:52.51" />
                    <SPLIT distance="1100" swimtime="00:16:39.23" />
                    <SPLIT distance="1150" swimtime="00:17:25.01" />
                    <SPLIT distance="1200" swimtime="00:18:10.95" />
                    <SPLIT distance="1250" swimtime="00:18:55.81" />
                    <SPLIT distance="1300" swimtime="00:19:41.62" />
                    <SPLIT distance="1350" swimtime="00:20:26.34" />
                    <SPLIT distance="1400" swimtime="00:21:11.30" />
                    <SPLIT distance="1450" swimtime="00:21:53.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="261" swimtime="00:00:37.51" resultid="21592" heatid="24333" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="1273" points="332" reactiontime="+43" swimtime="00:01:07.74" resultid="21593" heatid="24360" lane="0" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="307" reactiontime="+95" swimtime="00:00:33.01" resultid="21594" heatid="24393" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="1508" points="286" reactiontime="+69" swimtime="00:02:34.69" resultid="21595" heatid="24420" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="100" swimtime="00:01:13.30" />
                    <SPLIT distance="150" swimtime="00:01:54.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="280" reactiontime="+72" swimtime="00:05:36.08" resultid="21596" heatid="24479" lane="2" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.70" />
                    <SPLIT distance="100" swimtime="00:01:18.25" />
                    <SPLIT distance="150" swimtime="00:02:01.23" />
                    <SPLIT distance="200" swimtime="00:02:44.87" />
                    <SPLIT distance="250" swimtime="00:03:28.77" />
                    <SPLIT distance="300" swimtime="00:04:12.24" />
                    <SPLIT distance="350" swimtime="00:04:55.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAKO" nation="POL" region="WAR" clubid="21669" name="KS MAKO">
          <CONTACT city="Warszawa" email="ania.plywanie@gmail.com" name="Anna Dąbrowska" phone="601 480 280" />
          <ATHLETES>
            <ATHLETE birthdate="1967-07-11" firstname="Paweł" gender="M" lastname="Adamowicz" nation="POL" athleteid="21670">
              <RESULTS>
                <RESULT eventid="1079" points="164" reactiontime="+94" swimtime="00:00:38.17" resultid="21671" heatid="24285" lane="0" entrytime="00:00:38.92" />
                <RESULT eventid="1273" points="126" swimtime="00:01:33.35" resultid="21672" heatid="24355" lane="5" entrytime="00:01:32.67" />
                <RESULT eventid="1406" points="176" reactiontime="+60" swimtime="00:01:41.74" resultid="21673" heatid="24381" lane="4" entrytime="00:01:42.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="111" swimtime="00:03:32.20" resultid="21674" heatid="24417" lane="8" entrytime="00:03:28.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.10" />
                    <SPLIT distance="100" swimtime="00:01:45.22" />
                    <SPLIT distance="150" swimtime="00:02:42.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="200" swimtime="00:00:44.36" resultid="21675" heatid="24461" lane="2" entrytime="00:00:44.02" />
                <RESULT eventid="1744" points="108" reactiontime="+79" swimtime="00:07:41.28" resultid="21676" heatid="24475" lane="3" entrytime="00:08:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.11" />
                    <SPLIT distance="100" swimtime="00:01:53.64" />
                    <SPLIT distance="150" swimtime="00:02:54.91" />
                    <SPLIT distance="200" swimtime="00:03:53.90" />
                    <SPLIT distance="250" swimtime="00:04:51.97" />
                    <SPLIT distance="300" swimtime="00:05:49.43" />
                    <SPLIT distance="350" swimtime="00:06:47.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-22" firstname="Timea" gender="F" lastname="Balajcza" nation="POL" athleteid="21682">
              <RESULTS>
                <RESULT eventid="1096" points="225" reactiontime="+98" swimtime="00:03:27.10" resultid="21683" heatid="24298" lane="0" entrytime="00:03:28.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.68" />
                    <SPLIT distance="100" swimtime="00:01:41.83" />
                    <SPLIT distance="150" swimtime="00:02:37.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="206" reactiontime="+95" swimtime="00:13:40.20" resultid="21684" heatid="24311" lane="9" entrytime="00:13:46.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.03" />
                    <SPLIT distance="100" swimtime="00:01:34.08" />
                    <SPLIT distance="150" swimtime="00:02:24.19" />
                    <SPLIT distance="200" swimtime="00:03:15.66" />
                    <SPLIT distance="250" swimtime="00:04:06.70" />
                    <SPLIT distance="300" swimtime="00:04:58.54" />
                    <SPLIT distance="350" swimtime="00:05:50.51" />
                    <SPLIT distance="400" swimtime="00:06:42.93" />
                    <SPLIT distance="450" swimtime="00:07:35.71" />
                    <SPLIT distance="500" swimtime="00:08:28.98" />
                    <SPLIT distance="550" swimtime="00:09:22.26" />
                    <SPLIT distance="600" swimtime="00:10:15.35" />
                    <SPLIT distance="650" swimtime="00:11:07.09" />
                    <SPLIT distance="700" swimtime="00:11:59.04" />
                    <SPLIT distance="750" swimtime="00:12:51.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="267" reactiontime="+46" swimtime="00:03:35.79" resultid="21685" heatid="24339" lane="6" entrytime="00:03:30.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.44" />
                    <SPLIT distance="150" swimtime="00:02:41.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="201" swimtime="00:01:28.24" resultid="21686" heatid="24350" lane="8" entrytime="00:01:26.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="273" reactiontime="+79" swimtime="00:01:38.78" resultid="21687" heatid="24378" lane="3" entrytime="00:01:36.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="213" swimtime="00:03:08.92" resultid="21688" heatid="24412" lane="9" entrytime="00:03:05.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.65" />
                    <SPLIT distance="100" swimtime="00:01:32.42" />
                    <SPLIT distance="150" swimtime="00:02:20.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="301" swimtime="00:00:43.83" resultid="21689" heatid="24457" lane="8" entrytime="00:00:43.45" />
                <RESULT eventid="1721" points="198" reactiontime="+42" swimtime="00:06:45.61" resultid="21690" heatid="24471" lane="5" entrytime="00:06:15.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.98" />
                    <SPLIT distance="100" swimtime="00:01:34.58" />
                    <SPLIT distance="150" swimtime="00:02:26.00" />
                    <SPLIT distance="200" swimtime="00:03:17.77" />
                    <SPLIT distance="300" swimtime="00:05:01.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-03-14" firstname="Jarek" gender="M" lastname="Bystry" nation="POL" athleteid="21677">
              <RESULTS>
                <RESULT eventid="1079" points="390" reactiontime="+70" swimtime="00:00:28.60" resultid="21678" heatid="24292" lane="3" entrytime="00:00:28.00" />
                <RESULT eventid="1273" points="401" swimtime="00:01:03.61" resultid="21679" heatid="24362" lane="6" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="351" swimtime="00:00:31.57" resultid="21680" heatid="24395" lane="0" entrytime="00:00:31.00" />
                <RESULT eventid="1681" points="348" reactiontime="+76" swimtime="00:00:36.89" resultid="21681" heatid="24464" lane="4" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-05-02" firstname="Marcin" gender="M" lastname="Kotlarski" nation="POL" athleteid="21706">
              <RESULTS>
                <RESULT eventid="1273" points="490" swimtime="00:00:59.50" resultid="21707" heatid="24363" lane="1" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="472" reactiontime="+81" swimtime="00:02:10.94" resultid="21708" heatid="24422" lane="4" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.28" />
                    <SPLIT distance="100" swimtime="00:01:03.70" />
                    <SPLIT distance="150" swimtime="00:01:36.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="473" swimtime="00:04:42.35" resultid="21709" heatid="24480" lane="5" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.09" />
                    <SPLIT distance="150" swimtime="00:01:43.41" />
                    <SPLIT distance="200" swimtime="00:02:18.91" />
                    <SPLIT distance="250" swimtime="00:02:55.24" />
                    <SPLIT distance="300" swimtime="00:03:31.01" />
                    <SPLIT distance="350" swimtime="00:04:07.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-08" firstname="Siergiej" gender="M" lastname="Kulinicz" nation="POL" athleteid="21691">
              <RESULTS>
                <RESULT eventid="1079" points="319" reactiontime="+79" swimtime="00:00:30.59" resultid="21692" heatid="24288" lane="9" entrytime="00:00:32.06" />
                <RESULT eventid="1273" points="260" reactiontime="+72" swimtime="00:01:13.41" resultid="21693" heatid="24357" lane="4" entrytime="00:01:13.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-06-20" firstname="Tomasz" gender="M" lastname="Matras" nation="POL" athleteid="21694">
              <RESULTS>
                <RESULT eventid="1079" points="362" reactiontime="+87" swimtime="00:00:29.32" resultid="21695" heatid="24292" lane="7" entrytime="00:00:28.00" />
                <RESULT eventid="1273" points="329" swimtime="00:01:07.92" resultid="21696" heatid="24361" lane="1" entrytime="00:01:04.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-07-13" firstname="Sebastian" gender="M" lastname="Ostapczuk" nation="POL" athleteid="21710">
              <RESULTS>
                <RESULT eventid="1273" points="187" reactiontime="+42" swimtime="00:01:21.94" resultid="21711" heatid="24356" lane="0" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="195" reactiontime="+88" swimtime="00:01:38.39" resultid="21712" heatid="24382" lane="8" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="175" reactiontime="+50" swimtime="00:03:02.04" resultid="21713" heatid="24417" lane="1" entrytime="00:03:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.53" />
                    <SPLIT distance="100" swimtime="00:01:25.88" />
                    <SPLIT distance="150" swimtime="00:02:14.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="230" reactiontime="+44" swimtime="00:00:42.33" resultid="21714" heatid="24461" lane="7" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-30" firstname="Piotr" gender="M" lastname="Safrończyk" nation="POL" athleteid="21701">
              <RESULTS>
                <RESULT eventid="1079" points="639" reactiontime="+70" swimtime="00:00:24.27" resultid="21702" heatid="24296" lane="3" entrytime="00:00:24.30" />
                <RESULT eventid="1239" points="621" swimtime="00:02:28.47" resultid="21703" heatid="24346" lane="5" entrytime="00:02:32.30">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="670" reactiontime="+66" swimtime="00:01:05.23" resultid="21704" heatid="24385" lane="3" entrytime="00:01:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="708" swimtime="00:00:29.11" resultid="21705" heatid="24466" lane="2" entrytime="00:00:29.29" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1381" points="248" reactiontime="+142" swimtime="00:02:28.65" resultid="21716" heatid="24373" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.67" />
                    <SPLIT distance="100" swimtime="00:01:22.83" />
                    <SPLIT distance="150" swimtime="00:01:54.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21694" number="1" reactiontime="+142" />
                    <RELAYPOSITION athleteid="21670" number="2" />
                    <RELAYPOSITION athleteid="21677" number="3" reactiontime="+14" />
                    <RELAYPOSITION athleteid="21710" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1548" points="489" reactiontime="+64" swimtime="00:01:47.63" resultid="21717" heatid="24427" lane="7" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.35" />
                    <SPLIT distance="100" swimtime="00:00:50.71" />
                    <SPLIT distance="150" swimtime="00:01:19.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21706" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="21701" number="2" />
                    <RELAYPOSITION athleteid="21691" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="21677" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MAPOL" nation="POL" region="DOL" clubid="21222" name="KS Masters">
          <CONTACT city="Polkowice" email="bogdan.jawor@gmail.com" name="Jawor Bogdan" phone="519102742" state="DOL" street="ul.Kolejowa6/5" zip="59-100" />
          <ATHLETES>
            <ATHLETE birthdate="1941-10-02" firstname="Emilia" gender="F" lastname="Kawula" nation="POL" athleteid="21223">
              <RESULTS>
                <RESULT eventid="1062" points="21" swimtime="00:01:24.71" resultid="21224" heatid="24275" lane="2" />
                <RESULT eventid="1256" points="8" swimtime="00:04:17.59" resultid="21225" heatid="24348" lane="9" />
                <RESULT eventid="1664" points="17" swimtime="00:01:54.16" resultid="21226" heatid="24454" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-09-11" firstname="Jerzy" gender="M" lastname="Marchlewski" nation="POL" athleteid="21239">
              <RESULTS>
                <RESULT eventid="1079" points="146" reactiontime="+96" swimtime="00:00:39.70" resultid="21240" heatid="24282" lane="3" />
                <RESULT eventid="1205" points="79" swimtime="00:00:55.74" resultid="21241" heatid="24328" lane="2" />
                <RESULT eventid="1273" points="86" reactiontime="+81" swimtime="00:01:46.02" resultid="21242" heatid="24354" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="108" reactiontime="+55" swimtime="00:01:59.77" resultid="21243" heatid="24380" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="40" reactiontime="+111" swimtime="00:02:31.30" resultid="21244" heatid="24403" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="109" reactiontime="+80" swimtime="00:00:54.20" resultid="21245" heatid="24459" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-02" firstname="Pavlo" gender="M" lastname="Vechirko" nation="POL" athleteid="21232">
              <RESULTS>
                <RESULT eventid="1113" reactiontime="+104" status="DNF" swimtime="00:00:00.00" resultid="21233" heatid="24305" lane="0" entrytime="00:02:49.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="302" swimtime="00:00:35.75" resultid="21234" heatid="24333" lane="5" entrytime="00:00:34.20" entrycourse="LCM" />
                <RESULT eventid="1239" points="314" reactiontime="+71" swimtime="00:03:06.28" resultid="21235" heatid="24345" lane="0" entrytime="00:03:03.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.10" />
                    <SPLIT distance="100" swimtime="00:01:31.48" />
                    <SPLIT distance="150" swimtime="00:02:18.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="305" reactiontime="+80" swimtime="00:01:24.76" resultid="21236" heatid="24383" lane="4" entrytime="00:01:22.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="270" reactiontime="+87" swimtime="00:02:53.08" resultid="21237" heatid="24450" lane="3" entrytime="00:02:47.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.67" />
                    <SPLIT distance="100" swimtime="00:01:26.31" />
                    <SPLIT distance="150" swimtime="00:02:09.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="326" reactiontime="+93" swimtime="00:00:37.70" resultid="21238" heatid="24463" lane="3" entrytime="00:00:37.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-11-16" firstname="Gizela" gender="F" lastname="Wójcik" nation="POL" athleteid="21227">
              <RESULTS>
                <RESULT eventid="1062" points="47" swimtime="00:01:05.52" resultid="21228" heatid="24275" lane="4" />
                <RESULT eventid="1222" points="76" swimtime="00:05:27.83" resultid="21229" heatid="24338" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.42" />
                    <SPLIT distance="100" swimtime="00:02:40.19" />
                    <SPLIT distance="150" swimtime="00:04:05.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="61" swimtime="00:02:42.04" resultid="21230" heatid="24376" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="60" swimtime="00:01:14.77" resultid="21231" heatid="24453" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02001" nation="POL" region="DOL" clubid="22984" name="KS Rekin Świebodzice">
          <CONTACT city="Świebodzice" email="winiar182@wp.pl" internet="www.klubrekin.pl" name="WINIARCZYK Krzysztof" phone="606626274" state="DOL" street="Mieszka Starego 4" zip="58-160" />
          <ATHLETES>
            <ATHLETE birthdate="1986-04-20" firstname="Veronica" gender="F" lastname="Campbell-Żemier" nation="POL" athleteid="22985">
              <RESULTS>
                <RESULT eventid="1062" points="563" reactiontime="+79" swimtime="00:00:28.65" resultid="22986" heatid="24281" lane="2" entrytime="00:00:28.90" entrycourse="SCM" />
                <RESULT eventid="1222" points="428" reactiontime="+83" swimtime="00:03:04.49" resultid="22987" heatid="24340" lane="3" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.69" />
                    <SPLIT distance="100" swimtime="00:01:25.44" />
                    <SPLIT distance="150" swimtime="00:02:13.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="521" reactiontime="+41" swimtime="00:01:04.23" resultid="22988" heatid="24350" lane="7" entrytime="00:01:23.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="455" swimtime="00:01:23.37" resultid="22989" heatid="24379" lane="6" entrytime="00:01:23.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="443" swimtime="00:02:28.19" resultid="22990" heatid="24414" lane="7" entrytime="00:02:23.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                    <SPLIT distance="100" swimtime="00:01:09.13" />
                    <SPLIT distance="150" swimtime="00:01:48.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="502" swimtime="00:00:36.99" resultid="22991" heatid="24458" lane="2" entrytime="00:00:37.90" />
                <RESULT eventid="1721" points="356" reactiontime="+84" swimtime="00:05:33.59" resultid="22992" heatid="24473" lane="3" entrytime="00:04:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                    <SPLIT distance="100" swimtime="00:01:17.24" />
                    <SPLIT distance="150" swimtime="00:01:59.35" />
                    <SPLIT distance="200" swimtime="00:02:42.96" />
                    <SPLIT distance="250" swimtime="00:03:26.63" />
                    <SPLIT distance="300" swimtime="00:04:09.74" />
                    <SPLIT distance="350" swimtime="00:04:52.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-06-21" firstname="Alfred" gender="M" lastname="Żemier" nation="POL" athleteid="22993">
              <RESULTS>
                <RESULT eventid="1079" points="466" reactiontime="+79" swimtime="00:00:26.96" resultid="22994" heatid="24295" lane="3" entrytime="00:00:25.90" entrycourse="SCM" />
                <RESULT eventid="1113" points="342" reactiontime="+83" swimtime="00:02:42.89" resultid="22995" heatid="24306" lane="3" entrytime="00:02:29.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.93" />
                    <SPLIT distance="100" swimtime="00:01:14.06" />
                    <SPLIT distance="150" swimtime="00:02:03.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="423" reactiontime="+117" swimtime="00:00:31.95" resultid="22996" heatid="24334" lane="4" entrytime="00:00:31.90" />
                <RESULT eventid="1273" points="455" reactiontime="+65" swimtime="00:01:00.97" resultid="22997" heatid="24362" lane="3" entrytime="00:00:59.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="465" swimtime="00:00:28.74" resultid="22998" heatid="24396" lane="2" entrytime="00:00:28.90" />
                <RESULT eventid="1474" points="399" reactiontime="+78" swimtime="00:01:10.41" resultid="22999" heatid="24408" lane="1" entrytime="00:01:05.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="391" swimtime="00:01:08.13" resultid="23000" heatid="24441" lane="5" entrytime="00:01:03.90" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="23001" heatid="24465" lane="0" entrytime="00:00:35.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-11-09" firstname="Karol" gender="M" lastname="Żemier" nation="POL" athleteid="23002">
              <RESULTS>
                <RESULT eventid="1079" points="500" reactiontime="+82" swimtime="00:00:26.34" resultid="23003" heatid="24294" lane="0" entrytime="00:00:26.90" entrycourse="SCM" />
                <RESULT eventid="1113" points="501" reactiontime="+81" swimtime="00:02:23.52" resultid="23004" heatid="24306" lane="6" entrytime="00:02:29.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.52" />
                    <SPLIT distance="100" swimtime="00:01:06.68" />
                    <SPLIT distance="150" swimtime="00:01:48.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="552" swimtime="00:00:29.24" resultid="23005" heatid="24335" lane="5" entrytime="00:00:29.90" />
                <RESULT eventid="1341" points="392" swimtime="00:02:32.36" resultid="23006" heatid="24371" lane="1" entrytime="00:02:29.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                    <SPLIT distance="100" swimtime="00:01:09.20" />
                    <SPLIT distance="150" swimtime="00:01:49.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="519" swimtime="00:00:27.71" resultid="23007" heatid="24396" lane="6" entrytime="00:00:28.90" />
                <RESULT eventid="1474" points="515" reactiontime="+64" swimtime="00:01:04.68" resultid="23008" heatid="24408" lane="2" entrytime="00:01:03.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="489" swimtime="00:01:03.20" resultid="23009" heatid="24441" lane="4" entrytime="00:01:02.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="463" swimtime="00:02:24.63" resultid="23010" heatid="24451" lane="5" entrytime="00:02:29.90">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KS WAR" nation="POL" region="WIE" clubid="22266" name="KS Warta Poznań">
          <CONTACT city="Poznań" email="jacek.thiem@gmail.com" name="Thiem Jacek" phone="502 499 565" state="WIE" street="osiedle Dębina 19 m 34" zip="61-450" />
          <ATHLETES>
            <ATHLETE birthdate="1957-10-01" firstname="Grażyna" gender="F" lastname="Drela" nation="POL" license="500115700493" athleteid="22281">
              <RESULTS>
                <RESULT eventid="1062" points="274" reactiontime="+86" swimtime="00:00:36.44" resultid="22282" heatid="24278" lane="8" entrytime="00:00:37.00" />
                <RESULT eventid="1222" points="275" reactiontime="+83" swimtime="00:03:33.77" resultid="22283" heatid="24339" lane="2" entrytime="00:03:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.72" />
                    <SPLIT distance="100" swimtime="00:01:44.01" />
                    <SPLIT distance="150" swimtime="00:02:40.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="299" reactiontime="+65" swimtime="00:01:35.80" resultid="22284" heatid="24378" lane="6" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="296" reactiontime="+87" swimtime="00:00:44.07" resultid="22285" heatid="24456" lane="4" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-05-08" firstname="Anna" gender="F" lastname="Kotecka" nation="POL" license="100115600357" athleteid="22286">
              <RESULTS>
                <RESULT eventid="1147" points="218" swimtime="00:13:25.17" resultid="22287" heatid="24311" lane="0" entrytime="00:13:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.43" />
                    <SPLIT distance="100" swimtime="00:01:34.06" />
                    <SPLIT distance="150" swimtime="00:02:24.25" />
                    <SPLIT distance="200" swimtime="00:03:14.20" />
                    <SPLIT distance="250" swimtime="00:04:04.86" />
                    <SPLIT distance="300" swimtime="00:04:55.57" />
                    <SPLIT distance="350" swimtime="00:05:46.55" />
                    <SPLIT distance="400" swimtime="00:06:38.16" />
                    <SPLIT distance="450" swimtime="00:07:28.98" />
                    <SPLIT distance="500" swimtime="00:08:19.33" />
                    <SPLIT distance="550" swimtime="00:09:10.76" />
                    <SPLIT distance="600" swimtime="00:10:02.59" />
                    <SPLIT distance="650" swimtime="00:10:53.68" />
                    <SPLIT distance="700" swimtime="00:11:45.04" />
                    <SPLIT distance="750" swimtime="00:12:35.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="163" swimtime="00:00:49.44" resultid="22288" heatid="24324" lane="4" entrytime="00:00:50.00" />
                <RESULT eventid="1256" points="192" swimtime="00:01:29.56" resultid="22289" heatid="24350" lane="0" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="169" reactiontime="+92" swimtime="00:01:44.86" resultid="22290" heatid="24400" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="213" swimtime="00:03:09.16" resultid="22291" heatid="24411" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="184" reactiontime="+43" swimtime="00:03:38.04" resultid="22292" heatid="24443" lane="5" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:48.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="207" swimtime="00:06:39.11" resultid="22293" heatid="24471" lane="7" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.31" />
                    <SPLIT distance="100" swimtime="00:01:35.73" />
                    <SPLIT distance="150" swimtime="00:02:24.84" />
                    <SPLIT distance="200" swimtime="00:03:16.27" />
                    <SPLIT distance="250" swimtime="00:04:07.09" />
                    <SPLIT distance="300" swimtime="00:04:59.51" />
                    <SPLIT distance="350" swimtime="00:05:50.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-07-11" firstname="Waldemar" gender="M" lastname="Krakowiak" nation="POL" license="100115700335" athleteid="22317">
              <RESULTS>
                <RESULT eventid="14189" points="401" reactiontime="+65" swimtime="00:10:12.91" resultid="22318" heatid="24317" lane="6" entrytime="00:10:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                    <SPLIT distance="100" swimtime="00:01:05.79" />
                    <SPLIT distance="150" swimtime="00:01:41.27" />
                    <SPLIT distance="200" swimtime="00:02:17.69" />
                    <SPLIT distance="250" swimtime="00:02:54.75" />
                    <SPLIT distance="300" swimtime="00:03:33.28" />
                    <SPLIT distance="350" swimtime="00:04:12.13" />
                    <SPLIT distance="400" swimtime="00:04:51.09" />
                    <SPLIT distance="450" swimtime="00:05:30.13" />
                    <SPLIT distance="550" swimtime="00:06:51.37" />
                    <SPLIT distance="600" swimtime="00:08:52.72" />
                    <SPLIT distance="650" swimtime="00:08:12.64" />
                    <SPLIT distance="700" swimtime="00:10:12.91" />
                    <SPLIT distance="750" swimtime="00:09:33.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="445" swimtime="00:05:19.28" resultid="22319" heatid="24433" lane="6" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.72" />
                    <SPLIT distance="100" swimtime="00:01:04.56" />
                    <SPLIT distance="150" swimtime="00:01:47.16" />
                    <SPLIT distance="200" swimtime="00:02:30.84" />
                    <SPLIT distance="250" swimtime="00:03:15.03" />
                    <SPLIT distance="300" swimtime="00:04:00.67" />
                    <SPLIT distance="350" swimtime="00:04:40.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-05-24" firstname="Anna" gender="F" lastname="Krupińska" nation="POL" license="500115600520" athleteid="22274">
              <RESULTS>
                <RESULT eventid="1062" points="136" reactiontime="+120" swimtime="00:00:45.93" resultid="22275" heatid="24276" lane="4" entrytime="00:00:46.00" />
                <RESULT eventid="1222" points="163" reactiontime="+81" swimtime="00:04:14.56" resultid="22276" heatid="24339" lane="9" entrytime="00:04:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.57" />
                    <SPLIT distance="100" swimtime="00:02:04.55" />
                    <SPLIT distance="150" swimtime="00:03:12.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="103" reactiontime="+106" swimtime="00:01:50.25" resultid="22277" heatid="24349" lane="8" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="165" reactiontime="+94" swimtime="00:01:56.77" resultid="22278" heatid="24377" lane="2" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="103" reactiontime="+116" swimtime="00:04:00.74" resultid="22279" heatid="24410" lane="4" entrytime="00:03:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.93" />
                    <SPLIT distance="100" swimtime="00:01:57.19" />
                    <SPLIT distance="150" swimtime="00:03:01.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="172" reactiontime="+82" swimtime="00:00:52.85" resultid="22280" heatid="24456" lane="9" entrytime="00:00:52.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-07-13" firstname="Paulina" gender="F" lastname="Mendowska" nation="POL" license="100115600340" athleteid="22362">
              <RESULTS>
                <RESULT eventid="1423" points="385" reactiontime="+70" swimtime="00:00:33.57" resultid="22363" heatid="24389" lane="2" entrytime="00:00:31.30" />
                <RESULT eventid="1457" points="413" reactiontime="+84" swimtime="00:01:17.83" resultid="22364" heatid="24402" lane="2" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="360" swimtime="00:01:17.93" resultid="22365" heatid="24436" lane="5" entrytime="00:01:09.00" />
                <RESULT eventid="1630" points="396" swimtime="00:02:48.94" resultid="22366" heatid="24445" lane="6" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.89" />
                    <SPLIT distance="100" swimtime="00:01:22.97" />
                    <SPLIT distance="150" swimtime="00:02:06.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-05" firstname="Filip" gender="M" lastname="Piotrowski" nation="POL" license="500115700522" athleteid="22320">
              <RESULTS>
                <RESULT eventid="1079" points="437" reactiontime="+67" swimtime="00:00:27.55" resultid="22321" heatid="24283" lane="9" entrytime="00:01:30.00" />
                <RESULT comment="G8 - Pływak ukończył wyścig w położeniu na piersiach. (Time: 16:38), Z-3" eventid="1113" reactiontime="+70" status="DSQ" swimtime="00:02:38.59" resultid="22322" heatid="24307" lane="8" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                    <SPLIT distance="100" swimtime="00:01:14.00" />
                    <SPLIT distance="150" swimtime="00:02:03.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="453" swimtime="00:01:01.04" resultid="22323" heatid="24362" lane="4" entrytime="00:00:59.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="399" swimtime="00:00:30.23" resultid="22324" heatid="24396" lane="4" entrytime="00:00:28.53" />
                <RESULT eventid="1508" points="405" swimtime="00:02:17.81" resultid="22325" heatid="24422" lane="6" entrytime="00:02:17.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.63" />
                    <SPLIT distance="100" swimtime="00:01:08.27" />
                    <SPLIT distance="150" swimtime="00:01:44.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="410" reactiontime="+70" swimtime="00:01:07.01" resultid="22326" heatid="24441" lane="8" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="395" reactiontime="+76" swimtime="00:04:59.79" resultid="22327" heatid="24480" lane="3" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.96" />
                    <SPLIT distance="100" swimtime="00:01:14.33" />
                    <SPLIT distance="150" swimtime="00:01:52.62" />
                    <SPLIT distance="200" swimtime="00:02:32.06" />
                    <SPLIT distance="250" swimtime="00:03:09.18" />
                    <SPLIT distance="300" swimtime="00:03:46.86" />
                    <SPLIT distance="350" swimtime="00:04:24.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-12" firstname="Marcin" gender="M" lastname="Szymkowiak" nation="POL" license="500115700523" athleteid="22328">
              <RESULTS>
                <RESULT eventid="1079" points="526" reactiontime="+73" swimtime="00:00:25.90" resultid="22329" heatid="24283" lane="8" entrytime="00:01:30.00" />
                <RESULT eventid="1113" points="482" reactiontime="+70" swimtime="00:02:25.36" resultid="22330" heatid="24307" lane="9" entrytime="00:02:26.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.56" />
                    <SPLIT distance="100" swimtime="00:01:11.36" />
                    <SPLIT distance="150" swimtime="00:01:51.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="544" swimtime="00:02:35.09" resultid="22331" heatid="24346" lane="6" entrytime="00:02:37.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.38" />
                    <SPLIT distance="100" swimtime="00:01:13.77" />
                    <SPLIT distance="150" swimtime="00:01:54.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="522" swimtime="00:00:58.24" resultid="22332" heatid="24364" lane="5" entrytime="00:00:57.85" />
                <RESULT eventid="1406" points="603" swimtime="00:01:07.57" resultid="22333" heatid="24385" lane="1" entrytime="00:01:08.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="482" swimtime="00:00:28.40" resultid="22334" heatid="24397" lane="1" entrytime="00:00:28.43" />
                <RESULT eventid="1681" points="614" swimtime="00:00:30.52" resultid="22335" heatid="24466" lane="0" entrytime="00:00:31.14" />
                <RESULT eventid="1744" points="425" swimtime="00:04:52.69" resultid="22336" heatid="24481" lane="2" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                    <SPLIT distance="100" swimtime="00:01:10.45" />
                    <SPLIT distance="150" swimtime="00:01:48.26" />
                    <SPLIT distance="200" swimtime="00:02:26.38" />
                    <SPLIT distance="250" swimtime="00:03:04.57" />
                    <SPLIT distance="300" swimtime="00:03:42.62" />
                    <SPLIT distance="350" swimtime="00:04:19.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-02-17" firstname="Jacek" gender="M" lastname="Thiem" nation="POL" license="100115700345" athleteid="22267">
              <RESULTS>
                <RESULT eventid="14207" reactiontime="+116" status="OTL" swimtime="00:27:04.00" resultid="22268" heatid="24320" lane="4" entrytime="00:26:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.93" />
                    <SPLIT distance="100" swimtime="00:01:37.38" />
                    <SPLIT distance="150" swimtime="00:02:31.52" />
                    <SPLIT distance="200" swimtime="00:03:25.16" />
                    <SPLIT distance="250" swimtime="00:04:19.10" />
                    <SPLIT distance="300" swimtime="00:05:13.94" />
                    <SPLIT distance="350" swimtime="00:06:08.05" />
                    <SPLIT distance="400" swimtime="00:07:02.97" />
                    <SPLIT distance="450" swimtime="00:07:57.64" />
                    <SPLIT distance="500" swimtime="00:08:51.92" />
                    <SPLIT distance="550" swimtime="00:09:46.14" />
                    <SPLIT distance="600" swimtime="00:10:41.11" />
                    <SPLIT distance="650" swimtime="00:11:36.22" />
                    <SPLIT distance="700" swimtime="00:12:30.77" />
                    <SPLIT distance="750" swimtime="00:13:25.91" />
                    <SPLIT distance="800" swimtime="00:14:21.61" />
                    <SPLIT distance="850" swimtime="00:15:17.29" />
                    <SPLIT distance="900" swimtime="00:16:11.88" />
                    <SPLIT distance="950" swimtime="00:17:06.85" />
                    <SPLIT distance="1000" swimtime="00:18:01.63" />
                    <SPLIT distance="1050" swimtime="00:18:57.09" />
                    <SPLIT distance="1100" swimtime="00:19:53.00" />
                    <SPLIT distance="1150" swimtime="00:20:49.09" />
                    <SPLIT distance="1200" swimtime="00:21:43.86" />
                    <SPLIT distance="1250" swimtime="00:22:38.32" />
                    <SPLIT distance="1300" swimtime="00:23:33.05" />
                    <SPLIT distance="1350" swimtime="00:24:27.36" />
                    <SPLIT distance="1400" swimtime="00:25:20.32" />
                    <SPLIT distance="1450" swimtime="00:26:14.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="149" reactiontime="+98" swimtime="00:03:30.06" resultid="22269" heatid="24370" lane="0" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.70" />
                    <SPLIT distance="100" swimtime="00:01:41.74" />
                    <SPLIT distance="150" swimtime="00:02:35.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="162" reactiontime="+86" swimtime="00:00:40.80" resultid="22270" heatid="24392" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="1508" points="153" reactiontime="+85" swimtime="00:03:10.38" resultid="22271" heatid="24418" lane="1" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.54" />
                    <SPLIT distance="100" swimtime="00:01:33.36" />
                    <SPLIT distance="150" swimtime="00:02:24.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="159" reactiontime="+84" swimtime="00:01:31.91" resultid="22272" heatid="24439" lane="6" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="22273" heatid="24477" lane="2" entrytime="00:06:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-10-08" firstname="Błażej" gender="M" lastname="Wachowski" nation="POL" license="100115700545" athleteid="22354">
              <RESULTS>
                <RESULT eventid="1079" points="353" reactiontime="+84" swimtime="00:00:29.58" resultid="22355" heatid="24291" lane="4" entrytime="00:00:28.69" />
                <RESULT eventid="14189" points="320" reactiontime="+109" swimtime="00:11:00.43" resultid="22356" heatid="24317" lane="1" entrytime="00:10:29.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.09" />
                    <SPLIT distance="150" swimtime="00:01:58.20" />
                    <SPLIT distance="200" swimtime="00:02:39.40" />
                    <SPLIT distance="250" swimtime="00:03:20.70" />
                    <SPLIT distance="300" swimtime="00:04:02.74" />
                    <SPLIT distance="350" swimtime="00:04:44.94" />
                    <SPLIT distance="400" swimtime="00:05:27.27" />
                    <SPLIT distance="450" swimtime="00:06:09.26" />
                    <SPLIT distance="500" swimtime="00:06:50.05" />
                    <SPLIT distance="550" swimtime="00:07:32.89" />
                    <SPLIT distance="650" swimtime="00:08:56.98" />
                    <SPLIT distance="700" swimtime="00:09:38.25" />
                    <SPLIT distance="750" swimtime="00:10:20.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="279" reactiontime="+44" swimtime="00:02:50.59" resultid="22357" heatid="24370" lane="5" entrytime="00:02:49.30">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="317" reactiontime="+47" swimtime="00:02:29.50" resultid="22358" heatid="24421" lane="4" entrytime="00:02:22.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                    <SPLIT distance="100" swimtime="00:01:13.23" />
                    <SPLIT distance="150" swimtime="00:01:52.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="236" reactiontime="+48" swimtime="00:06:34.37" resultid="22359" heatid="24432" lane="0" entrytime="00:06:28.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                    <SPLIT distance="100" swimtime="00:01:27.80" />
                    <SPLIT distance="150" swimtime="00:02:22.58" />
                    <SPLIT distance="200" swimtime="00:05:11.28" />
                    <SPLIT distance="250" swimtime="00:04:13.47" />
                    <SPLIT distance="350" swimtime="00:05:54.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="283" reactiontime="+83" swimtime="00:01:15.83" resultid="22360" heatid="24440" lane="7" entrytime="00:01:13.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="313" reactiontime="+52" swimtime="00:05:23.80" resultid="22361" heatid="24480" lane="4" entrytime="00:05:08.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                    <SPLIT distance="100" swimtime="00:01:17.04" />
                    <SPLIT distance="150" swimtime="00:01:58.60" />
                    <SPLIT distance="200" swimtime="00:02:39.93" />
                    <SPLIT distance="250" swimtime="00:03:21.63" />
                    <SPLIT distance="300" swimtime="00:04:03.22" />
                    <SPLIT distance="350" swimtime="00:04:45.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-19" firstname="Przemysław" gender="M" lastname="Waraczewski" nation="POL" license="100115700344" athleteid="22312">
              <RESULTS>
                <RESULT eventid="1113" points="235" reactiontime="+90" swimtime="00:03:04.67" resultid="22313" heatid="24304" lane="9" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.00" />
                    <SPLIT distance="100" swimtime="00:01:31.25" />
                    <SPLIT distance="150" swimtime="00:02:22.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="267" reactiontime="+93" swimtime="00:03:16.64" resultid="22314" heatid="24344" lane="7" entrytime="00:03:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.95" />
                    <SPLIT distance="100" swimtime="00:01:32.97" />
                    <SPLIT distance="150" swimtime="00:02:25.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="245" reactiontime="+46" swimtime="00:01:31.13" resultid="22315" heatid="24383" lane="0" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="289" swimtime="00:00:39.24" resultid="22316" heatid="24462" lane="6" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-03-12" firstname="Włodzimierz" gender="M" lastname="Wiatr" nation="POL" athleteid="22303">
              <RESULTS>
                <RESULT eventid="1113" points="119" reactiontime="+111" swimtime="00:03:51.32" resultid="22304" heatid="24302" lane="2" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.05" />
                    <SPLIT distance="100" swimtime="00:01:57.88" />
                    <SPLIT distance="150" swimtime="00:03:01.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14207" points="141" reactiontime="+110" swimtime="00:27:51.74" resultid="22305" heatid="24320" lane="5" entrytime="00:27:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.05" />
                    <SPLIT distance="100" swimtime="00:01:37.88" />
                    <SPLIT distance="150" swimtime="00:02:32.41" />
                    <SPLIT distance="200" swimtime="00:03:28.11" />
                    <SPLIT distance="250" swimtime="00:04:23.38" />
                    <SPLIT distance="300" swimtime="00:05:20.16" />
                    <SPLIT distance="350" swimtime="00:06:15.13" />
                    <SPLIT distance="400" swimtime="00:07:11.85" />
                    <SPLIT distance="450" swimtime="00:08:08.08" />
                    <SPLIT distance="500" swimtime="00:09:05.21" />
                    <SPLIT distance="550" swimtime="00:10:00.92" />
                    <SPLIT distance="600" swimtime="00:10:57.69" />
                    <SPLIT distance="650" swimtime="00:11:53.03" />
                    <SPLIT distance="700" swimtime="00:12:50.09" />
                    <SPLIT distance="750" swimtime="00:13:46.75" />
                    <SPLIT distance="800" swimtime="00:14:44.29" />
                    <SPLIT distance="850" swimtime="00:15:40.34" />
                    <SPLIT distance="900" swimtime="00:16:37.08" />
                    <SPLIT distance="950" swimtime="00:17:32.86" />
                    <SPLIT distance="1000" swimtime="00:18:30.51" />
                    <SPLIT distance="1050" swimtime="00:19:26.52" />
                    <SPLIT distance="1100" swimtime="00:20:22.76" />
                    <SPLIT distance="1150" swimtime="00:21:18.16" />
                    <SPLIT distance="1200" swimtime="00:22:14.94" />
                    <SPLIT distance="1250" swimtime="00:23:11.18" />
                    <SPLIT distance="1300" swimtime="00:26:01.05" />
                    <SPLIT distance="1350" swimtime="00:25:05.47" />
                    <SPLIT distance="1450" swimtime="00:26:57.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="76" swimtime="00:00:56.48" resultid="22306" heatid="24330" lane="1" entrytime="00:00:50.25" />
                <RESULT eventid="1239" points="137" reactiontime="+109" swimtime="00:04:05.64" resultid="22307" heatid="24342" lane="4" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.81" />
                    <SPLIT distance="100" swimtime="00:01:59.36" />
                    <SPLIT distance="150" swimtime="00:03:02.31" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="M7 - Pływak wykonał naprzemienne lub nierównoczesne ruchy nóg. (Time: 16:53)" eventid="1440" reactiontime="+66" status="DSQ" swimtime="00:00:49.64" resultid="22308" heatid="24391" lane="8" entrytime="00:00:48.00" />
                <RESULT eventid="1508" points="138" reactiontime="+69" swimtime="00:03:17.17" resultid="22309" heatid="24417" lane="3" entrytime="00:03:18.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.88" />
                    <SPLIT distance="100" swimtime="00:01:35.45" />
                    <SPLIT distance="150" swimtime="00:02:27.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="22310" heatid="24447" lane="3" entrytime="00:04:20.00" />
                <RESULT eventid="1744" points="140" reactiontime="+79" swimtime="00:07:03.23" resultid="22311" heatid="24476" lane="6" entrytime="00:06:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.28" />
                    <SPLIT distance="100" swimtime="00:01:39.14" />
                    <SPLIT distance="150" swimtime="00:02:32.95" />
                    <SPLIT distance="200" swimtime="00:03:28.02" />
                    <SPLIT distance="250" swimtime="00:04:23.14" />
                    <SPLIT distance="300" swimtime="00:05:18.41" />
                    <SPLIT distance="350" swimtime="00:06:12.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-09-08" firstname="Szymon" gender="M" lastname="Wieja" nation="POL" license="500115700467" athleteid="22337">
              <RESULTS>
                <RESULT eventid="1079" points="460" reactiontime="+77" swimtime="00:00:27.08" resultid="22338" heatid="24283" lane="0" entrytime="00:01:30.00" />
                <RESULT eventid="1113" points="427" reactiontime="+82" swimtime="00:02:31.30" resultid="22339" heatid="24307" lane="1" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.21" />
                    <SPLIT distance="100" swimtime="00:01:10.95" />
                    <SPLIT distance="150" swimtime="00:01:57.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="431" swimtime="00:00:31.77" resultid="22340" heatid="24330" lane="7" entrytime="00:00:50.00" />
                <RESULT eventid="1273" points="492" swimtime="00:00:59.40" resultid="22341" heatid="24364" lane="1" entrytime="00:00:58.00" />
                <RESULT eventid="1474" points="397" reactiontime="+63" swimtime="00:01:10.50" resultid="22342" heatid="24404" lane="8" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="364" swimtime="00:02:22.81" resultid="22343" heatid="24423" lane="6" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.77" />
                    <SPLIT distance="100" swimtime="00:01:08.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="370" reactiontime="+78" swimtime="00:02:35.77" resultid="22344" heatid="24452" lane="0" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.04" />
                    <SPLIT distance="100" swimtime="00:01:16.13" />
                    <SPLIT distance="150" swimtime="00:01:56.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="362" swimtime="00:00:36.41" resultid="22345" heatid="24465" lane="2" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-10-01" firstname="Natalia" gender="F" lastname="Wiśniewska" nation="POL" license="500115600544" athleteid="22294">
              <RESULTS>
                <RESULT eventid="1096" points="531" reactiontime="+87" swimtime="00:02:35.74" resultid="22295" heatid="24299" lane="3" entrytime="00:02:37.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                    <SPLIT distance="100" swimtime="00:01:14.16" />
                    <SPLIT distance="150" swimtime="00:01:56.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="463" reactiontime="+84" swimtime="00:10:26.34" resultid="22296" heatid="24312" lane="6" entrytime="00:10:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                    <SPLIT distance="100" swimtime="00:01:13.18" />
                    <SPLIT distance="150" swimtime="00:01:52.79" />
                    <SPLIT distance="200" swimtime="00:02:32.41" />
                    <SPLIT distance="250" swimtime="00:03:11.49" />
                    <SPLIT distance="300" swimtime="00:03:51.35" />
                    <SPLIT distance="350" swimtime="00:04:30.77" />
                    <SPLIT distance="400" swimtime="00:05:10.01" />
                    <SPLIT distance="450" swimtime="00:05:50.22" />
                    <SPLIT distance="500" swimtime="00:06:29.77" />
                    <SPLIT distance="550" swimtime="00:07:09.58" />
                    <SPLIT distance="600" swimtime="00:09:08.39" />
                    <SPLIT distance="650" swimtime="00:08:28.88" />
                    <SPLIT distance="750" swimtime="00:09:48.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="555" swimtime="00:02:49.27" resultid="22297" heatid="24340" lane="5" entrytime="00:02:51.60">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="454" reactiontime="+76" swimtime="00:01:07.27" resultid="22298" heatid="24353" lane="8" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="558" reactiontime="+85" swimtime="00:01:17.88" resultid="22299" heatid="24379" lane="3" entrytime="00:01:22.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="505" reactiontime="+78" swimtime="00:05:34.38" resultid="22300" heatid="24429" lane="4" entrytime="00:05:45.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.84" />
                    <SPLIT distance="100" swimtime="00:01:13.00" />
                    <SPLIT distance="150" swimtime="00:01:59.18" />
                    <SPLIT distance="200" swimtime="00:02:43.40" />
                    <SPLIT distance="250" swimtime="00:03:28.02" />
                    <SPLIT distance="300" swimtime="00:04:13.44" />
                    <SPLIT distance="350" swimtime="00:04:54.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="559" reactiontime="+80" swimtime="00:00:35.68" resultid="22301" heatid="24458" lane="4" entrytime="00:00:34.73" />
                <RESULT eventid="1721" points="460" swimtime="00:05:06.10" resultid="22302" heatid="24473" lane="8" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                    <SPLIT distance="100" swimtime="00:01:12.82" />
                    <SPLIT distance="150" swimtime="00:01:52.08" />
                    <SPLIT distance="200" swimtime="00:02:31.84" />
                    <SPLIT distance="250" swimtime="00:03:11.45" />
                    <SPLIT distance="300" swimtime="00:03:51.31" />
                    <SPLIT distance="350" swimtime="00:04:29.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Warta Młodzi 1" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="450" reactiontime="+65" swimtime="00:02:01.89" resultid="22367" heatid="24374" lane="3" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                    <SPLIT distance="100" swimtime="00:01:03.41" />
                    <SPLIT distance="150" swimtime="00:01:33.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22337" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="22328" number="2" />
                    <RELAYPOSITION athleteid="22320" number="3" reactiontime="+6" />
                    <RELAYPOSITION athleteid="22354" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="Warta 2" number="2">
              <RESULTS>
                <RESULT eventid="1381" status="DNS" swimtime="00:00:00.00" resultid="22368" heatid="24373" lane="3" entrytime="00:02:38.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22303" number="1" />
                    <RELAYPOSITION athleteid="22312" number="2" />
                    <RELAYPOSITION athleteid="22267" number="3" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="Warta Młodzi 3" number="3">
              <RESULTS>
                <RESULT eventid="1548" points="479" swimtime="00:01:48.40" resultid="22369" heatid="24427" lane="5" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22337" number="1" />
                    <RELAYPOSITION athleteid="22320" number="2" />
                    <RELAYPOSITION athleteid="22354" number="3" />
                    <RELAYPOSITION athleteid="22328" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="Warta 4" number="4">
              <RESULTS>
                <RESULT eventid="1548" status="DNS" swimtime="00:00:00.00" resultid="22370" heatid="24426" lane="6" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.29" />
                    <SPLIT distance="100" swimtime="00:01:03.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22303" number="1" />
                    <RELAYPOSITION athleteid="22312" number="2" />
                    <RELAYPOSITION athleteid="22267" number="3" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Warta 5 mixed dow" number="5">
              <RESULTS>
                <RESULT eventid="1130" swimtime="00:02:33.50" resultid="22371" heatid="24308" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.65" />
                    <SPLIT distance="100" swimtime="00:01:22.07" />
                    <SPLIT distance="150" swimtime="00:01:59.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22286" number="1" />
                    <RELAYPOSITION athleteid="22281" number="2" />
                    <RELAYPOSITION athleteid="22267" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="22312" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" name="Warta 5 mixed dow" number="6">
              <RESULTS>
                <RESULT eventid="1698" reactiontime="+45" swimtime="00:02:50.61" resultid="22372" heatid="24468" lane="9" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.37" />
                    <SPLIT distance="100" swimtime="00:01:33.78" />
                    <SPLIT distance="150" swimtime="00:02:17.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22286" number="1" reactiontime="+45" />
                    <RELAYPOSITION athleteid="22281" number="2" />
                    <RELAYPOSITION athleteid="22267" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="22312" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="NZWAW" nation="POL" region="WA" clubid="20689" name="KS_Niezrzeszeni_pl">
          <CONTACT name="KS_Niezrzeszeni_pl" />
          <ATHLETES>
            <ATHLETE birthdate="1959-12-27" firstname="Wojciech" gender="M" lastname="Korpetta" nation="POL" athleteid="20690">
              <RESULTS>
                <RESULT eventid="1079" points="196" reactiontime="+114" swimtime="00:00:35.99" resultid="20691" heatid="24286" lane="0" entrytime="00:00:35.13" />
                <RESULT eventid="14189" points="190" reactiontime="+103" swimtime="00:13:05.94" resultid="20692" heatid="24315" lane="7" entrytime="00:12:54.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.75" />
                    <SPLIT distance="100" swimtime="00:01:31.53" />
                    <SPLIT distance="150" swimtime="00:02:21.88" />
                    <SPLIT distance="200" swimtime="00:03:12.84" />
                    <SPLIT distance="250" swimtime="00:04:04.02" />
                    <SPLIT distance="300" swimtime="00:04:55.38" />
                    <SPLIT distance="350" swimtime="00:05:46.49" />
                    <SPLIT distance="400" swimtime="00:06:37.34" />
                    <SPLIT distance="450" swimtime="00:07:28.10" />
                    <SPLIT distance="500" swimtime="00:08:18.56" />
                    <SPLIT distance="550" swimtime="00:09:08.91" />
                    <SPLIT distance="650" swimtime="00:10:48.86" />
                    <SPLIT distance="700" swimtime="00:09:59.07" />
                    <SPLIT distance="750" swimtime="00:12:24.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="200" reactiontime="+60" swimtime="00:01:20.20" resultid="20693" heatid="24357" lane="0" entrytime="00:01:18.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="178" reactiontime="+98" swimtime="00:03:01.17" resultid="20694" heatid="24418" lane="5" entrytime="00:02:58.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.51" />
                    <SPLIT distance="100" swimtime="00:01:30.02" />
                    <SPLIT distance="150" swimtime="00:02:17.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="177" reactiontime="+70" swimtime="00:03:19.20" resultid="20695" heatid="24449" lane="1" entrytime="00:03:12.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:30.01" />
                    <SPLIT distance="100" swimtime="00:01:38.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="180" reactiontime="+74" swimtime="00:06:29.06" resultid="20696" heatid="24477" lane="3" entrytime="00:06:23.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.87" />
                    <SPLIT distance="100" swimtime="00:01:33.82" />
                    <SPLIT distance="150" swimtime="00:02:25.12" />
                    <SPLIT distance="200" swimtime="00:03:16.93" />
                    <SPLIT distance="250" swimtime="00:04:07.23" />
                    <SPLIT distance="350" swimtime="00:05:45.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="039" nation="POL" region="SLA" clubid="20765" name="KU AZS PWSZ Racibórz">
          <CONTACT city="Racibórz" email="m.kunicki@vp.pl" name="Kunicki Marcin" phone="504233267" state="ŚLĄSK" street="Słowackiego 55" zip="47-400" />
          <ATHLETES>
            <ATHLETE birthdate="1998-06-14" firstname="Wiktoria" gender="F" lastname="Kolbe" nation="POL" license="103911600023" athleteid="20766">
              <RESULTS>
                <RESULT eventid="1062" points="558" reactiontime="+82" swimtime="00:00:28.74" resultid="20767" heatid="24281" lane="7" entrytime="00:00:29.00" entrycourse="LCM" />
                <RESULT eventid="1256" points="506" reactiontime="+74" swimtime="00:01:04.87" resultid="20768" heatid="24353" lane="7" entrytime="00:01:05.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="552" swimtime="00:00:29.78" resultid="20769" heatid="24389" lane="5" entrytime="00:00:29.50" entrycourse="LCM" />
                <RESULT eventid="1595" points="411" reactiontime="+41" swimtime="00:01:14.61" resultid="20770" heatid="24436" lane="2" entrytime="00:01:12.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="556" swimtime="00:00:35.74" resultid="20771" heatid="24458" lane="5" entrytime="00:00:36.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-10-02" firstname="Agnieszka" gender="F" lastname="Ostrowska" nation="POL" license="103911600016" athleteid="20774">
              <RESULTS>
                <RESULT eventid="1096" points="606" reactiontime="+76" swimtime="00:02:28.98" resultid="20775" heatid="24299" lane="5" entrytime="00:02:35.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="618" reactiontime="+78" swimtime="00:02:43.26" resultid="20776" heatid="24340" lane="4" entrytime="00:02:44.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                    <SPLIT distance="100" swimtime="00:01:18.84" />
                    <SPLIT distance="150" swimtime="00:02:00.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="629" reactiontime="+76" swimtime="00:01:14.82" resultid="20777" heatid="24379" lane="4" entrytime="00:01:18.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-02-24" firstname="Maciej" gender="M" lastname="Sudenis" nation="POL" license="103911700019" athleteid="20772">
              <RESULTS>
                <RESULT eventid="1079" points="494" reactiontime="+72" swimtime="00:00:26.45" resultid="20773" heatid="24295" lane="7" entrytime="00:00:26.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LCGW" nation="POL" region="LBS" clubid="20679" name="LC Gorzów Wlkp.">
          <CONTACT city="Os. Poznanskie" email="stan_ley@poczta.fm" name="Kaczmarek" phone="600277732" state="LUBUS" street="Liliowa" street2="9" zip="66-446" />
          <ATHLETES>
            <ATHLETE birthdate="1979-01-26" firstname="Stanislaw" gender="M" lastname="Kaczmarek" nation="POL" athleteid="20680">
              <RESULTS>
                <RESULT eventid="1113" points="483" reactiontime="+79" swimtime="00:02:25.26" resultid="20681" heatid="24307" lane="2" entrytime="00:02:23.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.21" />
                    <SPLIT distance="100" swimtime="00:01:09.82" />
                    <SPLIT distance="150" swimtime="00:01:51.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14189" points="462" reactiontime="+75" swimtime="00:09:44.58" resultid="20682" heatid="24317" lane="5" entrytime="00:09:20.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.18" />
                    <SPLIT distance="100" swimtime="00:01:08.87" />
                    <SPLIT distance="150" swimtime="00:01:55.22" />
                    <SPLIT distance="200" swimtime="00:02:21.31" />
                    <SPLIT distance="250" swimtime="00:02:58.06" />
                    <SPLIT distance="300" swimtime="00:03:35.17" />
                    <SPLIT distance="350" swimtime="00:04:12.03" />
                    <SPLIT distance="400" swimtime="00:04:49.54" />
                    <SPLIT distance="450" swimtime="00:05:26.54" />
                    <SPLIT distance="500" swimtime="00:06:04.03" />
                    <SPLIT distance="550" swimtime="00:06:41.44" />
                    <SPLIT distance="600" swimtime="00:07:18.72" />
                    <SPLIT distance="650" swimtime="00:07:55.43" />
                    <SPLIT distance="700" swimtime="00:08:32.39" />
                    <SPLIT distance="750" swimtime="00:09:08.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="441" reactiontime="+65" swimtime="00:02:46.35" resultid="20683" heatid="24346" lane="7" entrytime="00:02:43.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                    <SPLIT distance="100" swimtime="00:01:20.31" />
                    <SPLIT distance="150" swimtime="00:02:03.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="409" reactiontime="+72" swimtime="00:02:30.22" resultid="20684" heatid="24371" lane="2" entrytime="00:02:21.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                    <SPLIT distance="100" swimtime="00:01:11.46" />
                    <SPLIT distance="150" swimtime="00:01:51.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="466" swimtime="00:02:11.49" resultid="20685" heatid="24424" lane="9" entrytime="00:02:07.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.78" />
                    <SPLIT distance="100" swimtime="00:01:04.06" />
                    <SPLIT distance="150" swimtime="00:01:37.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="455" reactiontime="+43" swimtime="00:05:16.84" resultid="20686" heatid="24433" lane="3" entrytime="00:05:09.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.41" />
                    <SPLIT distance="100" swimtime="00:01:08.37" />
                    <SPLIT distance="150" swimtime="00:01:53.01" />
                    <SPLIT distance="200" swimtime="00:02:36.50" />
                    <SPLIT distance="250" swimtime="00:03:21.38" />
                    <SPLIT distance="300" swimtime="00:04:07.64" />
                    <SPLIT distance="350" swimtime="00:04:43.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="449" swimtime="00:01:05.04" resultid="20687" heatid="24442" lane="0" entrytime="00:01:02.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="483" swimtime="00:04:40.42" resultid="20688" heatid="24482" lane="6" entrytime="00:04:29.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.47" />
                    <SPLIT distance="100" swimtime="00:01:06.17" />
                    <SPLIT distance="150" swimtime="00:01:41.53" />
                    <SPLIT distance="200" swimtime="00:02:17.57" />
                    <SPLIT distance="250" swimtime="00:02:53.16" />
                    <SPLIT distance="300" swimtime="00:03:29.68" />
                    <SPLIT distance="350" swimtime="00:04:05.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="MAZ" clubid="21566" name="Legia Warszawa">
          <CONTACT email="agnieszka.kaczmarek85@gmail.com" name="Kaczmarek" phone="531799855" />
          <ATHLETES>
            <ATHLETE birthdate="1953-05-05" firstname="Bogdan" gender="M" lastname="Dubiński" nation="POL" athleteid="23426">
              <RESULTS>
                <RESULT eventid="1079" points="218" reactiontime="+99" swimtime="00:00:34.71" resultid="23427" heatid="24287" lane="0" entrytime="00:00:34.00" />
                <RESULT eventid="14189" points="175" reactiontime="+103" swimtime="00:13:27.64" resultid="23428" heatid="24314" lane="3" entrytime="00:15:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.33" />
                    <SPLIT distance="100" swimtime="00:01:28.15" />
                    <SPLIT distance="150" swimtime="00:02:19.16" />
                    <SPLIT distance="200" swimtime="00:03:11.22" />
                    <SPLIT distance="250" swimtime="00:04:02.33" />
                    <SPLIT distance="300" swimtime="00:04:54.94" />
                    <SPLIT distance="350" swimtime="00:05:47.09" />
                    <SPLIT distance="400" swimtime="00:06:40.16" />
                    <SPLIT distance="450" swimtime="00:07:32.38" />
                    <SPLIT distance="500" swimtime="00:08:25.34" />
                    <SPLIT distance="550" swimtime="00:09:17.46" />
                    <SPLIT distance="600" swimtime="00:10:09.07" />
                    <SPLIT distance="650" swimtime="00:11:00.36" />
                    <SPLIT distance="700" swimtime="00:11:51.51" />
                    <SPLIT distance="750" swimtime="00:12:41.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="211" swimtime="00:00:40.27" resultid="23429" heatid="24331" lane="3" entrytime="00:00:43.00" />
                <RESULT eventid="1341" points="78" reactiontime="+69" swimtime="00:04:20.71" resultid="23430" heatid="24369" lane="9" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.56" />
                    <SPLIT distance="100" swimtime="00:02:04.78" />
                    <SPLIT distance="150" swimtime="00:03:14.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="170" reactiontime="+84" swimtime="00:01:33.59" resultid="23431" heatid="24405" lane="9" entrytime="00:01:34.00" />
                <RESULT eventid="1578" points="134" reactiontime="+95" swimtime="00:07:55.58" resultid="23432" heatid="24431" lane="8" entrytime="00:07:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.78" />
                    <SPLIT distance="100" swimtime="00:02:04.43" />
                    <SPLIT distance="150" swimtime="00:03:04.54" />
                    <SPLIT distance="200" swimtime="00:04:03.29" />
                    <SPLIT distance="250" swimtime="00:05:15.30" />
                    <SPLIT distance="300" swimtime="00:06:23.20" />
                    <SPLIT distance="350" swimtime="00:07:12.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="153" swimtime="00:03:28.98" resultid="23433" heatid="24448" lane="6" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.87" />
                    <SPLIT distance="100" swimtime="00:01:44.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="170" reactiontime="+61" swimtime="00:06:37.11" resultid="23434" heatid="24477" lane="0" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.80" />
                    <SPLIT distance="100" swimtime="00:01:31.33" />
                    <SPLIT distance="150" swimtime="00:02:24.07" />
                    <SPLIT distance="200" swimtime="00:03:18.17" />
                    <SPLIT distance="250" swimtime="00:04:10.62" />
                    <SPLIT distance="300" swimtime="00:05:01.59" />
                    <SPLIT distance="350" swimtime="00:05:51.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-08-13" firstname="Romuald" gender="M" lastname="Kozlowski" nation="POL" athleteid="21571">
              <RESULTS>
                <RESULT eventid="1079" points="379" reactiontime="+79" swimtime="00:00:28.87" resultid="21572" heatid="24291" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="1239" points="355" reactiontime="+51" swimtime="00:02:58.79" resultid="21573" heatid="24341" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.34" />
                    <SPLIT distance="100" swimtime="00:01:24.23" />
                    <SPLIT distance="150" swimtime="00:02:10.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="351" reactiontime="+45" swimtime="00:01:20.90" resultid="21574" heatid="24384" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="21575" heatid="24396" lane="7" entrytime="00:00:29.00" />
                <RESULT eventid="1681" points="413" reactiontime="+43" swimtime="00:00:34.83" resultid="21576" heatid="24464" lane="2" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-04" firstname="Hubert" gender="M" lastname="Markowski" nation="POL" athleteid="21577">
              <RESULTS>
                <RESULT eventid="1113" points="376" reactiontime="+78" swimtime="00:02:37.87" resultid="21578" heatid="24305" lane="5" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                    <SPLIT distance="100" swimtime="00:01:15.62" />
                    <SPLIT distance="150" swimtime="00:02:01.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" status="DNS" swimtime="00:00:00.00" resultid="21579" heatid="24371" lane="9" entrytime="00:02:38.00" />
                <RESULT eventid="1474" points="342" reactiontime="+74" swimtime="00:01:14.14" resultid="21580" heatid="24407" lane="1" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="340" reactiontime="+73" swimtime="00:05:49.25" resultid="21581" heatid="24432" lane="7" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                    <SPLIT distance="100" swimtime="00:01:21.43" />
                    <SPLIT distance="150" swimtime="00:02:07.49" />
                    <SPLIT distance="200" swimtime="00:02:52.16" />
                    <SPLIT distance="250" swimtime="00:03:41.77" />
                    <SPLIT distance="300" swimtime="00:04:31.77" />
                    <SPLIT distance="350" swimtime="00:05:11.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="400" swimtime="00:01:07.61" resultid="21582" heatid="24440" lane="4" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="325" reactiontime="+119" swimtime="00:02:42.77" resultid="21583" heatid="24450" lane="4" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.89" />
                    <SPLIT distance="100" swimtime="00:01:21.06" />
                    <SPLIT distance="150" swimtime="00:02:02.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-07-12" firstname="Filip" gender="M" lastname="Rowinski" nation="POL" athleteid="21567">
              <RESULTS>
                <RESULT eventid="1406" points="521" swimtime="00:01:10.96" resultid="21568" heatid="24385" lane="6" entrytime="00:01:06.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="534" swimtime="00:00:27.44" resultid="21569" heatid="24398" lane="9" entrytime="00:00:26.99" />
                <RESULT eventid="1681" points="606" reactiontime="+65" swimtime="00:00:30.66" resultid="21570" heatid="24466" lane="7" entrytime="00:00:29.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-11-23" firstname="Katarzyna" gender="F" lastname="Żołnowska" nation="POL" athleteid="21584">
              <RESULTS>
                <RESULT eventid="1165" points="519" reactiontime="+82" swimtime="00:19:05.39" resultid="21585" heatid="24319" lane="4" entrytime="00:18:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                    <SPLIT distance="100" swimtime="00:01:09.64" />
                    <SPLIT distance="150" swimtime="00:01:46.94" />
                    <SPLIT distance="200" swimtime="00:02:24.75" />
                    <SPLIT distance="250" swimtime="00:03:03.24" />
                    <SPLIT distance="300" swimtime="00:03:41.58" />
                    <SPLIT distance="350" swimtime="00:04:20.64" />
                    <SPLIT distance="400" swimtime="00:04:59.29" />
                    <SPLIT distance="450" swimtime="00:05:37.87" />
                    <SPLIT distance="500" swimtime="00:06:15.86" />
                    <SPLIT distance="550" swimtime="00:06:54.19" />
                    <SPLIT distance="600" swimtime="00:07:32.64" />
                    <SPLIT distance="650" swimtime="00:08:11.39" />
                    <SPLIT distance="700" swimtime="00:08:49.57" />
                    <SPLIT distance="750" swimtime="00:09:28.27" />
                    <SPLIT distance="800" swimtime="00:10:06.64" />
                    <SPLIT distance="850" swimtime="00:10:45.58" />
                    <SPLIT distance="900" swimtime="00:11:24.25" />
                    <SPLIT distance="950" swimtime="00:12:03.25" />
                    <SPLIT distance="1000" swimtime="00:12:41.63" />
                    <SPLIT distance="1050" swimtime="00:13:20.40" />
                    <SPLIT distance="1100" swimtime="00:13:58.82" />
                    <SPLIT distance="1150" swimtime="00:14:37.82" />
                    <SPLIT distance="1200" swimtime="00:15:16.26" />
                    <SPLIT distance="1250" swimtime="00:15:55.47" />
                    <SPLIT distance="1300" swimtime="00:16:33.75" />
                    <SPLIT distance="1350" swimtime="00:17:12.95" />
                    <SPLIT distance="1400" swimtime="00:17:51.77" />
                    <SPLIT distance="1450" swimtime="00:18:29.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="552" swimtime="00:01:03.02" resultid="21586" heatid="24353" lane="5" entrytime="00:01:01.00" />
                <RESULT eventid="1491" points="562" swimtime="00:02:16.83" resultid="21587" heatid="24414" lane="5" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="517" reactiontime="+84" swimtime="00:04:54.50" resultid="21588" heatid="24473" lane="4" entrytime="00:04:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.08" />
                    <SPLIT distance="100" swimtime="00:01:10.13" />
                    <SPLIT distance="150" swimtime="00:01:47.26" />
                    <SPLIT distance="200" swimtime="00:02:25.34" />
                    <SPLIT distance="250" swimtime="00:03:03.54" />
                    <SPLIT distance="300" swimtime="00:03:41.45" />
                    <SPLIT distance="350" swimtime="00:04:18.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="20250" name="Masters Białystok">
          <CONTACT email="mbzgloszenia@gmail.com" name="DM" />
          <ATHLETES>
            <ATHLETE birthdate="1979-01-01" firstname="Dominika" gender="F" lastname="Michalik" nation="POL" athleteid="20257">
              <RESULTS>
                <RESULT eventid="1147" points="442" reactiontime="+83" swimtime="00:10:36.32" resultid="20258" heatid="24312" lane="5" entrytime="00:10:24.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                    <SPLIT distance="100" swimtime="00:01:12.05" />
                    <SPLIT distance="150" swimtime="00:01:51.71" />
                    <SPLIT distance="200" swimtime="00:02:31.45" />
                    <SPLIT distance="250" swimtime="00:03:11.59" />
                    <SPLIT distance="300" swimtime="00:03:51.19" />
                    <SPLIT distance="350" swimtime="00:04:31.44" />
                    <SPLIT distance="400" swimtime="00:05:11.75" />
                    <SPLIT distance="450" swimtime="00:05:52.08" />
                    <SPLIT distance="500" swimtime="00:06:32.22" />
                    <SPLIT distance="550" swimtime="00:07:13.08" />
                    <SPLIT distance="600" swimtime="00:07:53.25" />
                    <SPLIT distance="650" swimtime="00:08:34.32" />
                    <SPLIT distance="700" swimtime="00:09:15.59" />
                    <SPLIT distance="750" swimtime="00:09:56.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="501" swimtime="00:01:05.08" resultid="20259" heatid="24353" lane="1" entrytime="00:01:05.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="501" reactiontime="+72" swimtime="00:02:22.24" resultid="20260" heatid="24414" lane="2" entrytime="00:02:22.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.93" />
                    <SPLIT distance="100" swimtime="00:01:08.83" />
                    <SPLIT distance="150" swimtime="00:01:45.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="472" reactiontime="+74" swimtime="00:05:03.59" resultid="20261" heatid="24473" lane="7" entrytime="00:05:01.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                    <SPLIT distance="100" swimtime="00:01:12.28" />
                    <SPLIT distance="150" swimtime="00:01:50.62" />
                    <SPLIT distance="200" swimtime="00:02:29.26" />
                    <SPLIT distance="250" swimtime="00:03:07.90" />
                    <SPLIT distance="300" swimtime="00:03:46.52" />
                    <SPLIT distance="350" swimtime="00:04:25.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-01-01" firstname="Andrzej" gender="M" lastname="Twarowski" nation="POL" athleteid="20251">
              <RESULTS>
                <RESULT eventid="14207" reactiontime="+103" status="OTL" swimtime="00:25:30.91" resultid="20252" heatid="24321" lane="7" entrytime="00:25:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.58" />
                    <SPLIT distance="100" swimtime="00:01:32.59" />
                    <SPLIT distance="150" swimtime="00:02:23.51" />
                    <SPLIT distance="200" swimtime="00:03:15.48" />
                    <SPLIT distance="250" swimtime="00:04:07.34" />
                    <SPLIT distance="300" swimtime="00:04:59.76" />
                    <SPLIT distance="350" swimtime="00:05:51.72" />
                    <SPLIT distance="400" swimtime="00:06:44.89" />
                    <SPLIT distance="450" swimtime="00:07:36.44" />
                    <SPLIT distance="500" swimtime="00:08:27.97" />
                    <SPLIT distance="550" swimtime="00:09:19.94" />
                    <SPLIT distance="600" swimtime="00:10:12.00" />
                    <SPLIT distance="650" swimtime="00:11:04.71" />
                    <SPLIT distance="700" swimtime="00:11:56.95" />
                    <SPLIT distance="750" swimtime="00:12:49.06" />
                    <SPLIT distance="800" swimtime="00:13:39.33" />
                    <SPLIT distance="850" swimtime="00:14:31.35" />
                    <SPLIT distance="900" swimtime="00:15:22.95" />
                    <SPLIT distance="950" swimtime="00:16:14.45" />
                    <SPLIT distance="1000" swimtime="00:17:05.21" />
                    <SPLIT distance="1050" swimtime="00:17:57.29" />
                    <SPLIT distance="1100" swimtime="00:18:49.21" />
                    <SPLIT distance="1150" swimtime="00:19:41.29" />
                    <SPLIT distance="1200" swimtime="00:20:32.16" />
                    <SPLIT distance="1250" swimtime="00:21:24.66" />
                    <SPLIT distance="1300" swimtime="00:22:14.83" />
                    <SPLIT distance="1350" swimtime="00:23:06.12" />
                    <SPLIT distance="1400" swimtime="00:23:56.20" />
                    <SPLIT distance="1450" swimtime="00:24:45.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="207" reactiontime="+72" swimtime="00:03:34.04" resultid="20253" heatid="24343" lane="3" entrytime="00:03:29.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.72" />
                    <SPLIT distance="100" swimtime="00:01:41.32" />
                    <SPLIT distance="150" swimtime="00:02:37.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="122" reactiontime="+65" swimtime="00:03:44.83" resultid="20254" heatid="24369" lane="5" entrytime="00:03:42.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:50.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="163" reactiontime="+78" swimtime="00:07:26.28" resultid="20255" heatid="24431" lane="3" entrytime="00:07:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.78" />
                    <SPLIT distance="100" swimtime="00:01:48.57" />
                    <SPLIT distance="150" swimtime="00:02:44.01" />
                    <SPLIT distance="200" swimtime="00:03:40.05" />
                    <SPLIT distance="250" swimtime="00:04:40.32" />
                    <SPLIT distance="300" swimtime="00:05:41.93" />
                    <SPLIT distance="350" swimtime="00:06:35.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="169" swimtime="00:03:22.19" resultid="20256" heatid="24449" lane="8" entrytime="00:03:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.54" />
                    <SPLIT distance="100" swimtime="00:01:40.10" />
                    <SPLIT distance="150" swimtime="00:02:34.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LUB" nation="POL" region="LBL" clubid="22239" name="MASTERS Lublin">
          <CONTACT city="Lublin" email="masters_lublin@wp.pl" name="Wójcicki" phone="+48501794954" state="LUBEL" street="Stanisława Lema 18" zip="20-445" />
          <ATHLETES>
            <ATHLETE birthdate="1975-05-28" firstname="Anna" gender="F" lastname="Michalska" nation="POL" license="103503600002" athleteid="22255">
              <RESULTS>
                <RESULT eventid="1096" points="277" reactiontime="+105" swimtime="00:03:13.47" resultid="22256" heatid="24298" lane="2" entrytime="00:03:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.29" />
                    <SPLIT distance="100" swimtime="00:01:29.47" />
                    <SPLIT distance="150" swimtime="00:02:24.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="345" swimtime="00:00:38.57" resultid="22257" heatid="24326" lane="2" entrytime="00:00:38.09" entrycourse="LCM" />
                <RESULT eventid="1457" points="329" reactiontime="+93" swimtime="00:01:23.95" resultid="22258" heatid="24401" lane="5" entrytime="00:01:22.01" entrycourse="LCM" />
                <RESULT eventid="1630" points="296" reactiontime="+91" swimtime="00:03:06.03" resultid="22259" heatid="24445" lane="0" entrytime="00:03:01.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.31" />
                    <SPLIT distance="100" swimtime="00:01:28.27" />
                    <SPLIT distance="150" swimtime="00:02:17.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-12-11" firstname="Mirosław" gender="M" lastname="Molenda" nation="POL" license="103503700012" athleteid="22249">
              <RESULTS>
                <RESULT eventid="14189" reactiontime="+153" status="OTL" swimtime="00:13:31.91" resultid="22250" heatid="24315" lane="0" entrytime="00:13:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.61" />
                    <SPLIT distance="100" swimtime="00:01:26.38" />
                    <SPLIT distance="150" swimtime="00:02:15.56" />
                    <SPLIT distance="200" swimtime="00:03:06.90" />
                    <SPLIT distance="250" swimtime="00:03:57.91" />
                    <SPLIT distance="300" swimtime="00:04:50.38" />
                    <SPLIT distance="350" swimtime="00:05:42.17" />
                    <SPLIT distance="400" swimtime="00:06:35.58" />
                    <SPLIT distance="450" swimtime="00:07:28.36" />
                    <SPLIT distance="500" swimtime="00:08:21.64" />
                    <SPLIT distance="550" swimtime="00:09:14.58" />
                    <SPLIT distance="600" swimtime="00:10:07.75" />
                    <SPLIT distance="700" swimtime="00:11:53.30" />
                    <SPLIT distance="750" swimtime="00:12:45.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-10-21" firstname="Adam" gender="M" lastname="Pietrzak" nation="POL" license="103503700011" athleteid="22243">
              <RESULTS>
                <RESULT eventid="1079" points="318" reactiontime="+89" swimtime="00:00:30.63" resultid="22244" heatid="24288" lane="5" entrytime="00:00:31.17" entrycourse="LCM" />
                <RESULT eventid="1239" points="288" reactiontime="+76" swimtime="00:03:11.70" resultid="22245" heatid="24345" lane="3" entrytime="00:02:58.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.25" />
                    <SPLIT distance="100" swimtime="00:01:29.79" />
                    <SPLIT distance="150" swimtime="00:02:21.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="296" reactiontime="+74" swimtime="00:01:25.64" resultid="22246" heatid="24383" lane="3" entrytime="00:01:24.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="275" reactiontime="+69" swimtime="00:01:19.70" resultid="22247" heatid="24406" lane="9" entrytime="00:01:22.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="228" reactiontime="+90" swimtime="00:03:03.05" resultid="22248" heatid="24450" lane="1" entrytime="00:02:53.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.99" />
                    <SPLIT distance="100" swimtime="00:01:30.05" />
                    <SPLIT distance="150" swimtime="00:02:18.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-04-28" firstname="Rafał" gender="M" lastname="Wójcicki" nation="POL" license="103503700001" athleteid="22251">
              <RESULTS>
                <RESULT eventid="1205" points="241" swimtime="00:00:38.54" resultid="22252" heatid="24333" lane="0" entrytime="00:00:36.88" entrycourse="LCM" />
                <RESULT eventid="1474" points="250" reactiontime="+78" swimtime="00:01:22.24" resultid="22253" heatid="24406" lane="0" entrytime="00:01:20.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="273" swimtime="00:00:40.00" resultid="22254" heatid="24462" lane="5" entrytime="00:00:40.32" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-11-07" firstname="Konrad" gender="M" lastname="Ćwikła" nation="POL" license="103503700005" athleteid="22240">
              <RESULTS>
                <RESULT eventid="1273" points="344" swimtime="00:01:06.92" resultid="22241" heatid="24359" lane="7" entrytime="00:01:08.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="262" reactiontime="+88" swimtime="00:02:39.29" resultid="22242" heatid="24420" lane="7" entrytime="00:02:35.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.27" />
                    <SPLIT distance="150" swimtime="00:01:58.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="20915" name="Masters V Łomianki">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1964-03-12" firstname="Robert" gender="M" lastname="Dziudziek" nation="POL" athleteid="20916">
              <RESULTS>
                <RESULT eventid="14189" points="217" reactiontime="+119" swimtime="00:12:31.87" resultid="20917" heatid="24315" lane="4" entrytime="00:12:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.16" />
                    <SPLIT distance="100" swimtime="00:01:26.41" />
                    <SPLIT distance="150" swimtime="00:02:12.34" />
                    <SPLIT distance="200" swimtime="00:02:58.17" />
                    <SPLIT distance="250" swimtime="00:03:44.46" />
                    <SPLIT distance="300" swimtime="00:04:31.05" />
                    <SPLIT distance="350" swimtime="00:05:17.78" />
                    <SPLIT distance="400" swimtime="00:06:05.41" />
                    <SPLIT distance="450" swimtime="00:06:52.77" />
                    <SPLIT distance="500" swimtime="00:07:41.00" />
                    <SPLIT distance="550" swimtime="00:08:29.32" />
                    <SPLIT distance="600" swimtime="00:09:17.58" />
                    <SPLIT distance="650" swimtime="00:10:06.33" />
                    <SPLIT distance="700" swimtime="00:10:54.80" />
                    <SPLIT distance="750" swimtime="00:11:43.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="115" reactiontime="+101" swimtime="00:03:48.73" resultid="20918" heatid="24369" lane="4" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.51" />
                    <SPLIT distance="100" swimtime="00:01:46.95" />
                    <SPLIT distance="150" swimtime="00:02:47.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="20919" heatid="24420" lane="5" entrytime="00:02:35.00" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="20920" heatid="24438" lane="4" entrytime="00:01:35.00" />
                <RESULT eventid="1744" points="241" reactiontime="+77" swimtime="00:05:53.21" resultid="20921" heatid="24479" lane="1" entrytime="00:05:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                    <SPLIT distance="100" swimtime="00:01:22.04" />
                    <SPLIT distance="150" swimtime="00:02:05.77" />
                    <SPLIT distance="200" swimtime="00:02:50.97" />
                    <SPLIT distance="250" swimtime="00:03:35.96" />
                    <SPLIT distance="300" swimtime="00:04:21.77" />
                    <SPLIT distance="350" swimtime="00:05:07.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WIKRA" nation="POL" region="MAL" clubid="20697" name="Masters Wisła Kraków">
          <CONTACT email="wislaplywanie@gmail.com" internet="http://www.wislaplywanie.pl/sekcja-masters/" name="Tomasz Doniec" phone="693703490" />
          <ATHLETES>
            <ATHLETE birthdate="1957-02-26" firstname="Iwona" gender="F" lastname="Bednarczyk" nation="POL" license="501806600060" athleteid="20706">
              <RESULTS>
                <RESULT eventid="1096" points="67" reactiontime="+112" swimtime="00:05:10.39" resultid="20707" heatid="24297" lane="2" entrytime="00:04:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.03" />
                    <SPLIT distance="100" swimtime="00:02:38.71" />
                    <SPLIT distance="150" swimtime="00:03:57.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" status="OTL" swimtime="00:37:13.19" resultid="20708" heatid="24318" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.91" />
                    <SPLIT distance="100" swimtime="00:02:04.92" />
                    <SPLIT distance="150" swimtime="00:03:16.42" />
                    <SPLIT distance="200" swimtime="00:04:30.33" />
                    <SPLIT distance="250" swimtime="00:05:42.09" />
                    <SPLIT distance="300" swimtime="00:06:55.82" />
                    <SPLIT distance="350" swimtime="00:08:10.02" />
                    <SPLIT distance="400" swimtime="00:09:23.46" />
                    <SPLIT distance="450" swimtime="00:10:35.98" />
                    <SPLIT distance="500" swimtime="00:11:49.01" />
                    <SPLIT distance="550" swimtime="00:13:03.84" />
                    <SPLIT distance="600" swimtime="00:14:17.60" />
                    <SPLIT distance="650" swimtime="00:15:33.04" />
                    <SPLIT distance="700" swimtime="00:16:46.96" />
                    <SPLIT distance="750" swimtime="00:18:02.46" />
                    <SPLIT distance="800" swimtime="00:19:17.83" />
                    <SPLIT distance="850" swimtime="00:23:05.98" />
                    <SPLIT distance="900" swimtime="00:21:48.21" />
                    <SPLIT distance="1000" swimtime="00:24:22.54" />
                    <SPLIT distance="1050" swimtime="00:25:39.05" />
                    <SPLIT distance="1100" swimtime="00:26:55.70" />
                    <SPLIT distance="1150" swimtime="00:28:12.78" />
                    <SPLIT distance="1200" swimtime="00:29:29.47" />
                    <SPLIT distance="1250" swimtime="00:30:47.41" />
                    <SPLIT distance="1300" swimtime="00:32:02.58" />
                    <SPLIT distance="1350" swimtime="00:33:23.62" />
                    <SPLIT distance="1400" swimtime="00:34:40.35" />
                    <SPLIT distance="1450" swimtime="00:35:58.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="66" reactiontime="+105" swimtime="00:02:07.68" resultid="20709" heatid="24349" lane="9" entrytime="00:01:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="47" reactiontime="+120" swimtime="00:01:07.59" resultid="20710" heatid="24386" lane="2" entrytime="00:01:00.00" entrycourse="LCM" />
                <RESULT eventid="1491" points="76" reactiontime="+126" swimtime="00:04:25.75" resultid="20711" heatid="24410" lane="5" entrytime="00:04:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:04.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="102" reactiontime="+107" swimtime="00:01:02.82" resultid="20712" heatid="24455" lane="7" entrytime="00:01:00.00" entrycourse="LCM" />
                <RESULT eventid="1721" points="79" reactiontime="+114" swimtime="00:09:09.11" resultid="20713" heatid="24470" lane="1" entrytime="00:08:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.70" />
                    <SPLIT distance="100" swimtime="00:02:01.72" />
                    <SPLIT distance="150" swimtime="00:03:11.09" />
                    <SPLIT distance="200" swimtime="00:04:23.10" />
                    <SPLIT distance="250" swimtime="00:05:35.80" />
                    <SPLIT distance="300" swimtime="00:06:47.92" />
                    <SPLIT distance="350" swimtime="00:08:00.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1930-05-04" firstname="Stanisław" gender="M" lastname="Krokoszyński" nation="POL" athleteid="20698">
              <RESULTS>
                <RESULT eventid="1079" points="78" reactiontime="+127" swimtime="00:00:48.76" resultid="20699" heatid="24283" lane="3" entrytime="00:00:50.00" entrycourse="LCM" />
                <RESULT eventid="1113" points="47" reactiontime="+136" swimtime="00:05:13.73" resultid="20700" heatid="24301" lane="0" entrytime="00:05:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:04:10.52" />
                    <SPLIT distance="100" swimtime="00:02:44.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="57" swimtime="00:01:02.25" resultid="20701" heatid="24329" lane="9" entrytime="00:01:05.00" entrycourse="LCM" />
                <RESULT eventid="1273" points="71" reactiontime="+107" swimtime="00:01:53.18" resultid="20702" heatid="24355" lane="1" entrytime="00:01:58.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="53" reactiontime="+159" swimtime="00:02:31.12" resultid="20703" heatid="24381" lane="0" entrytime="00:02:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="65" reactiontime="+138" swimtime="00:04:12.74" resultid="20704" heatid="24416" lane="3" entrytime="00:03:58.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.81" />
                    <SPLIT distance="100" swimtime="00:02:01.00" />
                    <SPLIT distance="150" swimtime="00:03:06.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="51" swimtime="00:01:09.68" resultid="20705" heatid="24460" lane="8" entrytime="00:01:05.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-03-06" firstname="Ewa" gender="F" lastname="Rupp" nation="POL" athleteid="20714">
              <RESULTS>
                <RESULT eventid="1096" status="DNS" swimtime="00:00:00.00" resultid="20715" heatid="24297" lane="1" entrytime="00:04:36.40" entrycourse="LCM" />
                <RESULT eventid="1147" points="98" reactiontime="+123" swimtime="00:17:29.88" resultid="20716" heatid="24310" lane="6" entrytime="00:17:21.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:56.32" />
                    <SPLIT distance="250" swimtime="00:09:43.25" />
                    <SPLIT distance="300" swimtime="00:08:37.08" />
                    <SPLIT distance="350" swimtime="00:14:14.23" />
                    <SPLIT distance="400" swimtime="00:10:50.90" />
                    <SPLIT distance="450" swimtime="00:16:27.07" />
                    <SPLIT distance="500" swimtime="00:13:07.68" />
                    <SPLIT distance="600" swimtime="00:15:20.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="101" swimtime="00:00:58.00" resultid="20717" heatid="24324" lane="6" entrytime="00:00:56.16" entrycourse="LCM" />
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="20718" heatid="24349" lane="0" entrytime="00:01:48.10" entrycourse="LCM" />
                <RESULT eventid="1423" points="52" reactiontime="+87" swimtime="00:01:05.36" resultid="20719" heatid="24386" lane="7" entrytime="00:01:02.10" entrycourse="LCM" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="20720" heatid="24410" lane="3" entrytime="00:04:02.50" entrycourse="LCM" />
                <RESULT eventid="1595" points="47" reactiontime="+99" swimtime="00:02:33.63" resultid="20721" heatid="24434" lane="5" entrytime="00:02:19.00" entrycourse="LCM" />
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="20722" heatid="24470" lane="3" entrytime="00:08:20.10" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="20213" name="Masters Wrocław">
          <CONTACT name="Ostrasz" />
          <ATHLETES>
            <ATHLETE birthdate="1970-03-11" firstname="Anna" gender="F" lastname="Głowiak" nation="POL" athleteid="20214">
              <RESULTS>
                <RESULT eventid="1062" points="367" reactiontime="+87" swimtime="00:00:33.04" resultid="20215" heatid="24279" lane="1" entrytime="00:00:33.21" entrycourse="SCM" />
                <RESULT eventid="1147" points="313" reactiontime="+81" swimtime="00:11:53.57" resultid="20216" heatid="24312" lane="8" entrytime="00:11:54.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                    <SPLIT distance="100" swimtime="00:01:16.63" />
                    <SPLIT distance="150" swimtime="00:01:59.61" />
                    <SPLIT distance="200" swimtime="00:02:44.43" />
                    <SPLIT distance="250" swimtime="00:03:29.80" />
                    <SPLIT distance="300" swimtime="00:04:15.24" />
                    <SPLIT distance="350" swimtime="00:05:01.18" />
                    <SPLIT distance="400" swimtime="00:05:47.60" />
                    <SPLIT distance="450" swimtime="00:06:33.83" />
                    <SPLIT distance="500" swimtime="00:07:20.35" />
                    <SPLIT distance="550" swimtime="00:08:06.14" />
                    <SPLIT distance="600" swimtime="00:08:52.13" />
                    <SPLIT distance="650" swimtime="00:09:38.24" />
                    <SPLIT distance="750" swimtime="00:11:09.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="309" swimtime="00:00:40.01" resultid="20217" heatid="24325" lane="5" entrytime="00:00:41.01" entrycourse="SCM" />
                <RESULT eventid="1256" points="353" reactiontime="+62" swimtime="00:01:13.11" resultid="20218" heatid="24352" lane="9" entrytime="00:01:13.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="297" reactiontime="+98" swimtime="00:01:26.93" resultid="20219" heatid="24400" lane="4" entrytime="00:01:33.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="330" swimtime="00:02:43.35" resultid="20220" heatid="24413" lane="6" entrytime="00:02:39.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                    <SPLIT distance="100" swimtime="00:01:19.22" />
                    <SPLIT distance="150" swimtime="00:02:02.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="291" reactiontime="+92" swimtime="00:03:07.15" resultid="20221" heatid="24444" lane="1" entrytime="00:03:19.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.08" />
                    <SPLIT distance="100" swimtime="00:01:29.90" />
                    <SPLIT distance="150" swimtime="00:02:19.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="303" reactiontime="+79" swimtime="00:05:51.91" resultid="20222" heatid="24472" lane="3" entrytime="00:05:42.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.27" />
                    <SPLIT distance="100" swimtime="00:01:20.84" />
                    <SPLIT distance="150" swimtime="00:02:05.39" />
                    <SPLIT distance="200" swimtime="00:02:50.96" />
                    <SPLIT distance="250" swimtime="00:03:37.03" />
                    <SPLIT distance="300" swimtime="00:04:23.23" />
                    <SPLIT distance="350" swimtime="00:05:07.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-06-29" firstname="Piotr" gender="M" lastname="Krzekotowski" nation="POL" athleteid="20223">
              <RESULTS>
                <RESULT eventid="1079" points="161" reactiontime="+92" swimtime="00:00:38.39" resultid="20224" heatid="24285" lane="7" entrytime="00:00:37.90" entrycourse="SCM" />
                <RESULT eventid="1113" points="110" reactiontime="+105" swimtime="00:03:57.38" resultid="20225" heatid="24302" lane="1" entrytime="00:03:59.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.38" />
                    <SPLIT distance="100" swimtime="00:02:01.87" />
                    <SPLIT distance="150" swimtime="00:03:05.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="79" swimtime="00:00:55.71" resultid="20226" heatid="24329" lane="2" entrytime="00:00:59.00" entrycourse="SCM" />
                <RESULT eventid="1341" points="70" reactiontime="+93" swimtime="00:04:30.36" resultid="20227" heatid="24369" lane="7" entrytime="00:03:59.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.75" />
                    <SPLIT distance="100" swimtime="00:02:07.06" />
                    <SPLIT distance="150" swimtime="00:03:19.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="85" reactiontime="+91" swimtime="00:00:50.50" resultid="20228" heatid="24390" lane="3" entrytime="00:00:55.00" entrycourse="SCM" />
                <RESULT eventid="1578" points="100" reactiontime="+65" swimtime="00:08:43.92" resultid="20229" heatid="24431" lane="0" entrytime="00:08:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.16" />
                    <SPLIT distance="100" swimtime="00:02:11.21" />
                    <SPLIT distance="150" swimtime="00:03:27.35" />
                    <SPLIT distance="200" swimtime="00:04:43.54" />
                    <SPLIT distance="250" swimtime="00:05:47.78" />
                    <SPLIT distance="300" swimtime="00:06:53.71" />
                    <SPLIT distance="350" swimtime="00:07:49.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="66" swimtime="00:02:03.12" resultid="20230" heatid="24438" lane="9" entrytime="00:01:59.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="117" reactiontime="+63" swimtime="00:00:52.99" resultid="20231" heatid="24460" lane="6" entrytime="00:00:51.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-07-25" firstname="Piotr" gender="M" lastname="Ostrasz" nation="POL" athleteid="20232">
              <RESULTS>
                <RESULT eventid="1079" points="495" reactiontime="+75" swimtime="00:00:26.43" resultid="20233" heatid="24296" lane="0" entrytime="00:00:25.50" entrycourse="SCM" />
                <RESULT eventid="1273" points="481" reactiontime="+61" swimtime="00:00:59.86" resultid="20234" heatid="24363" lane="7" entrytime="00:00:59.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="442" swimtime="00:00:29.22" resultid="20235" heatid="24397" lane="8" entrytime="00:00:28.50" entrycourse="SCM" />
                <RESULT eventid="1681" points="428" swimtime="00:00:34.41" resultid="20236" heatid="24465" lane="6" entrytime="00:00:33.90" entrycourse="SCM" />
                <RESULT eventid="1744" points="279" swimtime="00:05:36.46" resultid="20237" heatid="24481" lane="7" entrytime="00:04:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                    <SPLIT distance="100" swimtime="00:01:11.70" />
                    <SPLIT distance="150" swimtime="00:01:51.56" />
                    <SPLIT distance="200" swimtime="00:02:33.52" />
                    <SPLIT distance="250" swimtime="00:03:17.71" />
                    <SPLIT distance="300" swimtime="00:04:03.68" />
                    <SPLIT distance="350" swimtime="00:04:50.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="21719" name="MASTERS Zdzieszowice">
          <CONTACT email="masters.zdzieszowice@gmail.com" name="Jajuga" phone="505127695" />
          <ATHLETES>
            <ATHLETE birthdate="1979-10-05" firstname="Ewelina" gender="F" lastname="Cuch" nation="POL" athleteid="21753">
              <RESULTS>
                <RESULT eventid="1222" points="250" reactiontime="+69" swimtime="00:03:40.70" resultid="21754" heatid="24339" lane="8" entrytime="00:03:42.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.39" />
                    <SPLIT distance="100" swimtime="00:01:46.15" />
                    <SPLIT distance="150" swimtime="00:02:41.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="257" swimtime="00:01:21.25" resultid="21755" heatid="24350" lane="5" entrytime="00:01:21.33" />
                <RESULT eventid="1388" points="253" reactiontime="+81" swimtime="00:01:41.32" resultid="21756" heatid="24378" lane="2" entrytime="00:01:39.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="255" swimtime="00:00:38.49" resultid="21757" heatid="24387" lane="5" entrytime="00:00:39.88" />
                <RESULT eventid="1595" status="DNS" swimtime="00:00:00.00" resultid="21758" heatid="24435" lane="3" entrytime="00:01:37.55" />
                <RESULT eventid="1664" points="265" reactiontime="+90" swimtime="00:00:45.76" resultid="21759" heatid="24456" lane="3" entrytime="00:00:45.36" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-11-02" firstname="Katarzyna" gender="F" lastname="Gniot" nation="POL" athleteid="21760">
              <RESULTS>
                <RESULT eventid="1062" status="DNS" swimtime="00:00:00.00" resultid="21761" heatid="24277" lane="6" entrytime="00:00:39.00" />
                <RESULT eventid="1096" status="DNS" swimtime="00:00:00.00" resultid="21762" heatid="24299" lane="9" entrytime="00:03:00.00" />
                <RESULT eventid="1388" status="DNS" swimtime="00:00:00.00" resultid="21763" heatid="24377" lane="6" entrytime="00:01:50.00" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="21764" heatid="24412" lane="0" entrytime="00:03:00.00" />
                <RESULT eventid="1630" status="DNS" swimtime="00:00:00.00" resultid="21765" heatid="24444" lane="9" entrytime="00:03:30.00" />
                <RESULT eventid="1664" status="DNS" swimtime="00:00:00.00" resultid="21766" heatid="24456" lane="8" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-15" firstname="Dawid" gender="M" lastname="Jajuga" nation="POL" athleteid="21720">
              <RESULTS>
                <RESULT eventid="1113" points="486" reactiontime="+84" swimtime="00:02:24.99" resultid="21721" heatid="24307" lane="0" entrytime="00:02:26.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.72" />
                    <SPLIT distance="100" swimtime="00:01:08.85" />
                    <SPLIT distance="150" swimtime="00:01:51.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14189" points="404" reactiontime="+81" swimtime="00:10:11.35" resultid="21722" heatid="24316" lane="6" entrytime="00:11:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                    <SPLIT distance="100" swimtime="00:01:11.25" />
                    <SPLIT distance="150" swimtime="00:01:49.60" />
                    <SPLIT distance="200" swimtime="00:02:28.12" />
                    <SPLIT distance="250" swimtime="00:03:06.49" />
                    <SPLIT distance="300" swimtime="00:03:45.06" />
                    <SPLIT distance="350" swimtime="00:04:23.46" />
                    <SPLIT distance="400" swimtime="00:05:01.98" />
                    <SPLIT distance="450" swimtime="00:05:39.85" />
                    <SPLIT distance="500" swimtime="00:06:18.78" />
                    <SPLIT distance="550" swimtime="00:06:58.40" />
                    <SPLIT distance="600" swimtime="00:07:38.00" />
                    <SPLIT distance="650" swimtime="00:08:17.76" />
                    <SPLIT distance="700" swimtime="00:08:57.10" />
                    <SPLIT distance="750" swimtime="00:09:35.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="447" swimtime="00:02:45.65" resultid="21723" heatid="24346" lane="8" entrytime="00:02:44.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                    <SPLIT distance="100" swimtime="00:01:21.12" />
                    <SPLIT distance="150" swimtime="00:02:03.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="422" reactiontime="+67" swimtime="00:02:28.61" resultid="21724" heatid="24371" lane="7" entrytime="00:02:25.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.81" />
                    <SPLIT distance="100" swimtime="00:01:08.63" />
                    <SPLIT distance="150" swimtime="00:01:47.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="440" swimtime="00:01:15.05" resultid="21725" heatid="24385" lane="9" entrytime="00:01:14.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="451" swimtime="00:05:17.77" resultid="21726" heatid="24433" lane="2" entrytime="00:05:10.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.82" />
                    <SPLIT distance="100" swimtime="00:01:08.35" />
                    <SPLIT distance="150" swimtime="00:01:51.70" />
                    <SPLIT distance="200" swimtime="00:02:35.11" />
                    <SPLIT distance="250" swimtime="00:03:19.75" />
                    <SPLIT distance="300" swimtime="00:04:05.77" />
                    <SPLIT distance="350" swimtime="00:04:42.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="471" swimtime="00:01:03.99" resultid="21727" heatid="24442" lane="8" entrytime="00:01:01.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="21728" heatid="24482" lane="9" entrytime="00:04:46.55" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-06" firstname="Fortunata" gender="F" lastname="Marczuk" nation="POL" athleteid="21737">
              <RESULTS>
                <RESULT eventid="1096" points="310" reactiontime="+95" swimtime="00:03:06.26" resultid="21738" heatid="24298" lane="4" entrytime="00:03:01.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.72" />
                    <SPLIT distance="100" swimtime="00:01:29.16" />
                    <SPLIT distance="150" swimtime="00:02:19.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" reactiontime="+99" status="OTL" swimtime="00:13:00.30" resultid="21739" heatid="24311" lane="2" entrytime="00:12:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.23" />
                    <SPLIT distance="100" swimtime="00:01:25.61" />
                    <SPLIT distance="150" swimtime="00:02:13.02" />
                    <SPLIT distance="200" swimtime="00:03:02.30" />
                    <SPLIT distance="300" swimtime="00:04:42.26" />
                    <SPLIT distance="350" swimtime="00:05:32.89" />
                    <SPLIT distance="400" swimtime="00:06:23.67" />
                    <SPLIT distance="450" swimtime="00:07:14.25" />
                    <SPLIT distance="500" swimtime="00:08:05.03" />
                    <SPLIT distance="600" swimtime="00:09:44.35" />
                    <SPLIT distance="700" swimtime="00:11:23.20" />
                    <SPLIT distance="750" swimtime="00:12:12.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="356" reactiontime="+72" swimtime="00:03:16.24" resultid="21740" heatid="24340" lane="2" entrytime="00:03:11.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.24" />
                    <SPLIT distance="100" swimtime="00:01:32.74" />
                    <SPLIT distance="150" swimtime="00:02:24.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="187" reactiontime="+81" swimtime="00:03:32.98" resultid="21741" heatid="24367" lane="2" entrytime="00:03:10.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.95" />
                    <SPLIT distance="100" swimtime="00:01:42.52" />
                    <SPLIT distance="150" swimtime="00:02:38.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="335" reactiontime="+59" swimtime="00:01:32.27" resultid="21742" heatid="24379" lane="0" entrytime="00:01:26.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="304" reactiontime="+73" swimtime="00:06:35.86" resultid="21743" heatid="24429" lane="6" entrytime="00:06:30.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.41" />
                    <SPLIT distance="100" swimtime="00:01:34.64" />
                    <SPLIT distance="150" swimtime="00:02:26.06" />
                    <SPLIT distance="200" swimtime="00:03:19.50" />
                    <SPLIT distance="250" swimtime="00:04:09.31" />
                    <SPLIT distance="300" swimtime="00:05:01.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="214" reactiontime="+58" swimtime="00:01:32.64" resultid="21744" heatid="24435" lane="5" entrytime="00:01:36.99" />
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="21745" heatid="24472" lane="2" entrytime="00:05:45.55" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-04-03" firstname="Daria" gender="F" lastname="Szydłowska - Smętek" nation="POL" athleteid="21746">
              <RESULTS>
                <RESULT eventid="1062" points="422" reactiontime="+96" swimtime="00:00:31.54" resultid="21747" heatid="24279" lane="4" entrytime="00:00:32.45" />
                <RESULT eventid="1147" points="384" reactiontime="+97" swimtime="00:11:06.89" resultid="21748" heatid="24311" lane="1" entrytime="00:13:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.00" />
                    <SPLIT distance="100" swimtime="00:01:17.66" />
                    <SPLIT distance="150" swimtime="00:03:25.58" />
                    <SPLIT distance="200" swimtime="00:02:42.39" />
                    <SPLIT distance="250" swimtime="00:04:51.18" />
                    <SPLIT distance="300" swimtime="00:04:08.29" />
                    <SPLIT distance="350" swimtime="00:06:16.26" />
                    <SPLIT distance="400" swimtime="00:05:33.97" />
                    <SPLIT distance="450" swimtime="00:07:41.38" />
                    <SPLIT distance="500" swimtime="00:06:58.83" />
                    <SPLIT distance="550" swimtime="00:09:05.63" />
                    <SPLIT distance="600" swimtime="00:09:47.65" />
                    <SPLIT distance="650" swimtime="00:10:27.88" />
                    <SPLIT distance="700" swimtime="00:11:06.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="351" swimtime="00:00:38.34" resultid="21749" heatid="24325" lane="2" entrytime="00:00:42.34" />
                <RESULT eventid="1256" points="402" reactiontime="+57" swimtime="00:01:10.04" resultid="21750" heatid="24352" lane="0" entrytime="00:01:12.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="399" reactiontime="+66" swimtime="00:02:33.43" resultid="21751" heatid="24413" lane="2" entrytime="00:02:40.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                    <SPLIT distance="100" swimtime="00:01:14.24" />
                    <SPLIT distance="150" swimtime="00:01:55.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="389" reactiontime="+59" swimtime="00:05:23.78" resultid="21752" heatid="24473" lane="9" entrytime="00:05:35.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                    <SPLIT distance="100" swimtime="00:01:17.35" />
                    <SPLIT distance="150" swimtime="00:01:58.74" />
                    <SPLIT distance="200" swimtime="00:02:40.17" />
                    <SPLIT distance="250" swimtime="00:03:21.62" />
                    <SPLIT distance="300" swimtime="00:04:02.80" />
                    <SPLIT distance="350" swimtime="00:04:43.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-09-15" firstname="Dorota" gender="F" lastname="Woźniak" nation="POL" athleteid="21729">
              <RESULTS>
                <RESULT eventid="1096" points="314" reactiontime="+100" swimtime="00:03:05.54" resultid="21730" heatid="24298" lane="6" entrytime="00:03:08.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                    <SPLIT distance="100" swimtime="00:01:28.60" />
                    <SPLIT distance="150" swimtime="00:02:21.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="319" swimtime="00:00:39.57" resultid="21731" heatid="24326" lane="7" entrytime="00:00:38.22" />
                <RESULT eventid="1324" points="232" reactiontime="+83" swimtime="00:03:18.12" resultid="21732" heatid="24367" lane="7" entrytime="00:03:17.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.28" />
                    <SPLIT distance="100" swimtime="00:01:34.97" />
                    <SPLIT distance="150" swimtime="00:02:27.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="300" reactiontime="+80" swimtime="00:01:26.57" resultid="21733" heatid="24401" lane="7" entrytime="00:01:27.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="277" reactiontime="+109" swimtime="00:06:48.22" resultid="21734" heatid="24429" lane="8" entrytime="00:07:15.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.47" />
                    <SPLIT distance="100" swimtime="00:01:34.21" />
                    <SPLIT distance="150" swimtime="00:02:27.62" />
                    <SPLIT distance="200" swimtime="00:03:19.78" />
                    <SPLIT distance="250" swimtime="00:04:18.01" />
                    <SPLIT distance="300" swimtime="00:05:15.84" />
                    <SPLIT distance="350" swimtime="00:06:03.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="294" reactiontime="+81" swimtime="00:03:06.46" resultid="21735" heatid="24444" lane="2" entrytime="00:03:11.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.25" />
                    <SPLIT distance="100" swimtime="00:01:30.67" />
                    <SPLIT distance="150" swimtime="00:02:19.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="242" reactiontime="+80" swimtime="00:06:19.25" resultid="21736" heatid="24471" lane="2" entrytime="00:06:30.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.36" />
                    <SPLIT distance="100" swimtime="00:01:29.79" />
                    <SPLIT distance="150" swimtime="00:02:18.05" />
                    <SPLIT distance="200" swimtime="00:03:06.19" />
                    <SPLIT distance="250" swimtime="00:03:55.00" />
                    <SPLIT distance="300" swimtime="00:04:43.61" />
                    <SPLIT distance="350" swimtime="00:05:32.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1358" points="325" reactiontime="+75" swimtime="00:02:34.61" resultid="21767" heatid="24372" lane="5" entrytime="00:02:20.11">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21729" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="21737" number="2" />
                    <RELAYPOSITION athleteid="21753" number="3" reactiontime="+12" />
                    <RELAYPOSITION athleteid="21746" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1525" points="341" reactiontime="+60" swimtime="00:02:17.98" resultid="21768" heatid="24425" lane="3" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                    <SPLIT distance="100" swimtime="00:01:08.00" />
                    <SPLIT distance="150" swimtime="00:01:42.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21746" number="1" reactiontime="+60" />
                    <RELAYPOSITION athleteid="21753" number="2" />
                    <RELAYPOSITION athleteid="21729" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="21737" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="21532" name="Masters Łódź">
          <CONTACT email="sport@masterslodz.pl" internet="http://masterslodz.pl" name="Trudnos Rafał" phone="604184311" />
          <ATHLETES>
            <ATHLETE birthdate="1977-06-06" firstname="Monika" gender="F" lastname="Klarecka" nation="POL" license="503605600029" athleteid="21533">
              <RESULTS>
                <RESULT eventid="1096" points="142" reactiontime="+114" swimtime="00:04:01.44" resultid="21534" heatid="24297" lane="6" entrytime="00:04:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.38" />
                    <SPLIT distance="150" swimtime="00:03:09.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="165" reactiontime="+123" swimtime="00:04:13.27" resultid="21535" heatid="24338" lane="6" entrytime="00:04:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.87" />
                    <SPLIT distance="150" swimtime="00:03:10.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="109" reactiontime="+75" swimtime="00:04:14.40" resultid="21536" heatid="24366" lane="5" entrytime="00:04:22.00" />
                <RESULT eventid="1423" points="110" reactiontime="+92" swimtime="00:00:50.98" resultid="21537" heatid="24386" lane="6" entrytime="00:00:57.00" />
                <RESULT eventid="1555" points="134" reactiontime="+91" swimtime="00:08:39.59" resultid="21538" heatid="24428" lane="5" entrytime="00:09:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:58.37" />
                    <SPLIT distance="200" swimtime="00:04:32.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MASKRAS" nation="POL" region="LBL" clubid="20451" name="Masterskrasnik">
          <CONTACT city="Kraśnik" email="masterskrasnik@gmail.pl" internet="masterdkrasnik.cba.pl" name="Michalczyk Jerzy" phone="601698977" state="LUB" street="Żwirki i Wigury 2" zip="23-210" />
          <ATHLETES>
            <ATHLETE birthdate="1956-01-09" firstname="Jerzy" gender="M" lastname="MIchalczyk" nation="POL" athleteid="20459">
              <RESULTS>
                <RESULT eventid="1079" points="106" reactiontime="+106" swimtime="00:00:44.17" resultid="20460" heatid="24283" lane="5" entrytime="00:00:48.00" />
                <RESULT eventid="1113" points="77" reactiontime="+102" swimtime="00:04:26.92" resultid="20461" heatid="24301" lane="3" entrytime="00:04:38.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.25" />
                    <SPLIT distance="100" swimtime="00:02:08.56" />
                    <SPLIT distance="150" swimtime="00:03:26.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="94" swimtime="00:00:52.67" resultid="20462" heatid="24329" lane="6" entrytime="00:00:58.40" />
                <RESULT eventid="1273" points="99" reactiontime="+64" swimtime="00:01:41.38" resultid="20463" heatid="24355" lane="7" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="82" reactiontime="+70" swimtime="00:00:51.09" resultid="20464" heatid="24390" lane="2" entrytime="00:00:57.20" />
                <RESULT eventid="1613" points="48" reactiontime="+71" swimtime="00:02:16.38" resultid="20465" heatid="24437" lane="5" entrytime="00:02:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-11-05" firstname="Krzysztof" gender="M" lastname="Samonek" nation="POL" athleteid="20452">
              <RESULTS>
                <RESULT eventid="1113" points="100" reactiontime="+122" swimtime="00:04:04.85" resultid="20453" heatid="24301" lane="5" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.81" />
                    <SPLIT distance="100" swimtime="00:01:58.42" />
                    <SPLIT distance="150" swimtime="00:03:10.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14189" reactiontime="+127" status="OTL" swimtime="00:16:15.47" resultid="20454" heatid="24314" lane="6" entrytime="00:15:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.82" />
                    <SPLIT distance="100" swimtime="00:01:50.61" />
                    <SPLIT distance="150" swimtime="00:02:51.35" />
                    <SPLIT distance="200" swimtime="00:03:52.90" />
                    <SPLIT distance="250" swimtime="00:04:55.84" />
                    <SPLIT distance="300" swimtime="00:05:58.29" />
                    <SPLIT distance="350" swimtime="00:07:01.27" />
                    <SPLIT distance="400" swimtime="00:08:03.60" />
                    <SPLIT distance="450" swimtime="00:09:06.31" />
                    <SPLIT distance="500" swimtime="00:10:07.59" />
                    <SPLIT distance="550" swimtime="00:11:10.21" />
                    <SPLIT distance="600" swimtime="00:12:11.79" />
                    <SPLIT distance="650" swimtime="00:13:14.22" />
                    <SPLIT distance="700" swimtime="00:14:16.90" />
                    <SPLIT distance="750" swimtime="00:15:17.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="115" swimtime="00:00:49.31" resultid="20455" heatid="24329" lane="5" entrytime="00:00:54.00" />
                <RESULT eventid="1474" points="96" reactiontime="+96" swimtime="00:01:53.11" resultid="20456" heatid="24404" lane="0" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="90" reactiontime="+93" swimtime="00:09:04.08" resultid="20457" heatid="24430" lane="4" entrytime="00:08:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.79" />
                    <SPLIT distance="100" swimtime="00:02:12.64" />
                    <SPLIT distance="150" swimtime="00:03:26.34" />
                    <SPLIT distance="200" swimtime="00:04:33.91" />
                    <SPLIT distance="250" swimtime="00:05:52.33" />
                    <SPLIT distance="300" swimtime="00:07:10.45" />
                    <SPLIT distance="350" swimtime="00:08:08.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="99" reactiontime="+90" swimtime="00:04:01.76" resultid="20458" heatid="24447" lane="5" entrytime="00:04:12.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:59.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="20392" name="MKP Szczecin">
          <CONTACT email="windmuhle@wp.pl" name="Kowalczyk Piotr" />
          <ATHLETES>
            <ATHLETE birthdate="1953-09-25" firstname="Sławomir" gender="M" lastname="Grzeszewski" nation="POL" athleteid="20420">
              <RESULTS>
                <RESULT eventid="1113" points="164" reactiontime="+95" swimtime="00:03:27.95" resultid="20421" heatid="24303" lane="9" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.46" />
                    <SPLIT distance="100" swimtime="00:01:41.26" />
                    <SPLIT distance="150" swimtime="00:02:39.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="183" reactiontime="+53" swimtime="00:03:42.72" resultid="20422" heatid="24343" lane="1" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.89" />
                    <SPLIT distance="100" swimtime="00:01:49.04" />
                    <SPLIT distance="150" swimtime="00:02:47.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="183" reactiontime="+44" swimtime="00:01:40.47" resultid="20423" heatid="24382" lane="0" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="20424" heatid="24392" lane="6" entrytime="00:00:37.00" />
                <RESULT eventid="1681" points="242" reactiontime="+42" swimtime="00:00:41.63" resultid="20425" heatid="24462" lane="2" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-02" firstname="Piotr" gender="M" lastname="Kowalczyk" nation="POL" athleteid="20413">
              <RESULTS>
                <RESULT eventid="14207" points="362" reactiontime="+92" swimtime="00:20:21.70" resultid="20414" heatid="24322" lane="1" entrytime="00:20:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                    <SPLIT distance="100" swimtime="00:01:14.03" />
                    <SPLIT distance="150" swimtime="00:01:53.05" />
                    <SPLIT distance="200" swimtime="00:02:32.91" />
                    <SPLIT distance="250" swimtime="00:03:12.59" />
                    <SPLIT distance="300" swimtime="00:03:52.49" />
                    <SPLIT distance="350" swimtime="00:04:32.89" />
                    <SPLIT distance="400" swimtime="00:05:13.31" />
                    <SPLIT distance="450" swimtime="00:05:53.66" />
                    <SPLIT distance="500" swimtime="00:06:34.18" />
                    <SPLIT distance="550" swimtime="00:07:15.74" />
                    <SPLIT distance="600" swimtime="00:07:57.27" />
                    <SPLIT distance="650" swimtime="00:08:38.77" />
                    <SPLIT distance="700" swimtime="00:09:19.98" />
                    <SPLIT distance="750" swimtime="00:10:01.34" />
                    <SPLIT distance="800" swimtime="00:10:42.51" />
                    <SPLIT distance="850" swimtime="00:11:23.60" />
                    <SPLIT distance="900" swimtime="00:12:04.67" />
                    <SPLIT distance="950" swimtime="00:12:46.05" />
                    <SPLIT distance="1000" swimtime="00:13:27.89" />
                    <SPLIT distance="1050" swimtime="00:14:09.88" />
                    <SPLIT distance="1100" swimtime="00:14:51.47" />
                    <SPLIT distance="1150" swimtime="00:15:33.40" />
                    <SPLIT distance="1200" swimtime="00:16:15.64" />
                    <SPLIT distance="1250" swimtime="00:16:57.29" />
                    <SPLIT distance="1300" swimtime="00:19:02.63" />
                    <SPLIT distance="1350" swimtime="00:18:21.01" />
                    <SPLIT distance="1450" swimtime="00:19:44.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="20415" heatid="24361" lane="2" entrytime="00:01:04.00" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="20416" heatid="24407" lane="9" entrytime="00:01:17.00" />
                <RESULT eventid="1508" points="381" reactiontime="+45" swimtime="00:02:20.64" resultid="20417" heatid="24422" lane="1" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.53" />
                    <SPLIT distance="100" swimtime="00:01:07.65" />
                    <SPLIT distance="150" swimtime="00:01:44.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="20418" heatid="24451" lane="9" entrytime="00:02:41.00" />
                <RESULT eventid="1744" points="381" reactiontime="+41" swimtime="00:05:03.41" resultid="20419" heatid="24481" lane="9" entrytime="00:05:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="100" swimtime="00:01:12.04" />
                    <SPLIT distance="150" swimtime="00:01:50.83" />
                    <SPLIT distance="200" swimtime="00:02:30.25" />
                    <SPLIT distance="250" swimtime="00:03:08.71" />
                    <SPLIT distance="300" swimtime="00:03:48.57" />
                    <SPLIT distance="350" swimtime="00:04:27.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1935-08-21" firstname="Stefania" gender="F" lastname="Noetzel" nation="POL" athleteid="20426">
              <RESULTS>
                <RESULT eventid="1187" points="28" swimtime="00:01:28.63" resultid="20427" heatid="24323" lane="3" entrytime="00:01:21.07" />
                <RESULT eventid="1222" points="59" swimtime="00:05:56.11" resultid="20428" heatid="24338" lane="0" entrytime="00:05:27.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:25.08" />
                    <SPLIT distance="100" swimtime="00:02:52.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="51" swimtime="00:02:52.29" resultid="20429" heatid="24376" lane="7" entrytime="00:02:33.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:22.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="57" swimtime="00:01:16.31" resultid="20430" heatid="24454" lane="4" entrytime="00:01:11.83" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-02-06" firstname="Lech" gender="M" lastname="Orecki" nation="POL" athleteid="20399">
              <RESULTS>
                <RESULT eventid="1079" points="280" reactiontime="+100" swimtime="00:00:31.95" resultid="20400" heatid="24289" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="14207" points="274" reactiontime="+101" swimtime="00:22:20.90" resultid="20401" heatid="24321" lane="5" entrytime="00:22:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.59" />
                    <SPLIT distance="100" swimtime="00:01:22.26" />
                    <SPLIT distance="150" swimtime="00:02:06.94" />
                    <SPLIT distance="200" swimtime="00:07:27.03" />
                    <SPLIT distance="250" swimtime="00:03:37.79" />
                    <SPLIT distance="300" swimtime="00:12:00.28" />
                    <SPLIT distance="350" swimtime="00:05:09.11" />
                    <SPLIT distance="400" swimtime="00:13:30.74" />
                    <SPLIT distance="450" swimtime="00:06:40.86" />
                    <SPLIT distance="500" swimtime="00:16:31.43" />
                    <SPLIT distance="550" swimtime="00:08:13.50" />
                    <SPLIT distance="650" swimtime="00:09:48.77" />
                    <SPLIT distance="750" swimtime="00:11:14.88" />
                    <SPLIT distance="850" swimtime="00:12:45.49" />
                    <SPLIT distance="950" swimtime="00:14:16.15" />
                    <SPLIT distance="1050" swimtime="00:15:45.73" />
                    <SPLIT distance="1150" swimtime="00:17:16.75" />
                    <SPLIT distance="1250" swimtime="00:18:46.93" />
                    <SPLIT distance="1350" swimtime="00:20:15.94" />
                    <SPLIT distance="1400" swimtime="00:20:59.56" />
                    <SPLIT distance="1450" swimtime="00:21:43.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="20402" heatid="24332" lane="7" entrytime="00:00:40.00" />
                <RESULT eventid="1273" points="297" swimtime="00:01:10.30" resultid="20403" heatid="24359" lane="6" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="20404" heatid="24405" lane="1" entrytime="00:01:30.00" />
                <RESULT eventid="1508" points="281" reactiontime="+41" swimtime="00:02:35.55" resultid="20405" heatid="24419" lane="5" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                    <SPLIT distance="100" swimtime="00:01:15.49" />
                    <SPLIT distance="150" swimtime="00:01:55.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="160" swimtime="00:03:26.02" resultid="20406" heatid="24449" lane="6" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.12" />
                    <SPLIT distance="100" swimtime="00:01:41.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="280" reactiontime="+48" swimtime="00:05:36.01" resultid="20407" heatid="24479" lane="0" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.49" />
                    <SPLIT distance="100" swimtime="00:01:21.49" />
                    <SPLIT distance="150" swimtime="00:02:05.01" />
                    <SPLIT distance="200" swimtime="00:02:50.00" />
                    <SPLIT distance="250" swimtime="00:03:33.89" />
                    <SPLIT distance="300" swimtime="00:04:17.19" />
                    <SPLIT distance="350" swimtime="00:04:58.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-06-07" firstname="Piotr" gender="M" lastname="Orłowski" nation="POL" athleteid="20431">
              <RESULTS>
                <RESULT eventid="1341" points="550" reactiontime="+82" swimtime="00:02:16.10" resultid="20432" heatid="24371" lane="3" entrytime="00:02:18.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.30" />
                    <SPLIT distance="100" swimtime="00:01:03.34" />
                    <SPLIT distance="150" swimtime="00:01:39.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="568" swimtime="00:00:26.89" resultid="20433" heatid="24398" lane="0" entrytime="00:00:26.76" />
                <RESULT eventid="1613" points="598" swimtime="00:00:59.13" resultid="20434" heatid="24442" lane="5" entrytime="00:00:59.58" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-08-10" firstname="Małgorzata" gender="F" lastname="Serbin" nation="POL" athleteid="20393">
              <RESULTS>
                <RESULT eventid="1165" points="388" reactiontime="+86" swimtime="00:21:01.35" resultid="20394" heatid="24319" lane="5" entrytime="00:20:20.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.30" />
                    <SPLIT distance="100" swimtime="00:01:16.71" />
                    <SPLIT distance="150" swimtime="00:01:57.57" />
                    <SPLIT distance="200" swimtime="00:02:38.77" />
                    <SPLIT distance="250" swimtime="00:03:20.00" />
                    <SPLIT distance="300" swimtime="00:04:01.56" />
                    <SPLIT distance="350" swimtime="00:04:43.37" />
                    <SPLIT distance="400" swimtime="00:05:25.05" />
                    <SPLIT distance="450" swimtime="00:06:07.00" />
                    <SPLIT distance="500" swimtime="00:06:49.14" />
                    <SPLIT distance="550" swimtime="00:07:31.14" />
                    <SPLIT distance="600" swimtime="00:08:13.51" />
                    <SPLIT distance="650" swimtime="00:08:55.69" />
                    <SPLIT distance="700" swimtime="00:09:38.02" />
                    <SPLIT distance="750" swimtime="00:10:20.20" />
                    <SPLIT distance="800" swimtime="00:11:02.43" />
                    <SPLIT distance="850" swimtime="00:11:45.10" />
                    <SPLIT distance="900" swimtime="00:12:27.71" />
                    <SPLIT distance="950" swimtime="00:13:10.36" />
                    <SPLIT distance="1000" swimtime="00:13:53.24" />
                    <SPLIT distance="1050" swimtime="00:14:36.92" />
                    <SPLIT distance="1100" swimtime="00:15:19.09" />
                    <SPLIT distance="1150" swimtime="00:16:02.04" />
                    <SPLIT distance="1200" swimtime="00:16:44.79" />
                    <SPLIT distance="1250" swimtime="00:17:27.91" />
                    <SPLIT distance="1300" swimtime="00:18:10.82" />
                    <SPLIT distance="1350" swimtime="00:18:53.59" />
                    <SPLIT distance="1400" swimtime="00:19:36.74" />
                    <SPLIT distance="1450" swimtime="00:20:19.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="405" reactiontime="+86" swimtime="00:01:09.86" resultid="20395" heatid="24352" lane="3" entrytime="00:01:09.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="405" swimtime="00:02:32.63" resultid="20396" heatid="24414" lane="9" entrytime="00:02:29.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.96" />
                    <SPLIT distance="100" swimtime="00:01:13.92" />
                    <SPLIT distance="150" swimtime="00:01:53.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="279" swimtime="00:03:09.77" resultid="20397" heatid="24445" lane="9" entrytime="00:03:04.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.56" />
                    <SPLIT distance="100" swimtime="00:01:32.73" />
                    <SPLIT distance="150" swimtime="00:02:21.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="416" swimtime="00:05:16.62" resultid="20398" heatid="24473" lane="0" entrytime="00:05:10.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                    <SPLIT distance="100" swimtime="00:01:16.58" />
                    <SPLIT distance="150" swimtime="00:01:56.55" />
                    <SPLIT distance="200" swimtime="00:02:36.90" />
                    <SPLIT distance="250" swimtime="00:03:17.07" />
                    <SPLIT distance="300" swimtime="00:03:57.67" />
                    <SPLIT distance="350" swimtime="00:04:37.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-10-02" firstname="Jadwiga" gender="F" lastname="Weber" nation="POL" athleteid="20408">
              <RESULTS>
                <RESULT eventid="1256" points="243" reactiontime="+85" swimtime="00:01:22.82" resultid="20409" heatid="24350" lane="3" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="258" reactiontime="+84" swimtime="00:01:31.02" resultid="20410" heatid="24401" lane="9" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="246" reactiontime="+87" swimtime="00:03:00.19" resultid="20411" heatid="24412" lane="1" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.03" />
                    <SPLIT distance="100" swimtime="00:01:26.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="258" swimtime="00:03:14.77" resultid="20412" heatid="24444" lane="6" entrytime="00:03:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.82" />
                    <SPLIT distance="100" swimtime="00:01:34.09" />
                    <SPLIT distance="150" swimtime="00:02:24.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="0811" nation="POL" region="SLA" clubid="21277" name="MKS Pałac Młodzieży Katowice">
          <CONTACT name="Jabczyk" phone="501341979" street="Mikołowska" />
          <ATHLETES>
            <ATHLETE birthdate="1997-08-04" firstname="Patrycja" gender="F" lastname="Bart" nation="POL" license="100811600172" athleteid="21287">
              <RESULTS>
                <RESULT eventid="1062" points="589" reactiontime="+79" swimtime="00:00:28.23" resultid="21288" heatid="24281" lane="5" entrytime="00:00:27.40" />
                <RESULT eventid="1096" points="598" reactiontime="+80" swimtime="00:02:29.66" resultid="21289" heatid="24299" lane="4" entrytime="00:02:30.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                    <SPLIT distance="100" swimtime="00:01:10.65" />
                    <SPLIT distance="150" swimtime="00:01:56.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="600" swimtime="00:00:32.07" resultid="21290" heatid="24327" lane="8" entrytime="00:00:35.44" />
                <RESULT eventid="1256" points="620" reactiontime="+79" swimtime="00:01:00.64" resultid="21291" heatid="24353" lane="4" entrytime="00:00:58.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="544" reactiontime="+71" swimtime="00:00:29.91" resultid="21292" heatid="24389" lane="3" entrytime="00:00:29.84" />
                <RESULT eventid="1491" points="642" reactiontime="+75" swimtime="00:02:10.96" resultid="21293" heatid="24414" lane="4" entrytime="00:02:07.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.61" />
                    <SPLIT distance="100" swimtime="00:01:03.68" />
                    <SPLIT distance="150" swimtime="00:01:37.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="532" reactiontime="+77" swimtime="00:01:08.43" resultid="21294" heatid="24436" lane="4" entrytime="00:01:06.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="466" reactiontime="+66" swimtime="00:00:37.91" resultid="21295" heatid="24454" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-05-15" firstname="Artur" gender="M" lastname="Pióro" nation="POL" license="100811700139" athleteid="21278">
              <RESULTS>
                <RESULT eventid="1113" points="563" reactiontime="+82" swimtime="00:02:18.03" resultid="21279" heatid="24307" lane="5" entrytime="00:02:15.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.37" />
                    <SPLIT distance="100" swimtime="00:01:04.24" />
                    <SPLIT distance="150" swimtime="00:01:46.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14189" points="615" reactiontime="+86" swimtime="00:08:51.62" resultid="21280" heatid="24317" lane="4" entrytime="00:08:30.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.11" />
                    <SPLIT distance="100" swimtime="00:01:02.22" />
                    <SPLIT distance="150" swimtime="00:01:34.75" />
                    <SPLIT distance="200" swimtime="00:02:07.48" />
                    <SPLIT distance="250" swimtime="00:02:40.33" />
                    <SPLIT distance="300" swimtime="00:03:13.56" />
                    <SPLIT distance="350" swimtime="00:03:46.82" />
                    <SPLIT distance="400" swimtime="00:04:20.31" />
                    <SPLIT distance="450" swimtime="00:04:54.11" />
                    <SPLIT distance="500" swimtime="00:05:28.28" />
                    <SPLIT distance="550" swimtime="00:06:01.61" />
                    <SPLIT distance="600" swimtime="00:06:36.00" />
                    <SPLIT distance="650" swimtime="00:07:09.89" />
                    <SPLIT distance="700" swimtime="00:07:44.08" />
                    <SPLIT distance="750" swimtime="00:08:18.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="515" reactiontime="+120" swimtime="00:00:29.93" resultid="21281" heatid="24335" lane="4" entrytime="00:00:29.06" />
                <RESULT eventid="1341" points="597" swimtime="00:02:12.40" resultid="21282" heatid="24371" lane="5" entrytime="00:02:17.43">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="517" reactiontime="+76" swimtime="00:00:27.73" resultid="21283" heatid="24397" lane="4" entrytime="00:00:27.29" />
                <RESULT eventid="1508" points="618" reactiontime="+74" swimtime="00:01:59.70" resultid="21284" heatid="24424" lane="4" entrytime="00:01:54.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.49" />
                    <SPLIT distance="100" swimtime="00:00:59.35" />
                    <SPLIT distance="150" swimtime="00:01:30.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="554" swimtime="00:01:00.63" resultid="21285" heatid="24442" lane="3" entrytime="00:00:59.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="654" reactiontime="+75" swimtime="00:04:13.52" resultid="21286" heatid="24482" lane="4" entrytime="00:04:03.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                    <SPLIT distance="100" swimtime="00:01:00.46" />
                    <SPLIT distance="150" swimtime="00:01:32.01" />
                    <SPLIT distance="200" swimtime="00:02:03.61" />
                    <SPLIT distance="250" swimtime="00:02:35.85" />
                    <SPLIT distance="300" swimtime="00:03:08.91" />
                    <SPLIT distance="350" swimtime="00:03:41.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SWDOL" nation="POL" region="DOL" clubid="20243" name="MKS Swim Academy Termy Jakuba Oława">
          <CONTACT city="Oława" email="biuro@swim-academy.pl" internet="www.swim-academy.pl" name="Grzegorz Fidala / Jacek Bereżnicki" phone="601316031 / 69643365" state="DOL" street="1 Maja 33a" zip="55-200" />
          <ATHLETES>
            <ATHLETE birthdate="1978-09-27" firstname="Magdalena" gender="F" lastname="Mruk" nation="POL" license="104501600044" athleteid="20244">
              <RESULTS>
                <RESULT eventid="1222" points="388" reactiontime="+77" swimtime="00:03:10.70" resultid="20245" heatid="24340" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.86" />
                    <SPLIT distance="100" swimtime="00:01:29.79" />
                    <SPLIT distance="150" swimtime="00:02:20.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="434" reactiontime="+77" swimtime="00:01:24.70" resultid="20246" heatid="24379" lane="1" entrytime="00:01:25.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="425" reactiontime="+73" swimtime="00:00:32.47" resultid="20247" heatid="24389" lane="0" entrytime="00:00:33.90" />
                <RESULT eventid="1595" points="336" reactiontime="+73" swimtime="00:01:19.78" resultid="20248" heatid="24436" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="450" reactiontime="+86" swimtime="00:00:38.35" resultid="20249" heatid="24458" lane="8" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="19927" name="MOSiR Ostrowiec Świętokrzyski">
          <CONTACT email="basen@mosir.ostrowiec.pl" name="Różalski Józef" phone="510-600-865" />
          <ATHLETES>
            <ATHLETE birthdate="1945-03-28" firstname="Józef" gender="M" lastname="Różalski" nation="POL" license="501012700001" athleteid="19928">
              <RESULTS>
                <RESULT eventid="1079" points="198" reactiontime="+99" swimtime="00:00:35.87" resultid="19929" heatid="24285" lane="2" entrytime="00:00:37.50" />
                <RESULT eventid="1113" points="123" reactiontime="+91" swimtime="00:03:48.87" resultid="19930" heatid="24302" lane="9" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.38" />
                    <SPLIT distance="100" swimtime="00:01:55.57" />
                    <SPLIT distance="150" swimtime="00:03:01.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="167" reactiontime="+86" swimtime="00:01:25.17" resultid="19931" heatid="24356" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="98" reactiontime="+53" swimtime="00:02:03.53" resultid="19932" heatid="24381" lane="5" entrytime="00:01:45.00" />
                <RESULT eventid="1440" points="185" reactiontime="+42" swimtime="00:00:39.04" resultid="19933" heatid="24391" lane="5" entrytime="00:00:40.50" />
                <RESULT eventid="1681" points="159" reactiontime="+41" swimtime="00:00:47.90" resultid="19934" heatid="24460" lane="5" entrytime="00:00:49.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOTYL" nation="POL" region="POM" clubid="20169" name="Motyl Mosir Stalowa Wola">
          <CONTACT city="Stalowa Wola" email="lorkowska@wp.pl" name="Chmielewski Andrzej" phone="600831914" street="Hutnicza 15" zip="37=450" />
          <ATHLETES>
            <ATHLETE birthdate="1973-01-14" firstname="Arkadiusz" gender="M" lastname="Berwecki" nation="POL" athleteid="20170">
              <RESULTS>
                <RESULT eventid="1079" points="471" reactiontime="+78" swimtime="00:00:26.86" resultid="20171" heatid="24294" lane="4" entrytime="00:00:26.49" />
                <RESULT eventid="1113" points="492" reactiontime="+75" swimtime="00:02:24.36" resultid="20172" heatid="24307" lane="6" entrytime="00:02:21.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.92" />
                    <SPLIT distance="100" swimtime="00:01:08.09" />
                    <SPLIT distance="150" swimtime="00:01:49.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="521" swimtime="00:00:58.27" resultid="20173" heatid="24365" lane="0" entrytime="00:00:56.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="480" swimtime="00:00:28.43" resultid="20174" heatid="24397" lane="2" entrytime="00:00:27.79" />
                <RESULT eventid="1508" points="512" reactiontime="+42" swimtime="00:02:07.44" resultid="20175" heatid="24424" lane="1" entrytime="00:02:06.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.44" />
                    <SPLIT distance="100" swimtime="00:01:02.97" />
                    <SPLIT distance="150" swimtime="00:01:35.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="523" swimtime="00:01:01.83" resultid="20176" heatid="24442" lane="7" entrytime="00:01:00.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="386" reactiontime="+85" swimtime="00:02:33.63" resultid="20177" heatid="24451" lane="3" entrytime="00:02:29.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                    <SPLIT distance="100" swimtime="00:01:14.13" />
                    <SPLIT distance="150" swimtime="00:01:54.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-02-27" firstname="Robert" gender="M" lastname="Lorkowski" nation="POL" athleteid="20178">
              <RESULTS>
                <RESULT eventid="1113" points="266" reactiontime="+96" swimtime="00:02:57.10" resultid="20179" heatid="24304" lane="0" entrytime="00:03:00.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                    <SPLIT distance="100" swimtime="00:01:24.78" />
                    <SPLIT distance="150" swimtime="00:02:17.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="176" reactiontime="+41" swimtime="00:03:18.79" resultid="20180" heatid="24370" lane="9" entrytime="00:03:27.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.00" />
                    <SPLIT distance="100" swimtime="00:01:32.73" />
                    <SPLIT distance="150" swimtime="00:02:26.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="262" reactiontime="+47" swimtime="00:02:39.34" resultid="20181" heatid="24419" lane="4" entrytime="00:02:38.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                    <SPLIT distance="100" swimtime="00:01:16.26" />
                    <SPLIT distance="150" swimtime="00:01:58.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="237" swimtime="00:06:33.54" resultid="20182" heatid="24432" lane="9" entrytime="00:06:34.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.26" />
                    <SPLIT distance="100" swimtime="00:01:33.32" />
                    <SPLIT distance="150" swimtime="00:02:22.94" />
                    <SPLIT distance="200" swimtime="00:03:12.70" />
                    <SPLIT distance="250" swimtime="00:04:09.68" />
                    <SPLIT distance="300" swimtime="00:05:05.93" />
                    <SPLIT distance="350" swimtime="00:05:51.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="227" reactiontime="+134" swimtime="00:03:03.42" resultid="20183" heatid="24449" lane="4" entrytime="00:03:02.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.43" />
                    <SPLIT distance="100" swimtime="00:01:29.55" />
                    <SPLIT distance="150" swimtime="00:02:17.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="20184" heatid="24478" lane="5" entrytime="00:05:54.03" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-07-07" firstname="Marcin" gender="M" lastname="Musialik" nation="POL" athleteid="20185">
              <RESULTS>
                <RESULT eventid="14207" points="438" reactiontime="+98" swimtime="00:19:06.80" resultid="20186" heatid="24322" lane="2" entrytime="00:19:15.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                    <SPLIT distance="100" swimtime="00:01:11.89" />
                    <SPLIT distance="150" swimtime="00:01:49.94" />
                    <SPLIT distance="200" swimtime="00:02:28.28" />
                    <SPLIT distance="250" swimtime="00:03:06.61" />
                    <SPLIT distance="300" swimtime="00:03:45.01" />
                    <SPLIT distance="350" swimtime="00:04:23.57" />
                    <SPLIT distance="400" swimtime="00:05:01.88" />
                    <SPLIT distance="450" swimtime="00:05:40.57" />
                    <SPLIT distance="500" swimtime="00:06:19.05" />
                    <SPLIT distance="550" swimtime="00:06:57.21" />
                    <SPLIT distance="600" swimtime="00:07:35.64" />
                    <SPLIT distance="650" swimtime="00:08:14.05" />
                    <SPLIT distance="700" swimtime="00:08:52.56" />
                    <SPLIT distance="750" swimtime="00:09:31.39" />
                    <SPLIT distance="800" swimtime="00:10:10.25" />
                    <SPLIT distance="850" swimtime="00:10:48.87" />
                    <SPLIT distance="900" swimtime="00:11:27.55" />
                    <SPLIT distance="950" swimtime="00:12:06.32" />
                    <SPLIT distance="1000" swimtime="00:12:45.07" />
                    <SPLIT distance="1050" swimtime="00:13:23.53" />
                    <SPLIT distance="1100" swimtime="00:14:02.11" />
                    <SPLIT distance="1150" swimtime="00:14:40.73" />
                    <SPLIT distance="1200" swimtime="00:15:19.59" />
                    <SPLIT distance="1250" swimtime="00:15:58.11" />
                    <SPLIT distance="1300" swimtime="00:16:36.77" />
                    <SPLIT distance="1350" swimtime="00:17:14.78" />
                    <SPLIT distance="1400" swimtime="00:17:52.84" />
                    <SPLIT distance="1450" swimtime="00:18:30.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="341" reactiontime="+89" swimtime="00:02:39.50" resultid="20187" heatid="24370" lane="4" entrytime="00:02:40.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                    <SPLIT distance="100" swimtime="00:01:16.02" />
                    <SPLIT distance="150" swimtime="00:01:57.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="453" swimtime="00:02:12.81" resultid="20188" heatid="24423" lane="9" entrytime="00:02:14.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.61" />
                    <SPLIT distance="100" swimtime="00:01:04.35" />
                    <SPLIT distance="150" swimtime="00:01:39.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="425" reactiontime="+41" swimtime="00:05:24.29" resultid="20189" heatid="24433" lane="1" entrytime="00:05:21.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                    <SPLIT distance="100" swimtime="00:01:12.03" />
                    <SPLIT distance="200" swimtime="00:02:35.60" />
                    <SPLIT distance="250" swimtime="00:03:23.36" />
                    <SPLIT distance="300" swimtime="00:04:10.95" />
                    <SPLIT distance="350" swimtime="00:04:48.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="403" reactiontime="+76" swimtime="00:02:31.46" resultid="20190" heatid="24451" lane="7" entrytime="00:02:34.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.07" />
                    <SPLIT distance="100" swimtime="00:01:14.38" />
                    <SPLIT distance="150" swimtime="00:01:53.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="455" swimtime="00:04:45.95" resultid="20191" heatid="24482" lane="0" entrytime="00:04:45.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                    <SPLIT distance="100" swimtime="00:01:07.82" />
                    <SPLIT distance="150" swimtime="00:01:43.19" />
                    <SPLIT distance="200" swimtime="00:02:19.49" />
                    <SPLIT distance="250" swimtime="00:02:55.43" />
                    <SPLIT distance="300" swimtime="00:03:32.88" />
                    <SPLIT distance="350" swimtime="00:04:09.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-26" firstname="Krzysztof" gender="M" lastname="Pawłowski" nation="POL" athleteid="20192">
              <RESULTS>
                <RESULT eventid="1079" points="352" reactiontime="+80" swimtime="00:00:29.61" resultid="20193" heatid="24289" lane="5" entrytime="00:00:30.27" />
                <RESULT eventid="14189" points="265" reactiontime="+87" swimtime="00:11:43.35" resultid="20194" heatid="24316" lane="2" entrytime="00:11:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                    <SPLIT distance="100" swimtime="00:01:17.71" />
                    <SPLIT distance="150" swimtime="00:02:01.77" />
                    <SPLIT distance="200" swimtime="00:02:46.65" />
                    <SPLIT distance="250" swimtime="00:03:31.78" />
                    <SPLIT distance="300" swimtime="00:04:16.87" />
                    <SPLIT distance="350" swimtime="00:05:02.10" />
                    <SPLIT distance="400" swimtime="00:05:47.22" />
                    <SPLIT distance="450" swimtime="00:06:32.22" />
                    <SPLIT distance="500" swimtime="00:07:17.41" />
                    <SPLIT distance="550" swimtime="00:08:02.83" />
                    <SPLIT distance="600" swimtime="00:08:48.14" />
                    <SPLIT distance="650" swimtime="00:09:32.81" />
                    <SPLIT distance="700" swimtime="00:10:17.26" />
                    <SPLIT distance="750" swimtime="00:11:01.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="342" swimtime="00:00:34.29" resultid="20195" heatid="24330" lane="9" entrytime="00:00:52.20" />
                <RESULT eventid="1239" points="313" swimtime="00:03:06.52" resultid="20196" heatid="24344" lane="2" entrytime="00:03:10.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.03" />
                    <SPLIT distance="100" swimtime="00:01:28.42" />
                    <SPLIT distance="150" swimtime="00:02:18.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="300" swimtime="00:01:25.28" resultid="20197" heatid="24383" lane="6" entrytime="00:01:25.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="320" reactiontime="+98" swimtime="00:01:15.78" resultid="20198" heatid="24407" lane="0" entrytime="00:01:16.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="320" reactiontime="+88" swimtime="00:02:43.55" resultid="20199" heatid="24449" lane="2" entrytime="00:03:10.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.56" />
                    <SPLIT distance="100" swimtime="00:01:18.75" />
                    <SPLIT distance="150" swimtime="00:02:01.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="365" reactiontime="+66" swimtime="00:00:36.30" resultid="20200" heatid="24464" lane="7" entrytime="00:00:36.32" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-04-17" firstname="Maria" gender="F" lastname="Petecka" nation="POL" athleteid="20201">
              <RESULTS>
                <RESULT eventid="1062" points="276" reactiontime="+97" swimtime="00:00:36.33" resultid="20202" heatid="24278" lane="2" entrytime="00:00:36.01" />
                <RESULT eventid="1096" points="257" reactiontime="+92" swimtime="00:03:18.35" resultid="20203" heatid="24298" lane="8" entrytime="00:03:16.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.41" />
                    <SPLIT distance="100" swimtime="00:01:38.43" />
                    <SPLIT distance="150" swimtime="00:02:33.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="235" reactiontime="+77" swimtime="00:03:45.14" resultid="20204" heatid="24339" lane="7" entrytime="00:03:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.90" />
                    <SPLIT distance="100" swimtime="00:01:50.69" />
                    <SPLIT distance="150" swimtime="00:02:48.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="218" reactiontime="+79" swimtime="00:01:46.51" resultid="20205" heatid="24378" lane="8" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="183" reactiontime="+78" swimtime="00:00:43.02" resultid="20206" heatid="24387" lane="6" entrytime="00:00:41.00" />
                <RESULT eventid="1595" points="173" reactiontime="+88" swimtime="00:01:39.50" resultid="20207" heatid="24435" lane="4" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="219" reactiontime="+79" swimtime="00:00:48.75" resultid="20208" heatid="24456" lane="2" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="19766" name="Nabaiji Team Decathlon">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1986-11-21" firstname="Laura" gender="F" lastname="Abucewicz" nation="POL" athleteid="21908">
              <RESULTS>
                <RESULT eventid="1062" points="122" reactiontime="+76" swimtime="00:00:47.68" resultid="21909" heatid="24276" lane="9" />
                <RESULT eventid="1187" points="125" swimtime="00:00:54.03" resultid="21910" heatid="24325" lane="1" entrytime="00:00:45.00" />
                <RESULT eventid="1664" points="106" reactiontime="+69" swimtime="00:01:02.04" resultid="21911" heatid="24453" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-06" firstname="Paweł" gender="M" lastname="Bednarczyk" nation="POL" athleteid="21928">
              <RESULTS>
                <RESULT eventid="1113" points="406" reactiontime="+77" swimtime="00:02:33.89" resultid="21929" heatid="24307" lane="7" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.31" />
                    <SPLIT distance="100" swimtime="00:01:10.18" />
                    <SPLIT distance="150" swimtime="00:01:54.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14189" reactiontime="+91" status="OTL" swimtime="00:11:17.16" resultid="21930" heatid="24317" lane="0" entrytime="00:10:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.28" />
                    <SPLIT distance="100" swimtime="00:01:12.16" />
                    <SPLIT distance="150" swimtime="00:01:50.51" />
                    <SPLIT distance="200" swimtime="00:02:31.37" />
                    <SPLIT distance="250" swimtime="00:03:12.62" />
                    <SPLIT distance="300" swimtime="00:03:55.74" />
                    <SPLIT distance="350" swimtime="00:04:38.87" />
                    <SPLIT distance="400" swimtime="00:05:22.94" />
                    <SPLIT distance="450" swimtime="00:06:07.02" />
                    <SPLIT distance="500" swimtime="00:06:51.88" />
                    <SPLIT distance="550" swimtime="00:07:36.06" />
                    <SPLIT distance="600" swimtime="00:08:19.91" />
                    <SPLIT distance="650" swimtime="00:09:03.90" />
                    <SPLIT distance="700" swimtime="00:09:48.51" />
                    <SPLIT distance="750" swimtime="00:10:33.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="532" swimtime="00:00:57.87" resultid="21931" heatid="24365" lane="6" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="561" swimtime="00:00:27.00" resultid="21932" heatid="24398" lane="6" entrytime="00:00:26.00" />
                <RESULT eventid="1578" points="344" swimtime="00:05:47.90" resultid="21933" heatid="24433" lane="0" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.26" />
                    <SPLIT distance="100" swimtime="00:01:08.40" />
                    <SPLIT distance="150" swimtime="00:01:54.87" />
                    <SPLIT distance="200" swimtime="00:02:41.47" />
                    <SPLIT distance="250" swimtime="00:03:30.73" />
                    <SPLIT distance="300" swimtime="00:04:22.09" />
                    <SPLIT distance="350" swimtime="00:05:05.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="21934" heatid="24442" lane="2" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-03-31" firstname="Agnieszka" gender="F" lastname="Dusza-Sabadasz" nation="POL" athleteid="21894">
              <RESULTS>
                <RESULT eventid="1062" points="230" reactiontime="+83" swimtime="00:00:38.58" resultid="21895" heatid="24278" lane="9" entrytime="00:00:37.55" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-04-06" firstname="Martyna" gender="F" lastname="Górajewska" nation="POL" athleteid="21899">
              <RESULTS>
                <RESULT eventid="1062" points="375" reactiontime="+94" swimtime="00:00:32.82" resultid="21900" heatid="24280" lane="0" entrytime="00:00:32.00" />
                <RESULT eventid="1664" points="331" reactiontime="+82" swimtime="00:00:42.49" resultid="21901" heatid="24457" lane="4" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-05-17" firstname="Zuzanna" gender="F" lastname="Kacalska" nation="POL" athleteid="21935">
              <RESULTS>
                <RESULT eventid="1062" points="430" reactiontime="+88" swimtime="00:00:31.34" resultid="21936" heatid="24280" lane="2" entrytime="00:00:30.80" />
                <RESULT eventid="1256" points="392" reactiontime="+81" swimtime="00:01:10.61" resultid="21937" heatid="24352" lane="8" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="388" reactiontime="+77" swimtime="00:02:34.81" resultid="21938" heatid="24413" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.83" />
                    <SPLIT distance="100" swimtime="00:01:14.44" />
                    <SPLIT distance="150" swimtime="00:01:55.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-08-27" firstname="Aneta" gender="F" lastname="Konkel" nation="POL" athleteid="21902">
              <RESULTS>
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="21903" heatid="24347" lane="4" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="21904" heatid="24409" lane="5" />
                <RESULT eventid="1222" points="124" reactiontime="+89" swimtime="00:04:38.44" resultid="24067" heatid="24337" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:13.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-10-02" firstname="Agnieszka" gender="F" lastname="Kos" nation="POL" athleteid="21951">
              <RESULTS>
                <RESULT eventid="1062" points="231" reactiontime="+87" swimtime="00:00:38.57" resultid="21952" heatid="24277" lane="2" entrytime="00:00:39.00" />
                <RESULT eventid="1256" points="180" reactiontime="+65" swimtime="00:01:31.43" resultid="21953" heatid="24349" lane="7" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-11-23" firstname="Filip" gender="M" lastname="Kołodziejski" nation="POL" athleteid="21954">
              <RESULTS>
                <RESULT eventid="1205" points="702" reactiontime="+67" swimtime="00:00:27.00" resultid="21955" heatid="24336" lane="5" entrytime="00:00:27.15" />
                <RESULT eventid="1474" points="675" reactiontime="+118" swimtime="00:00:59.10" resultid="21956" heatid="24408" lane="4" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="578" reactiontime="+112" swimtime="00:02:14.34" resultid="21957" heatid="24452" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.97" />
                    <SPLIT distance="100" swimtime="00:01:05.99" />
                    <SPLIT distance="150" swimtime="00:01:41.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-04-25" firstname="Mateusz" gender="M" lastname="Kołodziejski" nation="POL" athleteid="22618">
              <RESULTS>
                <RESULT eventid="1406" points="641" swimtime="00:01:06.20" resultid="22619" heatid="24385" lane="4" entrytime="00:01:05.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="592" swimtime="00:00:26.52" resultid="22620" heatid="24398" lane="5" entrytime="00:00:25.95" />
                <RESULT eventid="1681" points="670" swimtime="00:00:29.65" resultid="22621" heatid="24466" lane="6" entrytime="00:00:29.24" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-04-15" firstname="Rafał" gender="M" lastname="Krupiński" nation="POL" athleteid="21912">
              <RESULTS>
                <RESULT eventid="1273" points="155" reactiontime="+43" swimtime="00:01:27.29" resultid="21913" heatid="24354" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="124" reactiontime="+70" swimtime="00:03:24.19" resultid="21914" heatid="24416" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.26" />
                    <SPLIT distance="100" swimtime="00:01:35.38" />
                    <SPLIT distance="150" swimtime="00:02:31.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-04-02" firstname="Karolina" gender="F" lastname="Mazurek-Świstak" nation="POL" athleteid="21924">
              <RESULTS>
                <RESULT eventid="1187" points="508" swimtime="00:00:33.90" resultid="21925" heatid="24327" lane="9" entrytime="00:00:36.00" />
                <RESULT eventid="1388" points="446" reactiontime="+47" swimtime="00:01:23.89" resultid="21926" heatid="24379" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="493" swimtime="00:00:37.21" resultid="21927" heatid="24458" lane="1" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-04-07" firstname="Marzena" gender="F" lastname="Mikołajek" nation="POL" athleteid="21896">
              <RESULTS>
                <RESULT eventid="1256" points="279" reactiontime="+77" swimtime="00:01:19.10" resultid="21897" heatid="24351" lane="9" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="199" reactiontime="+99" swimtime="00:03:13.42" resultid="21898" heatid="24409" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.92" />
                    <SPLIT distance="100" swimtime="00:01:32.16" />
                    <SPLIT distance="150" swimtime="00:02:23.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-26" firstname="Bartosz" gender="M" lastname="Miller" nation="POL" athleteid="21915">
              <RESULTS>
                <RESULT eventid="1273" points="148" reactiontime="+58" swimtime="00:01:28.67" resultid="21916" heatid="24354" lane="5" />
                <RESULT eventid="1508" points="123" reactiontime="+90" swimtime="00:03:24.89" resultid="21917" heatid="24415" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.91" />
                    <SPLIT distance="100" swimtime="00:01:35.26" />
                    <SPLIT distance="150" swimtime="00:02:29.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-20" firstname="Kamila" gender="F" lastname="Popielarz" nation="POL" athleteid="21905">
              <RESULTS>
                <RESULT eventid="1062" points="101" reactiontime="+119" swimtime="00:00:50.71" resultid="21906" heatid="24276" lane="1" />
                <RESULT eventid="1256" points="73" reactiontime="+60" swimtime="00:02:03.32" resultid="21907" heatid="24348" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-11-04" firstname="Tomasz" gender="M" lastname="Sabadasz" nation="POL" athleteid="19767">
              <RESULTS>
                <RESULT eventid="1113" points="205" reactiontime="+84" swimtime="00:03:13.30" resultid="19768" heatid="24303" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.46" />
                    <SPLIT distance="100" swimtime="00:01:36.14" />
                    <SPLIT distance="150" swimtime="00:02:29.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="195" swimtime="00:07:00.35" resultid="19769" heatid="24431" lane="5" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.97" />
                    <SPLIT distance="100" swimtime="00:01:40.20" />
                    <SPLIT distance="200" swimtime="00:03:33.70" />
                    <SPLIT distance="250" swimtime="00:04:30.61" />
                    <SPLIT distance="300" swimtime="00:05:29.11" />
                    <SPLIT distance="350" swimtime="00:06:16.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-18" firstname="Emil" gender="M" lastname="Strumiński" nation="POL" athleteid="21918">
              <RESULTS>
                <RESULT eventid="1079" points="519" reactiontime="+73" swimtime="00:00:26.01" resultid="21919" heatid="24294" lane="6" entrytime="00:00:26.50" />
                <RESULT eventid="1273" points="564" swimtime="00:00:56.75" resultid="21920" heatid="24363" lane="5" entrytime="00:00:58.50" />
                <RESULT eventid="1440" points="523" reactiontime="+66" swimtime="00:00:27.64" resultid="21921" heatid="24396" lane="3" entrytime="00:00:28.80" />
                <RESULT eventid="1508" points="454" swimtime="00:02:12.70" resultid="21922" heatid="24423" lane="0" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.92" />
                    <SPLIT distance="100" swimtime="00:01:03.65" />
                    <SPLIT distance="150" swimtime="00:01:38.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="491" swimtime="00:01:03.15" resultid="21923" heatid="24441" lane="2" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-09-04" firstname="Mateusz" gender="M" lastname="Turowski" nation="POL" athleteid="21947">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="21948" heatid="24293" lane="4" entrytime="00:00:27.00" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="21949" heatid="24364" lane="8" entrytime="00:00:58.00" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="21950" heatid="24396" lane="9" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-01" firstname="Piotr" gender="M" lastname="Ławniczak" nation="POL" athleteid="21943">
              <RESULTS>
                <RESULT eventid="1079" points="378" reactiontime="+71" swimtime="00:00:28.90" resultid="21944" heatid="24294" lane="9" entrytime="00:00:27.00" />
                <RESULT eventid="1273" points="380" swimtime="00:01:04.76" resultid="21945" heatid="24364" lane="7" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="21946" heatid="24395" lane="4" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-03-18" firstname="Krystian" gender="M" lastname="Łukaszewicz" nation="POL" athleteid="21939">
              <RESULTS>
                <RESULT eventid="1079" points="446" reactiontime="+90" swimtime="00:00:27.35" resultid="21940" heatid="24293" lane="5" entrytime="00:00:27.00" />
                <RESULT eventid="1273" points="427" reactiontime="+88" swimtime="00:01:02.25" resultid="21941" heatid="24364" lane="2" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="21942" heatid="24398" lane="7" entrytime="00:00:26.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="366" reactiontime="+62" swimtime="00:02:10.54" resultid="21964" heatid="24373" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                    <SPLIT distance="100" swimtime="00:01:09.80" />
                    <SPLIT distance="150" swimtime="00:01:41.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21947" number="1" reactiontime="+62" />
                    <RELAYPOSITION athleteid="21928" number="2" />
                    <RELAYPOSITION athleteid="21918" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="21939" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1548" points="361" reactiontime="+80" swimtime="00:01:59.13" resultid="21966" heatid="24426" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.71" />
                    <SPLIT distance="100" swimtime="00:01:00.61" />
                    <SPLIT distance="150" swimtime="00:01:35.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21928" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="21918" number="2" />
                    <RELAYPOSITION athleteid="21912" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="22618" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" status="DNS" swimtime="00:00:00.00" resultid="21967" heatid="24426" lane="2">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21954" number="1" />
                    <RELAYPOSITION athleteid="21915" number="2" />
                    <RELAYPOSITION athleteid="21943" number="3" />
                    <RELAYPOSITION athleteid="21912" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1358" points="392" reactiontime="+79" swimtime="00:02:25.22" resultid="21961" heatid="24372" lane="3" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.12" />
                    <SPLIT distance="100" swimtime="00:01:15.93" />
                    <SPLIT distance="150" swimtime="00:01:52.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21924" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="21899" number="2" />
                    <RELAYPOSITION athleteid="21935" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="21896" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1525" points="440" reactiontime="+77" swimtime="00:02:06.77" resultid="21962" heatid="24425" lane="4" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                    <SPLIT distance="100" swimtime="00:01:03.62" />
                    <SPLIT distance="150" swimtime="00:01:35.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21924" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="21896" number="2" />
                    <RELAYPOSITION athleteid="21899" number="3" reactiontime="+12" />
                    <RELAYPOSITION athleteid="21935" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1525" points="111" swimtime="00:03:20.38" resultid="21963" heatid="24425" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.89" />
                    <SPLIT distance="100" swimtime="00:01:49.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21908" number="1" />
                    <RELAYPOSITION athleteid="21902" number="2" />
                    <RELAYPOSITION athleteid="21951" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="21905" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" reactiontime="+84" swimtime="00:02:08.16" resultid="21958" heatid="24309" lane="9" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                    <SPLIT distance="100" swimtime="00:01:11.62" />
                    <SPLIT distance="150" swimtime="00:01:39.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21899" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="21894" number="2" />
                    <RELAYPOSITION athleteid="21939" number="3" reactiontime="+79" />
                    <RELAYPOSITION athleteid="21943" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1130" status="DNS" swimtime="00:00:00.00" resultid="21959" heatid="24309" lane="4" entrytime="00:01:51.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21947" number="1" />
                    <RELAYPOSITION athleteid="21924" number="2" />
                    <RELAYPOSITION athleteid="21928" number="3" />
                    <RELAYPOSITION athleteid="21935" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" status="DNS" swimtime="00:00:00.00" resultid="21960" heatid="24467" lane="6">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21947" number="1" />
                    <RELAYPOSITION athleteid="21924" number="2" />
                    <RELAYPOSITION athleteid="21928" number="3" />
                    <RELAYPOSITION athleteid="21935" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="19755" name="Niezrzeszeni">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1965-07-28" firstname="Dorota" gender="F" lastname="Bernat" nation="POL" athleteid="23080">
              <RESULTS>
                <RESULT eventid="1222" points="97" reactiontime="+113" swimtime="00:05:02.38" resultid="23081" heatid="24338" lane="7" entrytime="00:05:02.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.83" />
                    <SPLIT distance="100" swimtime="00:02:25.81" />
                    <SPLIT distance="150" swimtime="00:03:45.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="46" reactiontime="+99" swimtime="00:02:23.79" resultid="23082" heatid="24348" lane="2" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="94" reactiontime="+79" swimtime="00:02:20.78" resultid="23083" heatid="24377" lane="9" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="43" reactiontime="+97" swimtime="00:05:20.07" resultid="23084" heatid="24410" lane="8" entrytime="00:05:06.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.84" />
                    <SPLIT distance="100" swimtime="00:02:38.37" />
                    <SPLIT distance="150" swimtime="00:04:03.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="91" reactiontime="+91" swimtime="00:01:05.18" resultid="23085" heatid="24455" lane="8" entrytime="00:01:02.70" />
                <RESULT eventid="1721" points="45" reactiontime="+94" swimtime="00:11:03.70" resultid="23086" heatid="24469" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.96" />
                    <SPLIT distance="100" swimtime="00:02:35.80" />
                    <SPLIT distance="150" swimtime="00:03:59.87" />
                    <SPLIT distance="200" swimtime="00:05:26.84" />
                    <SPLIT distance="250" swimtime="00:06:53.47" />
                    <SPLIT distance="300" swimtime="00:08:20.10" />
                    <SPLIT distance="350" swimtime="00:09:46.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-22" firstname="Piotr" gender="M" lastname="Burzyński" nation="POL" athleteid="19800">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="19801" heatid="24286" lane="4" entrytime="00:00:34.62" />
                <RESULT eventid="14207" status="DNS" swimtime="00:00:00.00" resultid="19802" heatid="24321" lane="9" entrytime="00:26:15.00" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="19803" heatid="24342" lane="5" entrytime="00:03:51.00" />
                <RESULT eventid="1341" status="DNS" swimtime="00:00:00.00" resultid="19804" heatid="24369" lane="8" entrytime="00:04:10.20" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="19805" heatid="24418" lane="9" entrytime="00:03:10.20" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="19806" heatid="24431" lane="1" entrytime="00:07:48.00" />
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="19807" heatid="24448" lane="0" entrytime="00:03:50.00" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="19808" heatid="24477" lane="5" entrytime="00:06:23.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-05-20" firstname="Ewa" gender="F" lastname="Cygan" nation="POL" athleteid="23853">
              <RESULTS>
                <RESULT eventid="1388" points="36" reactiontime="+149" swimtime="00:03:13.82" resultid="23854" heatid="24376" lane="5" entrytime="00:02:15.41" />
                <RESULT eventid="1256" points="20" reactiontime="+137" swimtime="00:03:09.33" resultid="23855" heatid="24347" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:25.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="25" swimtime="00:01:32.04" resultid="23856" heatid="24323" lane="7" />
                <RESULT eventid="1664" points="47" reactiontime="+129" swimtime="00:01:21.31" resultid="23857" heatid="24453" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="Bolesław" gender="M" lastname="Czyż" nation="POL" athleteid="22672">
              <RESULTS>
                <RESULT eventid="1341" points="56" reactiontime="+83" swimtime="00:04:51.43" resultid="22673" heatid="24368" lane="5" entrytime="00:04:46.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:19.25" />
                    <SPLIT distance="150" swimtime="00:03:37.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="87" reactiontime="+83" swimtime="00:09:08.97" resultid="22674" heatid="24430" lane="6" entrytime="00:09:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.19" />
                    <SPLIT distance="100" swimtime="00:02:16.94" />
                    <SPLIT distance="150" swimtime="00:03:27.66" />
                    <SPLIT distance="200" swimtime="00:04:35.11" />
                    <SPLIT distance="250" swimtime="00:05:50.57" />
                    <SPLIT distance="300" swimtime="00:07:03.61" />
                    <SPLIT distance="350" swimtime="00:08:07.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1941-11-21" firstname="Zbigniew" gender="M" lastname="Dymecki" nation="POL" athleteid="19935">
              <RESULTS>
                <RESULT eventid="1113" points="72" reactiontime="+135" swimtime="00:04:33.03" resultid="19936" heatid="24301" lane="2" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.95" />
                    <SPLIT distance="100" swimtime="00:02:19.46" />
                    <SPLIT distance="150" swimtime="00:03:33.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14189" points="72" reactiontime="+122" swimtime="00:18:04.97" resultid="19937" heatid="24313" lane="4" entrytime="00:18:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.34" />
                    <SPLIT distance="100" swimtime="00:02:05.86" />
                    <SPLIT distance="150" swimtime="00:03:13.09" />
                    <SPLIT distance="200" swimtime="00:04:23.88" />
                    <SPLIT distance="250" swimtime="00:05:31.47" />
                    <SPLIT distance="300" swimtime="00:06:41.01" />
                    <SPLIT distance="350" swimtime="00:07:50.05" />
                    <SPLIT distance="400" swimtime="00:08:59.38" />
                    <SPLIT distance="450" swimtime="00:10:09.59" />
                    <SPLIT distance="500" swimtime="00:11:17.82" />
                    <SPLIT distance="550" swimtime="00:12:27.72" />
                    <SPLIT distance="600" swimtime="00:13:35.35" />
                    <SPLIT distance="650" swimtime="00:14:45.97" />
                    <SPLIT distance="700" swimtime="00:15:53.27" />
                    <SPLIT distance="750" swimtime="00:16:59.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="70" reactiontime="+115" swimtime="00:05:05.93" resultid="19938" heatid="24341" lane="4" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.38" />
                    <SPLIT distance="100" swimtime="00:02:28.34" />
                    <SPLIT distance="150" swimtime="00:03:47.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="28" reactiontime="+109" swimtime="00:06:03.80" resultid="19939" heatid="24368" lane="6" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.51" />
                    <SPLIT distance="100" swimtime="00:02:47.11" />
                    <SPLIT distance="150" swimtime="00:04:28.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="67" reactiontime="+140" swimtime="00:02:20.26" resultid="19940" heatid="24380" lane="4" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="58" reactiontime="+88" swimtime="00:10:27.15" resultid="19941" heatid="24430" lane="1" entrytime="00:10:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.97" />
                    <SPLIT distance="100" swimtime="00:02:45.53" />
                    <SPLIT distance="150" swimtime="00:04:13.10" />
                    <SPLIT distance="200" swimtime="00:05:35.29" />
                    <SPLIT distance="250" swimtime="00:06:55.81" />
                    <SPLIT distance="300" swimtime="00:08:13.75" />
                    <SPLIT distance="350" swimtime="00:09:19.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="57" reactiontime="+111" swimtime="00:04:49.82" resultid="19942" heatid="24447" lane="0" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.22" />
                    <SPLIT distance="100" swimtime="00:02:19.80" />
                    <SPLIT distance="150" swimtime="00:03:35.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="77" reactiontime="+134" swimtime="00:08:37.09" resultid="19943" heatid="24475" lane="2" entrytime="00:08:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.47" />
                    <SPLIT distance="100" swimtime="00:01:59.52" />
                    <SPLIT distance="150" swimtime="00:03:06.18" />
                    <SPLIT distance="200" swimtime="00:04:13.91" />
                    <SPLIT distance="250" swimtime="00:05:21.47" />
                    <SPLIT distance="300" swimtime="00:06:29.82" />
                    <SPLIT distance="350" swimtime="00:07:34.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-11-29" firstname="Edward" gender="M" lastname="Dziekoński" nation="POL" athleteid="22622">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="22623" heatid="24284" lane="2" entrytime="00:00:41.00" />
                <RESULT eventid="14189" points="102" reactiontime="+134" swimtime="00:16:04.63" resultid="22624" heatid="24314" lane="2" entrytime="00:15:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.54" />
                    <SPLIT distance="100" swimtime="00:01:51.45" />
                    <SPLIT distance="150" swimtime="00:02:50.16" />
                    <SPLIT distance="200" swimtime="00:03:49.56" />
                    <SPLIT distance="250" swimtime="00:04:49.78" />
                    <SPLIT distance="300" swimtime="00:05:49.82" />
                    <SPLIT distance="350" swimtime="00:06:51.32" />
                    <SPLIT distance="400" swimtime="00:07:54.05" />
                    <SPLIT distance="450" swimtime="00:08:55.26" />
                    <SPLIT distance="500" swimtime="00:09:58.19" />
                    <SPLIT distance="550" swimtime="00:11:01.24" />
                    <SPLIT distance="600" swimtime="00:12:03.46" />
                    <SPLIT distance="650" swimtime="00:13:05.31" />
                    <SPLIT distance="700" swimtime="00:14:05.88" />
                    <SPLIT distance="750" swimtime="00:15:06.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="76" swimtime="00:00:56.63" resultid="22625" heatid="24330" lane="8" entrytime="00:00:52.00" />
                <RESULT eventid="1273" points="111" reactiontime="+73" swimtime="00:01:37.53" resultid="22626" heatid="24356" lane="9" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="107" reactiontime="+98" swimtime="00:00:46.87" resultid="22627" heatid="24391" lane="2" entrytime="00:00:44.00" />
                <RESULT eventid="1508" points="103" reactiontime="+76" swimtime="00:03:37.47" resultid="22628" heatid="24417" lane="7" entrytime="00:03:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.76" />
                    <SPLIT distance="100" swimtime="00:01:44.19" />
                    <SPLIT distance="150" swimtime="00:02:41.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="56" reactiontime="+104" swimtime="00:02:09.99" resultid="22629" heatid="24437" lane="4" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="100" reactiontime="+103" swimtime="00:07:53.34" resultid="22630" heatid="24476" lane="1" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.97" />
                    <SPLIT distance="100" swimtime="00:01:49.97" />
                    <SPLIT distance="150" swimtime="00:02:50.93" />
                    <SPLIT distance="200" swimtime="00:03:51.40" />
                    <SPLIT distance="250" swimtime="00:04:53.32" />
                    <SPLIT distance="300" swimtime="00:05:54.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-03" firstname="Piotr" gender="M" lastname="Fuliński" nation="POL" athleteid="19756">
              <RESULTS>
                <RESULT eventid="1079" points="470" reactiontime="+86" swimtime="00:00:26.88" resultid="19757" heatid="24294" lane="3" entrytime="00:00:26.50" />
                <RESULT eventid="1273" points="479" swimtime="00:00:59.92" resultid="19758" heatid="24362" lane="5" entrytime="00:00:59.80" />
                <RESULT eventid="1508" points="405" swimtime="00:02:17.78" resultid="19759" heatid="24422" lane="0" entrytime="00:02:19.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.42" />
                    <SPLIT distance="100" swimtime="00:01:05.50" />
                    <SPLIT distance="150" swimtime="00:01:41.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-05-26" firstname="Rafał" gender="M" lastname="Godlewski" nation="POL" athleteid="20967">
              <RESULTS>
                <RESULT eventid="1079" points="230" reactiontime="+72" swimtime="00:00:34.12" resultid="20968" heatid="24286" lane="9" entrytime="00:00:35.80" />
                <RESULT eventid="1239" points="370" swimtime="00:02:56.30" resultid="20969" heatid="24345" lane="1" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                    <SPLIT distance="100" swimtime="00:01:19.55" />
                    <SPLIT distance="150" swimtime="00:02:07.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="429" reactiontime="+64" swimtime="00:01:15.68" resultid="20970" heatid="24384" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="492" swimtime="00:00:32.86" resultid="20971" heatid="24465" lane="8" entrytime="00:00:35.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-08-29" firstname="Łukasz" gender="M" lastname="Grochowski" nation="POL" athleteid="20945">
              <RESULTS>
                <RESULT eventid="1113" points="289" reactiontime="+81" swimtime="00:02:52.38" resultid="20946" heatid="24304" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.04" />
                    <SPLIT distance="100" swimtime="00:01:22.30" />
                    <SPLIT distance="150" swimtime="00:02:10.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="252" swimtime="00:00:37.98" resultid="20947" heatid="24332" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1474" points="240" reactiontime="+64" swimtime="00:01:23.34" resultid="20948" heatid="24405" lane="7" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-05" firstname="Jarosław" gender="M" lastname="Guziński" nation="POL" athleteid="19809">
              <RESULTS>
                <RESULT eventid="1079" points="249" reactiontime="+109" swimtime="00:00:33.21" resultid="19810" heatid="24286" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1273" points="205" reactiontime="+110" swimtime="00:01:19.43" resultid="19811" heatid="24354" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="147" reactiontime="+86" swimtime="00:00:42.11" resultid="19812" heatid="24391" lane="7" entrytime="00:00:45.00" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="19813" heatid="24438" lane="0" entrytime="00:01:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-12-28" firstname="Andrzej" gender="M" lastname="Harenda" nation="POL" athleteid="20929">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="20930" heatid="24289" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="14189" points="202" reactiontime="+106" swimtime="00:12:50.28" resultid="20931" heatid="24315" lane="6" entrytime="00:12:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.73" />
                    <SPLIT distance="100" swimtime="00:01:25.09" />
                    <SPLIT distance="150" swimtime="00:02:11.40" />
                    <SPLIT distance="200" swimtime="00:02:58.95" />
                    <SPLIT distance="250" swimtime="00:03:47.33" />
                    <SPLIT distance="750" swimtime="00:12:05.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="294" reactiontime="+54" swimtime="00:01:10.53" resultid="20932" heatid="24359" lane="3" entrytime="00:01:07.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="20933" heatid="24393" lane="5" entrytime="00:00:34.00" />
                <RESULT eventid="1508" points="215" reactiontime="+76" swimtime="00:02:50.16" resultid="20934" heatid="24420" lane="8" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.24" />
                    <SPLIT distance="150" swimtime="00:02:07.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="229" reactiontime="+84" swimtime="00:05:59.65" resultid="20935" heatid="24478" lane="4" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.34" />
                    <SPLIT distance="150" swimtime="00:02:08.87" />
                    <SPLIT distance="200" swimtime="00:02:56.84" />
                    <SPLIT distance="250" swimtime="00:03:44.16" />
                    <SPLIT distance="300" swimtime="00:04:29.86" />
                    <SPLIT distance="350" swimtime="00:05:17.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-09-27" firstname="Weronika" gender="F" lastname="Kabut" nation="POL" athleteid="23418">
              <RESULTS>
                <RESULT eventid="1062" points="417" reactiontime="+75" swimtime="00:00:31.66" resultid="23419" heatid="24280" lane="5" entrytime="00:00:30.19" />
                <RESULT eventid="1096" points="327" reactiontime="+78" swimtime="00:03:03.06" resultid="23420" heatid="24299" lane="8" entrytime="00:02:52.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.48" />
                    <SPLIT distance="100" swimtime="00:01:26.38" />
                    <SPLIT distance="150" swimtime="00:02:19.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="359" swimtime="00:01:12.73" resultid="23421" heatid="24353" lane="0" entrytime="00:01:06.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="290" swimtime="00:00:36.88" resultid="23422" heatid="24388" lane="5" entrytime="00:00:34.39" />
                <RESULT eventid="1491" points="317" reactiontime="+75" swimtime="00:02:45.57" resultid="23423" heatid="24413" lane="4" entrytime="00:02:31.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.40" />
                    <SPLIT distance="100" swimtime="00:01:16.41" />
                    <SPLIT distance="150" swimtime="00:02:00.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="301" reactiontime="+71" swimtime="00:00:43.83" resultid="23424" heatid="24457" lane="7" entrytime="00:00:42.70" />
                <RESULT eventid="1721" points="274" reactiontime="+71" swimtime="00:06:04.05" resultid="23425" heatid="24472" lane="4" entrytime="00:05:36.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.53" />
                    <SPLIT distance="100" swimtime="00:01:21.43" />
                    <SPLIT distance="150" swimtime="00:02:07.41" />
                    <SPLIT distance="200" swimtime="00:02:54.40" />
                    <SPLIT distance="250" swimtime="00:03:42.86" />
                    <SPLIT distance="300" swimtime="00:04:30.88" />
                    <SPLIT distance="350" swimtime="00:05:19.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-06-11" firstname="Tomasz" gender="M" lastname="Karczewski" nation="POL" athleteid="20283">
              <RESULTS>
                <RESULT eventid="1079" points="338" reactiontime="+91" swimtime="00:00:30.01" resultid="20284" heatid="24289" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="14189" points="272" reactiontime="+97" swimtime="00:11:37.15" resultid="20285" heatid="24316" lane="0" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                    <SPLIT distance="100" swimtime="00:01:23.56" />
                    <SPLIT distance="150" swimtime="00:02:07.41" />
                    <SPLIT distance="200" swimtime="00:02:53.28" />
                    <SPLIT distance="250" swimtime="00:03:37.79" />
                    <SPLIT distance="300" swimtime="00:04:24.30" />
                    <SPLIT distance="350" swimtime="00:05:09.40" />
                    <SPLIT distance="400" swimtime="00:05:53.49" />
                    <SPLIT distance="450" swimtime="00:06:38.21" />
                    <SPLIT distance="500" swimtime="00:07:21.13" />
                    <SPLIT distance="550" swimtime="00:08:06.35" />
                    <SPLIT distance="600" swimtime="00:08:49.87" />
                    <SPLIT distance="650" swimtime="00:09:34.60" />
                    <SPLIT distance="700" swimtime="00:10:17.69" />
                    <SPLIT distance="750" swimtime="00:10:59.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="356" swimtime="00:01:06.17" resultid="20286" heatid="24358" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="361" swimtime="00:00:31.26" resultid="20287" heatid="24395" lane="9" entrytime="00:00:31.12" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-08-03" firstname="Lidia" gender="F" lastname="Kosek" nation="POL" athleteid="22636">
              <RESULTS>
                <RESULT eventid="1062" points="316" reactiontime="+76" swimtime="00:00:34.72" resultid="22637" heatid="24277" lane="4" entrytime="00:00:38.10" />
                <RESULT eventid="1222" points="220" reactiontime="+88" swimtime="00:03:50.23" resultid="22638" heatid="24338" lane="4" entrytime="00:04:05.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.45" />
                    <SPLIT distance="100" swimtime="00:01:51.88" />
                    <SPLIT distance="150" swimtime="00:02:50.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="237" reactiontime="+63" swimtime="00:03:02.52" resultid="22639" heatid="24411" lane="3" entrytime="00:03:20.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                    <SPLIT distance="100" swimtime="00:01:29.33" />
                    <SPLIT distance="150" swimtime="00:02:16.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="191" swimtime="00:06:50.40" resultid="22640" heatid="24471" lane="0" entrytime="00:07:15.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.27" />
                    <SPLIT distance="100" swimtime="00:01:35.45" />
                    <SPLIT distance="150" swimtime="00:02:28.25" />
                    <SPLIT distance="200" swimtime="00:03:21.26" />
                    <SPLIT distance="250" swimtime="00:04:16.22" />
                    <SPLIT distance="300" swimtime="00:05:09.79" />
                    <SPLIT distance="350" swimtime="00:06:02.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-08-12" firstname="Yevhenii" gender="M" lastname="Koshyl" nation="POL" athleteid="20306">
              <RESULTS>
                <RESULT eventid="1079" points="562" reactiontime="+86" swimtime="00:00:25.33" resultid="20307" heatid="24295" lane="4" entrytime="00:00:25.88" />
                <RESULT eventid="1273" points="582" swimtime="00:00:56.17" resultid="20308" heatid="24363" lane="2" entrytime="00:00:58.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="446" swimtime="00:02:13.44" resultid="20309" heatid="24423" lane="4" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.35" />
                    <SPLIT distance="100" swimtime="00:00:59.70" />
                    <SPLIT distance="150" swimtime="00:01:35.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="345" swimtime="00:01:10.99" resultid="20310" heatid="24441" lane="9" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-08-26" firstname="Adrian" gender="M" lastname="Kozioł" nation="POL" athleteid="22657">
              <RESULTS>
                <RESULT eventid="1079" points="406" reactiontime="+86" swimtime="00:00:28.22" resultid="22658" heatid="24292" lane="0" entrytime="00:00:28.50" />
                <RESULT eventid="1273" points="378" swimtime="00:01:04.84" resultid="22659" heatid="24360" lane="1" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="419" swimtime="00:00:29.74" resultid="22660" heatid="24395" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="22661" heatid="24440" lane="5" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-07-31" firstname="Piotr" gender="M" lastname="Krogulec" nation="POL" athleteid="22678">
              <RESULTS>
                <RESULT eventid="1079" points="441" reactiontime="+85" swimtime="00:00:27.46" resultid="22679" heatid="24292" lane="5" entrytime="00:00:28.00" />
                <RESULT eventid="1113" points="396" reactiontime="+85" swimtime="00:02:35.15" resultid="22680" heatid="24306" lane="9" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                    <SPLIT distance="100" swimtime="00:01:11.69" />
                    <SPLIT distance="150" swimtime="00:01:57.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="440" swimtime="00:00:31.55" resultid="22681" heatid="24334" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="22682" heatid="24361" lane="4" entrytime="00:01:03.00" />
                <RESULT eventid="1440" points="421" swimtime="00:00:29.70" resultid="22683" heatid="24394" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1474" points="389" swimtime="00:01:11.01" resultid="22684" heatid="24407" lane="3" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="22685" heatid="24451" lane="0" entrytime="00:02:40.00" />
                <RESULT eventid="1681" points="332" swimtime="00:00:37.46" resultid="22686" heatid="24465" lane="9" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-05-11" firstname="Joanna" gender="F" lastname="Krowicka" nation="POL" athleteid="23403">
              <RESULTS>
                <RESULT eventid="1222" status="DNS" swimtime="00:00:00.00" resultid="23404" heatid="24339" lane="0" entrytime="00:03:48.68" />
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="23405" heatid="24350" lane="9" entrytime="00:01:30.40" />
                <RESULT eventid="1388" status="DNS" swimtime="00:00:00.00" resultid="23406" heatid="24378" lane="0" entrytime="00:01:44.18" />
                <RESULT eventid="1423" status="DNS" swimtime="00:00:00.00" resultid="23407" heatid="24386" lane="4" entrytime="00:00:49.19" />
                <RESULT eventid="1664" status="DNS" swimtime="00:00:00.00" resultid="23408" heatid="24456" lane="7" entrytime="00:00:47.02" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-11-12" firstname="Jakub" gender="M" lastname="Kędzierski" nation="POL" athleteid="19784">
              <RESULTS>
                <RESULT eventid="1205" points="307" swimtime="00:00:35.54" resultid="19785" heatid="24332" lane="5" entrytime="00:00:38.00" />
                <RESULT eventid="1273" points="354" swimtime="00:01:06.31" resultid="19786" heatid="24357" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="287" swimtime="00:02:34.63" resultid="19787" heatid="24420" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.48" />
                    <SPLIT distance="100" swimtime="00:01:12.46" />
                    <SPLIT distance="150" swimtime="00:01:53.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-08-29" firstname="Hracki" gender="M" lastname="Libor" nation="CZE" athleteid="20266">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="20267" heatid="24288" lane="6" entrytime="00:00:31.50" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="20268" heatid="24345" lane="9" entrytime="00:03:05.00" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="20269" heatid="24359" lane="0" entrytime="00:01:09.50" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="20270" heatid="24383" lane="1" entrytime="00:01:27.50" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="20271" heatid="24420" lane="1" entrytime="00:02:35.50" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="20272" heatid="24462" lane="0" entrytime="00:00:42.25" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="20273" heatid="24479" lane="7" entrytime="00:05:36.25" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-10-24" firstname="Andrzej" gender="M" lastname="Marszałek" nation="POL" athleteid="19944">
              <RESULTS>
                <RESULT eventid="1079" points="118" reactiontime="+98" swimtime="00:00:42.63" resultid="19945" heatid="24284" lane="8" entrytime="00:00:44.00" />
                <RESULT eventid="14189" points="112" reactiontime="+102" swimtime="00:15:35.58" resultid="19946" heatid="24314" lane="7" entrytime="00:16:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.79" />
                    <SPLIT distance="100" swimtime="00:01:48.42" />
                    <SPLIT distance="150" swimtime="00:02:45.27" />
                    <SPLIT distance="200" swimtime="00:03:42.41" />
                    <SPLIT distance="250" swimtime="00:04:39.94" />
                    <SPLIT distance="300" swimtime="00:05:38.14" />
                    <SPLIT distance="350" swimtime="00:06:36.38" />
                    <SPLIT distance="400" swimtime="00:07:35.36" />
                    <SPLIT distance="450" swimtime="00:08:33.62" />
                    <SPLIT distance="500" swimtime="00:09:33.10" />
                    <SPLIT distance="550" swimtime="00:10:32.93" />
                    <SPLIT distance="600" swimtime="00:11:33.50" />
                    <SPLIT distance="650" swimtime="00:12:33.78" />
                    <SPLIT distance="700" swimtime="00:13:34.75" />
                    <SPLIT distance="750" swimtime="00:14:35.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="102" reactiontime="+79" swimtime="00:01:40.14" resultid="19947" heatid="24355" lane="3" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="69" reactiontime="+75" swimtime="00:00:54.15" resultid="19948" heatid="24391" lane="9" entrytime="00:00:49.00" />
                <RESULT eventid="1508" points="100" reactiontime="+74" swimtime="00:03:39.13" resultid="19949" heatid="24417" lane="0" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.68" />
                    <SPLIT distance="100" swimtime="00:01:45.13" />
                    <SPLIT distance="150" swimtime="00:02:43.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="108" reactiontime="+79" swimtime="00:07:40.72" resultid="19950" heatid="24476" lane="0" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.00" />
                    <SPLIT distance="100" swimtime="00:01:48.05" />
                    <SPLIT distance="150" swimtime="00:02:45.80" />
                    <SPLIT distance="200" swimtime="00:03:43.71" />
                    <SPLIT distance="250" swimtime="00:04:42.45" />
                    <SPLIT distance="300" swimtime="00:05:41.87" />
                    <SPLIT distance="350" swimtime="00:06:42.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-05-24" firstname="Bogdan" gender="M" lastname="Martyniuk" nation="POL" athleteid="22648">
              <RESULTS>
                <RESULT eventid="1079" points="183" reactiontime="+115" swimtime="00:00:36.79" resultid="22649" heatid="24282" lane="4" />
                <RESULT eventid="1113" points="96" reactiontime="+113" swimtime="00:04:08.81" resultid="22650" heatid="24300" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.65" />
                    <SPLIT distance="100" swimtime="00:02:05.84" />
                    <SPLIT distance="150" swimtime="00:03:16.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="99" swimtime="00:00:51.78" resultid="22651" heatid="24328" lane="1" />
                <RESULT eventid="1273" points="106" reactiontime="+83" swimtime="00:01:38.89" resultid="22652" heatid="24355" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="76" reactiontime="+69" swimtime="00:00:52.38" resultid="22653" heatid="24390" lane="8" />
                <RESULT eventid="1508" points="82" reactiontime="+78" swimtime="00:03:54.22" resultid="22654" heatid="24415" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:51.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="22655" heatid="24437" lane="0" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="22656" heatid="24459" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-03-09" firstname="Aleksandra" gender="F" lastname="Morkisz" nation="POL" athleteid="19788">
              <RESULTS>
                <RESULT eventid="1222" points="367" reactiontime="+84" swimtime="00:03:14.14" resultid="19789" heatid="24340" lane="8" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.62" />
                    <SPLIT distance="100" swimtime="00:01:33.78" />
                    <SPLIT distance="150" swimtime="00:02:25.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="370" reactiontime="+54" swimtime="00:01:29.26" resultid="19790" heatid="24378" lane="4" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="335" reactiontime="+67" swimtime="00:02:42.63" resultid="19791" heatid="24412" lane="6" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.95" />
                    <SPLIT distance="100" swimtime="00:01:18.98" />
                    <SPLIT distance="150" swimtime="00:02:01.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="364" swimtime="00:00:41.16" resultid="19792" heatid="24457" lane="1" entrytime="00:00:43.00" />
                <RESULT eventid="1721" points="326" reactiontime="+59" swimtime="00:05:43.38" resultid="19793" heatid="24472" lane="7" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.80" />
                    <SPLIT distance="100" swimtime="00:01:19.48" />
                    <SPLIT distance="150" swimtime="00:02:02.88" />
                    <SPLIT distance="200" swimtime="00:02:47.01" />
                    <SPLIT distance="250" swimtime="00:03:31.56" />
                    <SPLIT distance="300" swimtime="00:04:16.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-02-13" firstname="Steran" gender="M" lastname="Niedzielski" nation="POL" athleteid="19794">
              <RESULTS>
                <RESULT eventid="1079" points="145" reactiontime="+115" swimtime="00:00:39.80" resultid="19795" heatid="24285" lane="6" entrytime="00:00:37.00" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="19796" heatid="24330" lane="0" entrytime="00:00:52.00" />
                <RESULT eventid="1239" points="139" reactiontime="+76" swimtime="00:04:04.26" resultid="19797" heatid="24342" lane="6" entrytime="00:04:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.87" />
                    <SPLIT distance="100" swimtime="00:01:58.43" />
                    <SPLIT distance="150" swimtime="00:03:03.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="19798" heatid="24381" lane="7" entrytime="00:01:51.00" />
                <RESULT eventid="1681" points="150" reactiontime="+63" swimtime="00:00:48.75" resultid="19799" heatid="24460" lane="2" entrytime="00:00:52.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-09-24" firstname="Szymon" gender="M" lastname="Parafiniak" nation="POL" athleteid="22641">
              <RESULTS>
                <RESULT eventid="1079" points="304" reactiontime="+84" swimtime="00:00:31.08" resultid="22642" heatid="24290" lane="1" entrytime="00:00:29.90" />
                <RESULT eventid="1273" points="224" reactiontime="+77" swimtime="00:01:17.20" resultid="22643" heatid="24359" lane="4" entrytime="00:01:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="22644" heatid="24393" lane="0" entrytime="00:00:35.50" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="22645" heatid="24422" lane="9" entrytime="00:02:20.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-03-27" firstname="Jakub" gender="M" lastname="Pogorzelec" nation="POL" athleteid="21506">
              <RESULTS>
                <RESULT eventid="1079" points="474" reactiontime="+87" swimtime="00:00:26.80" resultid="21507" heatid="24292" lane="2" entrytime="00:00:28.00" />
                <RESULT eventid="1113" points="285" reactiontime="+97" swimtime="00:02:53.03" resultid="21508" heatid="24300" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.26" />
                    <SPLIT distance="100" swimtime="00:01:13.13" />
                    <SPLIT distance="150" swimtime="00:02:10.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="413" reactiontime="+80" swimtime="00:00:32.22" resultid="21509" heatid="24334" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="1273" points="477" swimtime="00:01:00.00" resultid="21510" heatid="24360" lane="6" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="409" swimtime="00:00:29.99" resultid="21511" heatid="24394" lane="0" entrytime="00:00:33.00" />
                <RESULT eventid="1508" points="327" swimtime="00:02:28.05" resultid="21512" heatid="24421" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                    <SPLIT distance="100" swimtime="00:01:08.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-10" firstname="Michał" gender="M" lastname="Rudziński" nation="POL" athleteid="20922">
              <RESULTS>
                <RESULT eventid="1079" points="168" reactiontime="+126" swimtime="00:00:37.88" resultid="20923" heatid="24285" lane="3" entrytime="00:00:36.82" />
                <RESULT eventid="1239" points="208" reactiontime="+88" swimtime="00:03:33.77" resultid="20924" heatid="24341" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.16" />
                    <SPLIT distance="100" swimtime="00:01:42.31" />
                    <SPLIT distance="150" swimtime="00:02:38.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="135" reactiontime="+87" swimtime="00:03:37.17" resultid="20925" heatid="24369" lane="3" entrytime="00:03:45.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.15" />
                    <SPLIT distance="100" swimtime="00:01:42.23" />
                    <SPLIT distance="150" swimtime="00:02:39.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="176" reactiontime="+44" swimtime="00:00:39.68" resultid="20926" heatid="24391" lane="4" entrytime="00:00:39.78" />
                <RESULT eventid="1613" points="160" reactiontime="+64" swimtime="00:01:31.65" resultid="20927" heatid="24438" lane="3" entrytime="00:01:35.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="132" reactiontime="+80" swimtime="00:07:11.79" resultid="20928" heatid="24476" lane="8" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.89" />
                    <SPLIT distance="100" swimtime="00:01:39.26" />
                    <SPLIT distance="150" swimtime="00:02:34.96" />
                    <SPLIT distance="200" swimtime="00:03:33.01" />
                    <SPLIT distance="250" swimtime="00:04:27.70" />
                    <SPLIT distance="300" swimtime="00:05:24.01" />
                    <SPLIT distance="350" swimtime="00:06:18.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-06-14" firstname="Andrzej" gender="M" lastname="Rusinowicz" nation="POL" athleteid="20936">
              <RESULTS>
                <RESULT eventid="1113" points="67" reactiontime="+109" swimtime="00:04:39.88" resultid="20937" heatid="24301" lane="7" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.39" />
                    <SPLIT distance="100" swimtime="00:02:14.36" />
                    <SPLIT distance="150" swimtime="00:03:32.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14207" reactiontime="+123" status="OTL" swimtime="00:36:30.91" resultid="20938" heatid="24320" lane="1" entrytime="00:35:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.96" />
                    <SPLIT distance="100" swimtime="00:02:13.94" />
                    <SPLIT distance="150" swimtime="00:03:26.97" />
                    <SPLIT distance="200" swimtime="00:04:38.76" />
                    <SPLIT distance="250" swimtime="00:05:51.56" />
                    <SPLIT distance="300" swimtime="00:07:02.49" />
                    <SPLIT distance="350" swimtime="00:08:15.50" />
                    <SPLIT distance="400" swimtime="00:09:29.30" />
                    <SPLIT distance="450" swimtime="00:10:43.63" />
                    <SPLIT distance="500" swimtime="00:11:59.77" />
                    <SPLIT distance="550" swimtime="00:13:12.75" />
                    <SPLIT distance="600" swimtime="00:14:25.18" />
                    <SPLIT distance="650" swimtime="00:15:39.73" />
                    <SPLIT distance="700" swimtime="00:16:51.66" />
                    <SPLIT distance="750" swimtime="00:18:05.75" />
                    <SPLIT distance="800" swimtime="00:19:17.43" />
                    <SPLIT distance="850" swimtime="00:20:32.13" />
                    <SPLIT distance="900" swimtime="00:21:43.72" />
                    <SPLIT distance="950" swimtime="00:22:58.73" />
                    <SPLIT distance="1000" swimtime="00:24:10.16" />
                    <SPLIT distance="1050" swimtime="00:25:24.66" />
                    <SPLIT distance="1100" swimtime="00:26:37.06" />
                    <SPLIT distance="1150" swimtime="00:27:51.61" />
                    <SPLIT distance="1200" swimtime="00:29:04.45" />
                    <SPLIT distance="1250" swimtime="00:30:19.70" />
                    <SPLIT distance="1350" swimtime="00:32:51.30" />
                    <SPLIT distance="1400" swimtime="00:34:02.85" />
                    <SPLIT distance="1450" swimtime="00:35:19.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="20939" heatid="24329" lane="3" entrytime="00:00:57.00" />
                <RESULT eventid="1239" points="69" reactiontime="+97" swimtime="00:05:07.99" resultid="20940" heatid="24342" lane="1" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.72" />
                    <SPLIT distance="100" swimtime="00:02:30.84" />
                    <SPLIT distance="150" swimtime="00:03:52.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="62" reactiontime="+80" swimtime="00:02:10.33" resultid="20941" heatid="24403" lane="3" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="57" reactiontime="+82" swimtime="00:10:31.79" resultid="20942" heatid="24430" lane="7" entrytime="00:10:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.41" />
                    <SPLIT distance="100" swimtime="00:02:30.91" />
                    <SPLIT distance="150" swimtime="00:03:55.04" />
                    <SPLIT distance="200" swimtime="00:05:20.86" />
                    <SPLIT distance="250" swimtime="00:06:46.22" />
                    <SPLIT distance="300" swimtime="00:08:09.19" />
                    <SPLIT distance="350" swimtime="00:09:22.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="60" reactiontime="+86" swimtime="00:04:45.24" resultid="20943" heatid="24447" lane="7" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.74" />
                    <SPLIT distance="100" swimtime="00:02:17.96" />
                    <SPLIT distance="150" swimtime="00:03:33.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="20944" heatid="24475" lane="7" entrytime="00:08:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-08-03" firstname="Roman" gender="M" lastname="Saienko" nation="POL" athleteid="20301">
              <RESULTS>
                <RESULT eventid="1079" points="521" reactiontime="+71" swimtime="00:00:25.97" resultid="20302" heatid="24295" lane="5" entrytime="00:00:25.89" />
                <RESULT eventid="1273" points="497" swimtime="00:00:59.21" resultid="20303" heatid="24363" lane="6" entrytime="00:00:58.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="410" reactiontime="+53" swimtime="00:02:17.24" resultid="20304" heatid="24423" lane="7" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.11" />
                    <SPLIT distance="100" swimtime="00:01:03.76" />
                    <SPLIT distance="150" swimtime="00:01:40.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="424" swimtime="00:01:06.31" resultid="20305" heatid="24441" lane="0" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-05" firstname="Tomasz" gender="M" lastname="Sitkowski" nation="POL" athleteid="23090">
              <RESULTS>
                <RESULT eventid="1079" points="374" reactiontime="+91" swimtime="00:00:29.00" resultid="23091" heatid="24291" lane="2" entrytime="00:00:29.00" />
                <RESULT eventid="1205" points="285" swimtime="00:00:36.44" resultid="23092" heatid="24333" lane="1" entrytime="00:00:36.30" />
                <RESULT eventid="1273" points="326" swimtime="00:01:08.15" resultid="23093" heatid="24360" lane="9" entrytime="00:01:07.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="248" reactiontime="+125" swimtime="00:01:22.44" resultid="23094" heatid="24405" lane="4" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-02-10" firstname="Jacek" gender="M" lastname="Sokulski" nation="POL" athleteid="22666">
              <RESULTS>
                <RESULT eventid="1079" points="654" reactiontime="+68" swimtime="00:00:24.08" resultid="22667" heatid="24296" lane="6" entrytime="00:00:24.50" />
                <RESULT eventid="1205" points="587" reactiontime="+64" swimtime="00:00:28.66" resultid="22668" heatid="24336" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="1273" points="678" reactiontime="+68" swimtime="00:00:53.38" resultid="22669" heatid="24365" lane="7" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="708" reactiontime="+72" swimtime="00:00:24.98" resultid="22670" heatid="24398" lane="3" entrytime="00:00:26.00" />
                <RESULT eventid="1613" points="612" swimtime="00:00:58.66" resultid="22671" heatid="24442" lane="6" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-07-22" firstname="Ireneusz" gender="M" lastname="Stachurski" nation="POL" athleteid="19980">
              <RESULTS>
                <RESULT eventid="1079" points="205" reactiontime="+103" swimtime="00:00:35.44" resultid="19981" heatid="24286" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="14189" points="165" reactiontime="+119" swimtime="00:13:43.92" resultid="19982" heatid="24313" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.10" />
                    <SPLIT distance="100" swimtime="00:01:31.50" />
                    <SPLIT distance="150" swimtime="00:02:23.45" />
                    <SPLIT distance="200" swimtime="00:03:16.08" />
                    <SPLIT distance="250" swimtime="00:04:09.43" />
                    <SPLIT distance="300" swimtime="00:05:01.75" />
                    <SPLIT distance="350" swimtime="00:05:55.65" />
                    <SPLIT distance="400" swimtime="00:06:48.84" />
                    <SPLIT distance="450" swimtime="00:07:42.00" />
                    <SPLIT distance="500" swimtime="00:08:34.19" />
                    <SPLIT distance="550" swimtime="00:09:27.64" />
                    <SPLIT distance="600" swimtime="00:10:20.55" />
                    <SPLIT distance="650" swimtime="00:11:12.98" />
                    <SPLIT distance="700" swimtime="00:12:05.15" />
                    <SPLIT distance="750" swimtime="00:12:56.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="19983" heatid="24390" lane="1" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="19984" heatid="24419" lane="0" entrytime="00:02:54.00" />
                <RESULT eventid="1613" points="107" reactiontime="+69" swimtime="00:01:44.75" resultid="19985" heatid="24438" lane="6" entrytime="00:01:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="171" reactiontime="+84" swimtime="00:06:35.87" resultid="19986" heatid="24477" lane="6" entrytime="00:06:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.64" />
                    <SPLIT distance="100" swimtime="00:01:30.26" />
                    <SPLIT distance="150" swimtime="00:02:20.44" />
                    <SPLIT distance="200" swimtime="00:03:12.65" />
                    <SPLIT distance="250" swimtime="00:04:03.65" />
                    <SPLIT distance="300" swimtime="00:04:55.95" />
                    <SPLIT distance="350" swimtime="00:05:47.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-07" firstname="Michał" gender="M" lastname="Urbański" nation="POL" athleteid="19951">
              <RESULTS>
                <RESULT eventid="14207" points="451" reactiontime="+84" swimtime="00:18:55.69" resultid="19952" heatid="24322" lane="4" entrytime="00:18:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.81" />
                    <SPLIT distance="100" swimtime="00:01:06.80" />
                    <SPLIT distance="150" swimtime="00:01:42.68" />
                    <SPLIT distance="200" swimtime="00:02:19.17" />
                    <SPLIT distance="250" swimtime="00:02:56.06" />
                    <SPLIT distance="300" swimtime="00:03:33.44" />
                    <SPLIT distance="350" swimtime="00:04:10.72" />
                    <SPLIT distance="400" swimtime="00:04:48.18" />
                    <SPLIT distance="450" swimtime="00:05:26.11" />
                    <SPLIT distance="500" swimtime="00:06:03.98" />
                    <SPLIT distance="550" swimtime="00:06:41.97" />
                    <SPLIT distance="600" swimtime="00:07:20.31" />
                    <SPLIT distance="650" swimtime="00:07:58.88" />
                    <SPLIT distance="700" swimtime="00:08:37.43" />
                    <SPLIT distance="750" swimtime="00:09:15.93" />
                    <SPLIT distance="800" swimtime="00:09:54.42" />
                    <SPLIT distance="850" swimtime="00:10:33.36" />
                    <SPLIT distance="900" swimtime="00:11:12.43" />
                    <SPLIT distance="950" swimtime="00:11:51.66" />
                    <SPLIT distance="1000" swimtime="00:12:30.56" />
                    <SPLIT distance="1050" swimtime="00:13:09.18" />
                    <SPLIT distance="1100" swimtime="00:13:47.39" />
                    <SPLIT distance="1150" swimtime="00:14:26.08" />
                    <SPLIT distance="1200" swimtime="00:15:04.78" />
                    <SPLIT distance="1250" swimtime="00:15:43.62" />
                    <SPLIT distance="1300" swimtime="00:16:22.18" />
                    <SPLIT distance="1350" swimtime="00:17:00.71" />
                    <SPLIT distance="1400" swimtime="00:17:39.84" />
                    <SPLIT distance="1450" swimtime="00:18:18.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="552" reactiontime="+68" swimtime="00:02:34.40" resultid="19953" heatid="24346" lane="4" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.89" />
                    <SPLIT distance="100" swimtime="00:01:14.07" />
                    <SPLIT distance="150" swimtime="00:01:53.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="19954" heatid="24424" lane="3" entrytime="00:02:01.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1938-04-28" firstname="Andrzej" gender="M" lastname="Wiśniewski" nation="POL" athleteid="22646">
              <RESULTS>
                <RESULT eventid="14207" points="65" reactiontime="+121" swimtime="00:35:55.33" resultid="22647" heatid="24320" lane="8" entrytime="00:41:37.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.12" />
                    <SPLIT distance="100" swimtime="00:02:13.23" />
                    <SPLIT distance="150" swimtime="00:03:24.23" />
                    <SPLIT distance="200" swimtime="00:04:36.00" />
                    <SPLIT distance="250" swimtime="00:05:46.24" />
                    <SPLIT distance="300" swimtime="00:06:57.07" />
                    <SPLIT distance="350" swimtime="00:08:07.98" />
                    <SPLIT distance="400" swimtime="00:09:18.76" />
                    <SPLIT distance="450" swimtime="00:10:29.78" />
                    <SPLIT distance="500" swimtime="00:11:40.48" />
                    <SPLIT distance="550" swimtime="00:12:51.24" />
                    <SPLIT distance="600" swimtime="00:14:02.05" />
                    <SPLIT distance="650" swimtime="00:15:13.71" />
                    <SPLIT distance="700" swimtime="00:16:25.51" />
                    <SPLIT distance="750" swimtime="00:17:37.01" />
                    <SPLIT distance="800" swimtime="00:18:50.01" />
                    <SPLIT distance="850" swimtime="00:20:02.46" />
                    <SPLIT distance="900" swimtime="00:21:15.51" />
                    <SPLIT distance="950" swimtime="00:22:27.53" />
                    <SPLIT distance="1000" swimtime="00:23:40.28" />
                    <SPLIT distance="1050" swimtime="00:24:53.06" />
                    <SPLIT distance="1100" swimtime="00:26:06.75" />
                    <SPLIT distance="1150" swimtime="00:27:21.78" />
                    <SPLIT distance="1200" swimtime="00:28:36.40" />
                    <SPLIT distance="1250" swimtime="00:29:49.78" />
                    <SPLIT distance="1300" swimtime="00:31:04.23" />
                    <SPLIT distance="1350" swimtime="00:32:17.99" />
                    <SPLIT distance="1400" swimtime="00:33:31.08" />
                    <SPLIT distance="1450" swimtime="00:34:43.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-12-04" firstname="Angelika" gender="F" lastname="Wróbel" nation="POL" athleteid="22662">
              <RESULTS>
                <RESULT eventid="1062" points="568" reactiontime="+84" swimtime="00:00:28.58" resultid="22663" heatid="24281" lane="6" entrytime="00:00:28.65" />
                <RESULT eventid="1256" points="564" reactiontime="+73" swimtime="00:01:02.56" resultid="22664" heatid="24353" lane="3" entrytime="00:01:01.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="502" reactiontime="+80" swimtime="00:02:22.08" resultid="22665" heatid="24414" lane="3" entrytime="00:02:15.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                    <SPLIT distance="100" swimtime="00:01:08.92" />
                    <SPLIT distance="150" swimtime="00:01:44.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-02-01" firstname="Jolanta" gender="F" lastname="Zawadzka" nation="POL" athleteid="22631">
              <RESULTS>
                <RESULT eventid="1096" points="208" reactiontime="+89" swimtime="00:03:32.84" resultid="22632" heatid="24298" lane="9" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.12" />
                    <SPLIT distance="100" swimtime="00:01:41.12" />
                    <SPLIT distance="150" swimtime="00:02:40.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="256" reactiontime="+65" swimtime="00:01:40.95" resultid="22633" heatid="24377" lane="4" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="222" reactiontime="+65" swimtime="00:00:40.34" resultid="22634" heatid="24387" lane="2" entrytime="00:00:41.00" />
                <RESULT eventid="1664" points="272" swimtime="00:00:45.33" resultid="22635" heatid="24457" lane="9" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-08-29" firstname="Leszek" gender="M" lastname="Zawadzki" nation="POL" athleteid="19779">
              <RESULTS>
                <RESULT eventid="1079" points="328" reactiontime="+112" swimtime="00:00:30.29" resultid="19780" heatid="24291" lane="7" entrytime="00:00:29.00" />
                <RESULT eventid="14207" reactiontime="+123" status="OTL" swimtime="00:23:26.67" resultid="19781" heatid="24322" lane="8" entrytime="00:20:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                    <SPLIT distance="100" swimtime="00:01:14.79" />
                    <SPLIT distance="150" swimtime="00:01:56.50" />
                    <SPLIT distance="200" swimtime="00:02:39.30" />
                    <SPLIT distance="250" swimtime="00:03:23.03" />
                    <SPLIT distance="300" swimtime="00:04:07.21" />
                    <SPLIT distance="350" swimtime="00:04:52.21" />
                    <SPLIT distance="400" swimtime="00:05:37.41" />
                    <SPLIT distance="450" swimtime="00:06:23.33" />
                    <SPLIT distance="500" swimtime="00:07:09.61" />
                    <SPLIT distance="550" swimtime="00:07:56.03" />
                    <SPLIT distance="600" swimtime="00:08:42.32" />
                    <SPLIT distance="650" swimtime="00:09:29.33" />
                    <SPLIT distance="700" swimtime="00:10:17.33" />
                    <SPLIT distance="750" swimtime="00:11:04.79" />
                    <SPLIT distance="800" swimtime="00:11:52.52" />
                    <SPLIT distance="850" swimtime="00:12:40.18" />
                    <SPLIT distance="900" swimtime="00:13:28.35" />
                    <SPLIT distance="950" swimtime="00:14:15.63" />
                    <SPLIT distance="1000" swimtime="00:15:04.07" />
                    <SPLIT distance="1050" swimtime="00:15:52.40" />
                    <SPLIT distance="1100" swimtime="00:16:40.96" />
                    <SPLIT distance="1150" swimtime="00:17:29.45" />
                    <SPLIT distance="1200" swimtime="00:18:18.63" />
                    <SPLIT distance="1250" swimtime="00:19:06.60" />
                    <SPLIT distance="1300" swimtime="00:19:54.19" />
                    <SPLIT distance="1350" swimtime="00:20:42.02" />
                    <SPLIT distance="1400" swimtime="00:21:28.13" />
                    <SPLIT distance="1450" swimtime="00:22:39.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="300" reactiontime="+90" swimtime="00:02:32.22" resultid="19782" heatid="24417" lane="5" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                    <SPLIT distance="100" swimtime="00:01:10.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="286" reactiontime="+106" swimtime="00:05:33.98" resultid="19783" heatid="24476" lane="7" entrytime="00:07:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                    <SPLIT distance="100" swimtime="00:01:14.31" />
                    <SPLIT distance="150" swimtime="00:01:55.78" />
                    <SPLIT distance="200" swimtime="00:02:38.59" />
                    <SPLIT distance="250" swimtime="00:03:22.24" />
                    <SPLIT distance="300" swimtime="00:04:07.37" />
                    <SPLIT distance="350" swimtime="00:04:52.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-11-08" firstname="Tomasz" gender="M" lastname="Zdebel" nation="POL" athleteid="23087">
              <RESULTS>
                <RESULT eventid="1406" points="291" reactiontime="+68" swimtime="00:01:26.12" resultid="23088" heatid="24382" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="23089" heatid="24464" lane="9" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-11-01" firstname="Stanisław" gender="M" lastname="Zejfert" nation="POL" athleteid="20262">
              <RESULTS>
                <RESULT eventid="1205" points="141" swimtime="00:00:46.10" resultid="20263" heatid="24328" lane="3" />
                <RESULT eventid="1474" points="127" reactiontime="+93" swimtime="00:01:42.98" resultid="20264" heatid="24403" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="115" reactiontime="+91" swimtime="00:03:49.83" resultid="20265" heatid="24446" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.45" />
                    <SPLIT distance="100" swimtime="00:01:54.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-04-24" firstname="Włodzimierz" gender="M" lastname="Zieleziński" nation="POL" athleteid="20958">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="20959" heatid="24286" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="14207" points="128" reactiontime="+142" swimtime="00:28:47.97" resultid="20960" heatid="24320" lane="2" entrytime="00:29:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.77" />
                    <SPLIT distance="100" swimtime="00:01:37.94" />
                    <SPLIT distance="150" swimtime="00:02:33.43" />
                    <SPLIT distance="200" swimtime="00:03:30.70" />
                    <SPLIT distance="250" swimtime="00:04:28.94" />
                    <SPLIT distance="300" swimtime="00:05:26.29" />
                    <SPLIT distance="350" swimtime="00:06:24.93" />
                    <SPLIT distance="400" swimtime="00:07:23.47" />
                    <SPLIT distance="450" swimtime="00:08:21.28" />
                    <SPLIT distance="500" swimtime="00:09:20.85" />
                    <SPLIT distance="550" swimtime="00:10:18.78" />
                    <SPLIT distance="600" swimtime="00:11:17.21" />
                    <SPLIT distance="650" swimtime="00:12:15.81" />
                    <SPLIT distance="700" swimtime="00:13:13.86" />
                    <SPLIT distance="750" swimtime="00:14:12.50" />
                    <SPLIT distance="800" swimtime="00:15:11.67" />
                    <SPLIT distance="850" swimtime="00:18:10.05" />
                    <SPLIT distance="900" swimtime="00:17:10.28" />
                    <SPLIT distance="950" swimtime="00:20:08.00" />
                    <SPLIT distance="1000" swimtime="00:19:08.42" />
                    <SPLIT distance="1050" swimtime="00:22:04.45" />
                    <SPLIT distance="1100" swimtime="00:21:06.37" />
                    <SPLIT distance="1150" swimtime="00:24:01.16" />
                    <SPLIT distance="1200" swimtime="00:23:02.91" />
                    <SPLIT distance="1250" swimtime="00:25:57.74" />
                    <SPLIT distance="1300" swimtime="00:25:01.49" />
                    <SPLIT distance="1350" swimtime="00:27:53.91" />
                    <SPLIT distance="1400" swimtime="00:26:55.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="20961" heatid="24331" lane="8" entrytime="00:00:44.00" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="20962" heatid="24356" lane="6" entrytime="00:01:25.00" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="20963" heatid="24404" lane="3" entrytime="00:01:40.00" />
                <RESULT eventid="1508" points="136" reactiontime="+93" swimtime="00:03:18.22" resultid="20964" heatid="24417" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                    <SPLIT distance="100" swimtime="00:01:30.22" />
                    <SPLIT distance="150" swimtime="00:02:24.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="20965" heatid="24448" lane="3" entrytime="00:03:40.00" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="20966" heatid="24477" lane="8" entrytime="00:06:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-02-03" firstname="Damian" gender="M" lastname="Ziółkowski" nation="POL" athleteid="20949">
              <RESULTS>
                <RESULT eventid="1079" points="380" reactiontime="+82" swimtime="00:00:28.85" resultid="20950" heatid="24287" lane="3" entrytime="00:00:32.90" />
                <RESULT eventid="1440" points="346" reactiontime="+69" swimtime="00:00:31.72" resultid="20951" heatid="24393" lane="2" entrytime="00:00:34.17" />
                <RESULT eventid="1508" points="318" reactiontime="+73" swimtime="00:02:29.41" resultid="20952" heatid="24420" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                    <SPLIT distance="100" swimtime="00:01:10.61" />
                    <SPLIT distance="150" swimtime="00:01:50.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="287" reactiontime="+71" swimtime="00:01:15.51" resultid="20953" heatid="24439" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-11-10" firstname="Andrzej" gender="M" lastname="Łopuszynski" nation="POL" athleteid="19814">
              <RESULTS>
                <RESULT eventid="1113" points="111" reactiontime="+105" swimtime="00:03:56.87" resultid="19815" heatid="24302" lane="8" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.33" />
                    <SPLIT distance="100" swimtime="00:01:52.83" />
                    <SPLIT distance="150" swimtime="00:02:54.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="104" reactiontime="+63" swimtime="00:03:56.44" resultid="19816" heatid="24369" lane="1" entrytime="00:04:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.15" />
                    <SPLIT distance="150" swimtime="00:02:55.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="110" reactiontime="+75" swimtime="00:08:27.57" resultid="19817" heatid="24430" lane="5" entrytime="00:08:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:50.53" />
                    <SPLIT distance="200" swimtime="00:04:08.01" />
                    <SPLIT distance="300" swimtime="00:06:21.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="101" reactiontime="+61" swimtime="00:01:46.75" resultid="19818" heatid="24438" lane="1" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-02-01" firstname="Ewa" gender="F" lastname="Łukasiuk" nation="POL" athleteid="20954">
              <RESULTS>
                <RESULT eventid="1062" points="371" reactiontime="+76" swimtime="00:00:32.92" resultid="20955" heatid="24279" lane="6" entrytime="00:00:32.90" />
                <RESULT eventid="1256" points="306" reactiontime="+44" swimtime="00:01:16.68" resultid="20956" heatid="24351" lane="1" entrytime="00:01:16.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="337" reactiontime="+42" swimtime="00:00:42.22" resultid="20957" heatid="24457" lane="2" entrytime="00:00:42.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-16" firstname="Wojciech" gender="M" lastname="Żmiejko" nation="POL" athleteid="20274">
              <RESULTS>
                <RESULT eventid="1079" points="390" reactiontime="+81" swimtime="00:00:28.61" resultid="20275" heatid="24291" lane="3" entrytime="00:00:28.95" />
                <RESULT eventid="1113" points="334" reactiontime="+83" swimtime="00:02:44.25" resultid="20276" heatid="24305" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.20" />
                    <SPLIT distance="100" swimtime="00:01:17.87" />
                    <SPLIT distance="150" swimtime="00:02:06.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="293" swimtime="00:00:36.10" resultid="20277" heatid="24333" lane="3" entrytime="00:00:35.95" />
                <RESULT eventid="1273" points="363" swimtime="00:01:05.73" resultid="20278" heatid="24361" lane="0" entrytime="00:01:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="372" swimtime="00:00:30.94" resultid="20279" heatid="24395" lane="1" entrytime="00:00:30.95" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="20280" heatid="24406" lane="6" entrytime="00:01:18.95" />
                <RESULT eventid="1613" points="326" swimtime="00:01:12.37" resultid="20281" heatid="24440" lane="2" entrytime="00:01:12.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="338" swimtime="00:00:37.23" resultid="20282" heatid="24463" lane="6" entrytime="00:00:37.95" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="356" reactiontime="+65" swimtime="00:02:11.74" resultid="22687" heatid="24374" lane="9" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                    <SPLIT distance="100" swimtime="00:01:09.72" />
                    <SPLIT distance="150" swimtime="00:01:40.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22678" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="22657" number="2" />
                    <RELAYPOSITION athleteid="23087" number="3" reactiontime="+2" />
                    <RELAYPOSITION athleteid="22641" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="397" swimtime="00:01:55.36" resultid="22688" heatid="24427" lane="8" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.32" />
                    <SPLIT distance="100" swimtime="00:00:55.36" />
                    <SPLIT distance="150" swimtime="00:01:24.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22657" number="1" />
                    <RELAYPOSITION athleteid="22678" number="2" />
                    <RELAYPOSITION athleteid="23087" number="3" reactiontime="+19" />
                    <RELAYPOSITION athleteid="22641" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="20742" name="Niezrzeszone JK TEAM">
          <CONTACT email="joanna.kwatera@gmail.com" name="Joanna Kwatera" phone="790611187" />
          <ATHLETES>
            <ATHLETE birthdate="1998-09-13" firstname="Karolina" gender="F" lastname="Dudziak" nation="POL" athleteid="20758">
              <RESULTS>
                <RESULT eventid="1147" reactiontime="+111" status="OTL" swimtime="00:13:11.57" resultid="20759" heatid="24312" lane="0" entrytime="00:11:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.75" />
                    <SPLIT distance="100" swimtime="00:01:27.76" />
                    <SPLIT distance="150" swimtime="00:02:14.68" />
                    <SPLIT distance="200" swimtime="00:03:03.32" />
                    <SPLIT distance="250" swimtime="00:03:52.98" />
                    <SPLIT distance="300" swimtime="00:04:42.78" />
                    <SPLIT distance="350" swimtime="00:05:33.49" />
                    <SPLIT distance="400" swimtime="00:06:24.23" />
                    <SPLIT distance="450" swimtime="00:07:15.87" />
                    <SPLIT distance="500" swimtime="00:08:07.67" />
                    <SPLIT distance="550" swimtime="00:08:59.06" />
                    <SPLIT distance="600" swimtime="00:09:50.42" />
                    <SPLIT distance="650" swimtime="00:10:41.84" />
                    <SPLIT distance="700" swimtime="00:11:32.96" />
                    <SPLIT distance="750" swimtime="00:12:23.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="243" reactiontime="+77" swimtime="00:01:22.77" resultid="20760" heatid="24350" lane="2" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="246" reactiontime="+82" swimtime="00:03:00.14" resultid="20761" heatid="24412" lane="2" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.16" />
                    <SPLIT distance="100" swimtime="00:01:27.40" />
                    <SPLIT distance="150" swimtime="00:02:14.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="239" reactiontime="+65" swimtime="00:06:20.71" resultid="20762" heatid="24472" lane="9" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.89" />
                    <SPLIT distance="100" swimtime="00:01:27.28" />
                    <SPLIT distance="150" swimtime="00:02:14.72" />
                    <SPLIT distance="200" swimtime="00:03:04.08" />
                    <SPLIT distance="250" swimtime="00:03:53.54" />
                    <SPLIT distance="300" swimtime="00:04:43.85" />
                    <SPLIT distance="350" swimtime="00:05:33.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-09-12" firstname="Joanna" gender="F" lastname="Kwatera" nation="POL" athleteid="20747">
              <RESULTS>
                <RESULT eventid="1222" points="320" reactiontime="+71" swimtime="00:03:23.32" resultid="20748" heatid="24339" lane="4" entrytime="00:03:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.54" />
                    <SPLIT distance="100" swimtime="00:01:39.44" />
                    <SPLIT distance="150" swimtime="00:02:31.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-05-27" firstname="Ada" gender="F" lastname="Malinowska" nation="POL" athleteid="20743">
              <RESULTS>
                <RESULT eventid="1256" points="463" swimtime="00:01:06.80" resultid="20744" heatid="24352" lane="5" entrytime="00:01:08.00" />
                <RESULT eventid="1388" points="376" swimtime="00:01:28.85" resultid="20745" heatid="24378" lane="7" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="447" swimtime="00:00:31.95" resultid="20746" heatid="24388" lane="6" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-04-04" firstname="Karolina" gender="F" lastname="Szkudlarek" nation="POL" athleteid="20749">
              <RESULTS>
                <RESULT eventid="1062" points="521" reactiontime="+82" swimtime="00:00:29.40" resultid="20750" heatid="24281" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="1147" points="409" reactiontime="+77" swimtime="00:10:52.58" resultid="20751" heatid="24312" lane="3" entrytime="00:10:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                    <SPLIT distance="100" swimtime="00:01:10.28" />
                    <SPLIT distance="150" swimtime="00:01:49.40" />
                    <SPLIT distance="200" swimtime="00:02:29.20" />
                    <SPLIT distance="250" swimtime="00:03:09.57" />
                    <SPLIT distance="300" swimtime="00:03:50.34" />
                    <SPLIT distance="350" swimtime="00:04:30.92" />
                    <SPLIT distance="400" swimtime="00:05:13.16" />
                    <SPLIT distance="450" swimtime="00:05:55.28" />
                    <SPLIT distance="500" swimtime="00:06:37.17" />
                    <SPLIT distance="550" swimtime="00:07:19.69" />
                    <SPLIT distance="600" swimtime="00:08:02.12" />
                    <SPLIT distance="650" swimtime="00:08:45.61" />
                    <SPLIT distance="700" swimtime="00:09:28.32" />
                    <SPLIT distance="750" swimtime="00:10:11.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="458" swimtime="00:00:35.10" resultid="20752" heatid="24327" lane="7" entrytime="00:00:34.00" />
                <RESULT eventid="1256" points="520" reactiontime="+71" swimtime="00:01:04.30" resultid="20753" heatid="24353" lane="6" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="448" reactiontime="+62" swimtime="00:01:15.79" resultid="20754" heatid="24402" lane="8" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="493" reactiontime="+71" swimtime="00:02:22.99" resultid="20755" heatid="24414" lane="6" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                    <SPLIT distance="100" swimtime="00:01:08.27" />
                    <SPLIT distance="150" swimtime="00:01:45.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="443" reactiontime="+71" swimtime="00:00:38.56" resultid="20756" heatid="24458" lane="6" entrytime="00:00:37.00" />
                <RESULT eventid="1721" points="449" reactiontime="+75" swimtime="00:05:08.60" resultid="20757" heatid="24473" lane="5" entrytime="00:04:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                    <SPLIT distance="100" swimtime="00:01:11.96" />
                    <SPLIT distance="150" swimtime="00:01:50.74" />
                    <SPLIT distance="200" swimtime="00:02:30.02" />
                    <SPLIT distance="250" swimtime="00:03:10.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-02-17" firstname="Nadia" gender="F" lastname="Świętek" nation="POL" athleteid="20763">
              <RESULTS>
                <RESULT eventid="1062" points="248" reactiontime="+107" swimtime="00:00:37.63" resultid="20764" heatid="24277" lane="1" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="CZE" region="SLPL" clubid="21270" name="Plavecký klub Slávia VŠ Plzeň z.s.">
          <CONTACT city="Plzeň" email="bazilova@plaveckyklubplzen.cz" internet="www.plaveckyklubplzen.cz" name="Radka Bažilová" phone="+420737037564" street="náměstí Generála Píky 42" zip="326 00" />
          <ATHLETES>
            <ATHLETE birthdate="1977-10-18" firstname="Kamila Dagmara" gender="F" lastname="Častoral" nation="CZE" athleteid="21271">
              <RESULTS>
                <RESULT eventid="1222" points="172" reactiontime="+91" swimtime="00:04:09.76" resultid="21272" heatid="24338" lane="2" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.04" />
                    <SPLIT distance="100" swimtime="00:02:03.38" />
                    <SPLIT distance="150" swimtime="00:03:06.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="33" reactiontime="+90" swimtime="00:06:17.90" resultid="21273" heatid="24366" lane="4" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:30.85" />
                    <SPLIT distance="100" swimtime="00:03:11.45" />
                    <SPLIT distance="150" swimtime="00:04:50.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="150" reactiontime="+83" swimtime="00:02:00.64" resultid="21274" heatid="24377" lane="1" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="28" reactiontime="+82" swimtime="00:03:01.63" resultid="21275" heatid="24435" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="152" reactiontime="+72" swimtime="00:00:55.08" resultid="21276" heatid="24455" lane="5" entrytime="00:00:55.00" />
                <RESULT eventid="1555" points="96" reactiontime="+98" swimtime="00:09:40.60" resultid="23435" heatid="24428" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.97" />
                    <SPLIT distance="150" swimtime="00:04:11.07" />
                    <SPLIT distance="200" swimtime="00:07:34.50" />
                    <SPLIT distance="250" swimtime="00:06:29.61" />
                    <SPLIT distance="350" swimtime="00:08:37.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="CZE" clubid="19955" name="Plavecký klub Zábřeh">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1973-06-01" firstname="Petr" gender="M" lastname="Horvat" nation="CZE" athleteid="19971">
              <RESULTS>
                <RESULT eventid="1079" points="292" reactiontime="+89" swimtime="00:00:31.49" resultid="19972" heatid="24289" lane="6" entrytime="00:00:30.73" />
                <RESULT eventid="14189" points="247" reactiontime="+84" swimtime="00:11:59.70" resultid="19973" heatid="24315" lane="5" entrytime="00:12:06.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.14" />
                    <SPLIT distance="100" swimtime="00:02:54.74" />
                    <SPLIT distance="150" swimtime="00:02:15.71" />
                    <SPLIT distance="250" swimtime="00:03:39.88" />
                    <SPLIT distance="300" swimtime="00:05:57.05" />
                    <SPLIT distance="350" swimtime="00:05:11.25" />
                    <SPLIT distance="400" swimtime="00:07:28.65" />
                    <SPLIT distance="450" swimtime="00:06:43.23" />
                    <SPLIT distance="550" swimtime="00:08:14.20" />
                    <SPLIT distance="650" swimtime="00:09:45.79" />
                    <SPLIT distance="750" swimtime="00:11:16.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="322" reactiontime="+79" swimtime="00:03:04.65" resultid="19974" heatid="24344" lane="4" entrytime="00:03:05.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.06" />
                    <SPLIT distance="100" swimtime="00:01:29.45" />
                    <SPLIT distance="150" swimtime="00:02:17.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="283" reactiontime="+43" swimtime="00:01:11.42" resultid="19975" heatid="24358" lane="2" entrytime="00:01:10.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="258" swimtime="00:00:34.94" resultid="19976" heatid="24393" lane="9" entrytime="00:00:35.71" />
                <RESULT eventid="1508" points="238" reactiontime="+68" swimtime="00:02:44.55" resultid="19977" heatid="24419" lane="7" entrytime="00:02:45.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.71" />
                    <SPLIT distance="100" swimtime="00:01:20.90" />
                    <SPLIT distance="150" swimtime="00:02:04.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="284" swimtime="00:00:39.46" resultid="19978" heatid="24463" lane="8" entrytime="00:00:38.59" />
                <RESULT eventid="1744" points="241" reactiontime="+78" swimtime="00:05:53.24" resultid="19979" heatid="24478" lane="3" entrytime="00:05:54.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.22" />
                    <SPLIT distance="100" swimtime="00:01:24.94" />
                    <SPLIT distance="150" swimtime="00:02:10.02" />
                    <SPLIT distance="200" swimtime="00:02:55.69" />
                    <SPLIT distance="250" swimtime="00:03:40.85" />
                    <SPLIT distance="300" swimtime="00:04:26.03" />
                    <SPLIT distance="350" swimtime="00:05:11.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-09-19" firstname="Jiri" gender="M" lastname="Sip" nation="CZE" athleteid="19963">
              <RESULTS>
                <RESULT eventid="1079" points="425" reactiontime="+92" swimtime="00:00:27.79" resultid="19964" heatid="24293" lane="8" entrytime="00:00:27.64" />
                <RESULT eventid="1113" points="395" reactiontime="+104" swimtime="00:02:35.33" resultid="19965" heatid="24306" lane="0" entrytime="00:02:34.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                    <SPLIT distance="100" swimtime="00:01:14.26" />
                    <SPLIT distance="150" swimtime="00:02:00.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="387" swimtime="00:00:32.93" resultid="19966" heatid="24334" lane="6" entrytime="00:00:32.79" />
                <RESULT eventid="1273" points="464" reactiontime="+81" swimtime="00:01:00.56" resultid="19967" heatid="24362" lane="7" entrytime="00:01:00.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="387" reactiontime="+144" swimtime="00:01:11.09" resultid="19968" heatid="24407" lane="6" entrytime="00:01:11.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="385" reactiontime="+90" swimtime="00:05:35.08" resultid="19969" heatid="24432" lane="4" entrytime="00:05:39.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                    <SPLIT distance="100" swimtime="00:01:14.13" />
                    <SPLIT distance="150" swimtime="00:01:58.78" />
                    <SPLIT distance="200" swimtime="00:02:42.41" />
                    <SPLIT distance="250" swimtime="00:03:31.16" />
                    <SPLIT distance="300" swimtime="00:04:19.31" />
                    <SPLIT distance="350" swimtime="00:04:59.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="351" reactiontime="+84" swimtime="00:02:38.54" resultid="19970" heatid="24451" lane="1" entrytime="00:02:37.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.21" />
                    <SPLIT distance="100" swimtime="00:01:16.77" />
                    <SPLIT distance="150" swimtime="00:01:58.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="GER" clubid="19844" name="Post SV Leipzig">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1985-01-01" firstname="Sven" gender="M" lastname="Lützkendorf" nation="GER" athleteid="19845">
              <RESULTS>
                <RESULT eventid="14207" points="481" reactiontime="+104" swimtime="00:18:31.01" resultid="19846" heatid="24322" lane="3" entrytime="00:18:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                    <SPLIT distance="100" swimtime="00:01:06.46" />
                    <SPLIT distance="150" swimtime="00:01:42.10" />
                    <SPLIT distance="200" swimtime="00:02:18.20" />
                    <SPLIT distance="250" swimtime="00:02:54.66" />
                    <SPLIT distance="300" swimtime="00:03:30.91" />
                    <SPLIT distance="350" swimtime="00:04:07.63" />
                    <SPLIT distance="400" swimtime="00:04:43.83" />
                    <SPLIT distance="450" swimtime="00:05:20.46" />
                    <SPLIT distance="500" swimtime="00:05:57.18" />
                    <SPLIT distance="550" swimtime="00:06:34.15" />
                    <SPLIT distance="600" swimtime="00:07:11.19" />
                    <SPLIT distance="650" swimtime="00:07:48.75" />
                    <SPLIT distance="700" swimtime="00:08:26.22" />
                    <SPLIT distance="750" swimtime="00:09:03.85" />
                    <SPLIT distance="800" swimtime="00:09:41.51" />
                    <SPLIT distance="850" swimtime="00:10:19.36" />
                    <SPLIT distance="900" swimtime="00:10:57.14" />
                    <SPLIT distance="950" swimtime="00:11:35.00" />
                    <SPLIT distance="1000" swimtime="00:12:12.40" />
                    <SPLIT distance="1050" swimtime="00:12:50.52" />
                    <SPLIT distance="1100" swimtime="00:13:27.95" />
                    <SPLIT distance="1150" swimtime="00:14:06.07" />
                    <SPLIT distance="1200" swimtime="00:14:43.74" />
                    <SPLIT distance="1250" swimtime="00:15:21.96" />
                    <SPLIT distance="1300" swimtime="00:15:59.49" />
                    <SPLIT distance="1350" swimtime="00:16:37.57" />
                    <SPLIT distance="1400" swimtime="00:17:15.69" />
                    <SPLIT distance="1450" swimtime="00:17:54.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="463" reactiontime="+66" swimtime="00:00:31.01" resultid="19847" heatid="24335" lane="9" entrytime="00:00:31.70" />
                <RESULT eventid="1273" points="468" reactiontime="+59" swimtime="00:01:00.41" resultid="19848" heatid="24364" lane="9" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="495" reactiontime="+74" swimtime="00:02:08.90" resultid="19849" heatid="24424" lane="6" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.63" />
                    <SPLIT distance="100" swimtime="00:01:02.03" />
                    <SPLIT distance="150" swimtime="00:01:35.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="460" reactiontime="+96" swimtime="00:05:15.84" resultid="19850" heatid="24433" lane="7" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="100" swimtime="00:01:09.51" />
                    <SPLIT distance="150" swimtime="00:01:50.41" />
                    <SPLIT distance="200" swimtime="00:02:31.26" />
                    <SPLIT distance="250" swimtime="00:03:16.40" />
                    <SPLIT distance="300" swimtime="00:04:01.79" />
                    <SPLIT distance="350" swimtime="00:04:39.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="SLA" clubid="20163" name="RMKS Rybnik">
          <CONTACT email="aniaduda0511@tlen.pl" name="Duda Anna" phone="792666159" />
          <ATHLETES>
            <ATHLETE birthdate="1981-04-15" firstname="Anna" gender="F" lastname="Duda" nation="POL" athleteid="20164">
              <RESULTS>
                <RESULT eventid="1062" status="DNS" swimtime="00:00:00.00" resultid="20165" heatid="24281" lane="3" entrytime="00:00:28.20" />
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="20166" heatid="24327" lane="0" entrytime="00:00:36.00" />
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="20167" heatid="24353" lane="2" entrytime="00:01:04.30" />
                <RESULT eventid="1423" status="DNS" swimtime="00:00:00.00" resultid="20168" heatid="24389" lane="4" entrytime="00:00:29.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ROYAL" nation="SVK" region="BAO" clubid="20209" name="ROYAL plavecký klub">
          <CONTACT city="Bratislava" email="schild@royalclub.sk" name="Schild Igor" phone="0911175865" street="Iľjušinová 6" zip="85101" />
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="20107" name="Rydułtowska Akademia Aktywnego Seniora">
          <CONTACT name="MARIAN" street="OTLIK" />
          <ATHLETES>
            <ATHLETE birthdate="1940-05-16" firstname="Rudolf" gender="M" lastname="Bugla" nation="POL" athleteid="20148">
              <RESULTS>
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="20149" heatid="24301" lane="6" entrytime="00:04:40.00" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="20150" heatid="24329" lane="7" entrytime="00:00:59.00" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="20151" heatid="24342" lane="7" entrytime="00:04:30.12" />
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="20152" heatid="24380" lane="5" entrytime="00:02:20.14" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="20153" heatid="24430" lane="2" entrytime="00:09:50.20" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="20154" heatid="24437" lane="2" entrytime="00:02:40.05" />
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="20155" heatid="24447" lane="8" entrytime="00:04:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-11-24" firstname="Jerzy" gender="M" lastname="Ciecior" nation="POL" athleteid="20139">
              <RESULTS>
                <RESULT eventid="1113" points="161" reactiontime="+87" swimtime="00:03:29.23" resultid="20140" heatid="24303" lane="0" entrytime="00:03:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.37" />
                    <SPLIT distance="100" swimtime="00:01:38.77" />
                    <SPLIT distance="150" swimtime="00:02:42.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14207" points="166" reactiontime="+96" swimtime="00:26:23.44" resultid="20141" heatid="24321" lane="1" entrytime="00:25:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.49" />
                    <SPLIT distance="100" swimtime="00:01:36.77" />
                    <SPLIT distance="150" swimtime="00:02:28.76" />
                    <SPLIT distance="200" swimtime="00:03:21.38" />
                    <SPLIT distance="250" swimtime="00:04:14.98" />
                    <SPLIT distance="300" swimtime="00:05:07.61" />
                    <SPLIT distance="350" swimtime="00:06:00.89" />
                    <SPLIT distance="400" swimtime="00:06:53.43" />
                    <SPLIT distance="450" swimtime="00:07:47.02" />
                    <SPLIT distance="500" swimtime="00:08:39.34" />
                    <SPLIT distance="550" swimtime="00:09:32.62" />
                    <SPLIT distance="600" swimtime="00:10:25.38" />
                    <SPLIT distance="650" swimtime="00:11:18.77" />
                    <SPLIT distance="700" swimtime="00:12:11.78" />
                    <SPLIT distance="750" swimtime="00:13:05.20" />
                    <SPLIT distance="800" swimtime="00:13:57.55" />
                    <SPLIT distance="850" swimtime="00:14:51.22" />
                    <SPLIT distance="900" swimtime="00:15:44.03" />
                    <SPLIT distance="950" swimtime="00:16:38.42" />
                    <SPLIT distance="1000" swimtime="00:17:30.93" />
                    <SPLIT distance="1050" swimtime="00:18:24.75" />
                    <SPLIT distance="1100" swimtime="00:19:18.06" />
                    <SPLIT distance="1150" swimtime="00:20:12.15" />
                    <SPLIT distance="1200" swimtime="00:21:05.78" />
                    <SPLIT distance="1250" swimtime="00:21:59.04" />
                    <SPLIT distance="1300" swimtime="00:22:52.79" />
                    <SPLIT distance="1350" swimtime="00:23:46.75" />
                    <SPLIT distance="1400" swimtime="00:24:39.55" />
                    <SPLIT distance="1450" swimtime="00:25:32.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="190" swimtime="00:00:41.69" resultid="20142" heatid="24331" lane="5" entrytime="00:00:41.00" />
                <RESULT eventid="1341" points="92" reactiontime="+68" swimtime="00:04:06.14" resultid="20143" heatid="24369" lane="2" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.99" />
                    <SPLIT distance="100" swimtime="00:01:56.38" />
                    <SPLIT distance="150" swimtime="00:03:03.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="145" reactiontime="+92" swimtime="00:01:38.50" resultid="20144" heatid="24405" lane="0" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="146" reactiontime="+80" swimtime="00:07:42.74" resultid="20145" heatid="24431" lane="2" entrytime="00:07:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.61" />
                    <SPLIT distance="100" swimtime="00:01:58.14" />
                    <SPLIT distance="150" swimtime="00:02:55.42" />
                    <SPLIT distance="200" swimtime="00:03:52.34" />
                    <SPLIT distance="250" swimtime="00:04:58.43" />
                    <SPLIT distance="300" swimtime="00:06:02.55" />
                    <SPLIT distance="350" swimtime="00:06:53.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="131" reactiontime="+66" swimtime="00:01:38.01" resultid="20146" heatid="24439" lane="7" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="155" reactiontime="+77" swimtime="00:03:27.94" resultid="20147" heatid="24448" lane="4" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.22" />
                    <SPLIT distance="100" swimtime="00:01:42.34" />
                    <SPLIT distance="150" swimtime="00:02:36.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-02-02" firstname="Maria" gender="F" lastname="Lippa" nation="POL" athleteid="20115">
              <RESULTS>
                <RESULT eventid="1062" points="20" swimtime="00:01:26.74" resultid="20116" heatid="24276" lane="8" />
                <RESULT eventid="1187" points="27" swimtime="00:01:29.25" resultid="20117" heatid="24323" lane="6" />
                <RESULT eventid="1256" points="29" swimtime="00:02:46.59" resultid="20118" heatid="24348" lane="7" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="28" reactiontime="+192" swimtime="00:03:10.02" resultid="20119" heatid="24399" lane="4" entrytime="00:03:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:30.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="32" swimtime="00:05:52.29" resultid="20120" heatid="24410" lane="0" entrytime="00:05:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.71" />
                    <SPLIT distance="100" swimtime="00:02:52.38" />
                    <SPLIT distance="150" swimtime="00:04:22.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="31" reactiontime="+180" swimtime="00:06:32.75" resultid="20121" heatid="24443" lane="7" entrytime="00:06:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:31.73" />
                    <SPLIT distance="100" swimtime="00:03:12.16" />
                    <SPLIT distance="150" swimtime="00:04:55.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="23" swimtime="00:01:43.12" resultid="20122" heatid="24454" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-08-21" firstname="Kądzioła" gender="M" lastname="Michał" nation="POL" athleteid="20108">
              <RESULTS>
                <RESULT eventid="1079" points="326" reactiontime="+79" swimtime="00:00:30.36" resultid="20109" heatid="24292" lane="9" entrytime="00:00:28.50" />
                <RESULT eventid="1205" points="320" reactiontime="+74" swimtime="00:00:35.06" resultid="20110" heatid="24334" lane="7" entrytime="00:00:33.20" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="20111" heatid="24361" lane="7" entrytime="00:01:04.00" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="20112" heatid="24395" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="20113" heatid="24407" lane="8" entrytime="00:01:14.00" />
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="20114" heatid="24450" lane="5" entrytime="00:02:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1945-12-07" firstname="Miron" gender="M" lastname="Starosta" nation="POL" athleteid="20130">
              <RESULTS>
                <RESULT eventid="1079" points="74" reactiontime="+91" swimtime="00:00:49.79" resultid="20131" heatid="24283" lane="4" entrytime="00:00:48.00" />
                <RESULT eventid="1113" points="60" reactiontime="+118" swimtime="00:04:50.61" resultid="20132" heatid="24301" lane="1" entrytime="00:04:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.85" />
                    <SPLIT distance="100" swimtime="00:02:19.22" />
                    <SPLIT distance="150" swimtime="00:03:43.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="61" reactiontime="+84" swimtime="00:05:21.07" resultid="20133" heatid="24342" lane="9" entrytime="00:05:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.36" />
                    <SPLIT distance="100" swimtime="00:02:38.14" />
                    <SPLIT distance="150" swimtime="00:04:01.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" status="DNS" swimtime="00:00:00.00" resultid="20134" heatid="24368" lane="2" />
                <RESULT eventid="1406" points="67" reactiontime="+41" swimtime="00:02:20.07" resultid="20135" heatid="24381" lane="9" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="20136" heatid="24430" lane="9" />
                <RESULT eventid="1613" points="27" reactiontime="+77" swimtime="00:02:45.34" resultid="20137" heatid="24437" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="76" reactiontime="+74" swimtime="00:01:01.03" resultid="20138" heatid="24460" lane="1" entrytime="00:01:02.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-05-26" firstname="Władysław" gender="M" lastname="Szurek" nation="POL" athleteid="20123">
              <RESULTS>
                <RESULT eventid="1205" points="11" swimtime="00:01:46.38" resultid="20124" heatid="24328" lane="6" />
                <RESULT eventid="1273" points="19" reactiontime="+94" swimtime="00:02:53.07" resultid="20125" heatid="24354" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:22.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="11" reactiontime="+103" swimtime="00:03:51.96" resultid="20126" heatid="24403" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:47.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="22" reactiontime="+91" swimtime="00:06:01.29" resultid="20127" heatid="24415" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.92" />
                    <SPLIT distance="150" swimtime="00:04:28.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="12" swimtime="00:08:08.65" resultid="20128" heatid="24446" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:46.71" />
                    <SPLIT distance="150" swimtime="00:05:59.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="20129" heatid="24474" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="22689" name="Sekcja Masters UKP Jedynka Elbląg">
          <CONTACT name="a" />
          <ATHLETES>
            <ATHLETE birthdate="1954-02-04" firstname="Ewa" gender="F" lastname="Kerner Mateusiak" nation="POL" athleteid="22690">
              <RESULTS>
                <RESULT eventid="1062" points="48" swimtime="00:01:04.91" resultid="22691" heatid="24276" lane="2" entrytime="00:01:00.00" />
                <RESULT eventid="1147" points="63" swimtime="00:20:15.12" resultid="22692" heatid="24310" lane="7" entrytime="00:20:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.26" />
                    <SPLIT distance="100" swimtime="00:02:21.20" />
                    <SPLIT distance="150" swimtime="00:03:39.53" />
                    <SPLIT distance="200" swimtime="00:04:56.28" />
                    <SPLIT distance="250" swimtime="00:06:13.37" />
                    <SPLIT distance="300" swimtime="00:07:29.41" />
                    <SPLIT distance="350" swimtime="00:08:45.40" />
                    <SPLIT distance="400" swimtime="00:10:03.00" />
                    <SPLIT distance="450" swimtime="00:11:18.85" />
                    <SPLIT distance="500" swimtime="00:12:35.59" />
                    <SPLIT distance="550" swimtime="00:13:51.52" />
                    <SPLIT distance="600" swimtime="00:15:08.99" />
                    <SPLIT distance="650" swimtime="00:16:25.65" />
                    <SPLIT distance="700" swimtime="00:17:42.79" />
                    <SPLIT distance="750" swimtime="00:18:59.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="55" swimtime="00:01:11.14" resultid="22693" heatid="24323" lane="4" entrytime="00:01:09.35" />
                <RESULT eventid="1256" points="50" swimtime="00:02:19.98" resultid="22694" heatid="24348" lane="5" entrytime="00:01:58.00" />
                <RESULT eventid="1457" points="45" swimtime="00:02:42.13" resultid="22695" heatid="24400" lane="8" entrytime="00:02:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="55" swimtime="00:04:55.45" resultid="22696" heatid="24410" lane="6" entrytime="00:04:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" status="DNF" swimtime="00:00:00.00" resultid="22697" heatid="24470" lane="0" entrytime="00:10:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.47" />
                    <SPLIT distance="100" swimtime="00:02:19.43" />
                    <SPLIT distance="150" swimtime="00:03:34.60" />
                    <SPLIT distance="300" swimtime="00:07:20.38" />
                    <SPLIT distance="350" swimtime="00:08:34.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="20737" name="Siemacha Kraków">
          <CONTACT email="joanna.kwatera@gmail.com" name="Joanna Kwatera" phone="790611187" />
          <ATHLETES>
            <ATHLETE birthdate="1980-02-23" firstname="Monika" gender="F" lastname="Kuc" nation="POL" athleteid="20738">
              <RESULTS>
                <RESULT eventid="1147" points="229" reactiontime="+105" swimtime="00:13:11.56" resultid="20739" heatid="24311" lane="7" entrytime="00:13:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.81" />
                    <SPLIT distance="100" swimtime="00:01:31.01" />
                    <SPLIT distance="150" swimtime="00:02:20.10" />
                    <SPLIT distance="200" swimtime="00:03:10.09" />
                    <SPLIT distance="250" swimtime="00:04:00.25" />
                    <SPLIT distance="300" swimtime="00:04:51.27" />
                    <SPLIT distance="350" swimtime="00:05:42.06" />
                    <SPLIT distance="400" swimtime="00:06:32.89" />
                    <SPLIT distance="450" swimtime="00:07:23.53" />
                    <SPLIT distance="500" swimtime="00:08:14.09" />
                    <SPLIT distance="550" swimtime="00:09:04.76" />
                    <SPLIT distance="600" swimtime="00:09:55.30" />
                    <SPLIT distance="650" swimtime="00:10:44.95" />
                    <SPLIT distance="700" swimtime="00:11:35.44" />
                    <SPLIT distance="750" swimtime="00:12:25.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-08" firstname="Karolina" gender="F" lastname="Spóła" nation="POL" athleteid="20740">
              <RESULTS>
                <RESULT eventid="1062" points="137" reactiontime="+92" swimtime="00:00:45.86" resultid="20741" heatid="24276" lane="6" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="21603" name="SIKRET Gliwice">
          <CONTACT city="Gliwice" email="joannaeco@tlen.pl" name="Joanna Zagała" phone="601427257" state="ŚLĄSK" street="Kościuszki 35" zip="44-100" />
          <ATHLETES>
            <ATHLETE birthdate="1958-02-05" firstname="Zofia" gender="F" lastname="Dąbrowska" nation="POL" athleteid="21613">
              <RESULTS>
                <RESULT eventid="1062" points="131" reactiontime="+86" swimtime="00:00:46.58" resultid="21614" heatid="24277" lane="0" entrytime="00:00:44.00" />
                <RESULT eventid="1147" points="116" reactiontime="+89" swimtime="00:16:32.36" resultid="21615" heatid="24310" lane="4" entrytime="00:16:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.31" />
                    <SPLIT distance="100" swimtime="00:01:51.00" />
                    <SPLIT distance="150" swimtime="00:02:52.25" />
                    <SPLIT distance="200" swimtime="00:03:53.80" />
                    <SPLIT distance="250" swimtime="00:04:55.54" />
                    <SPLIT distance="350" swimtime="00:06:59.84" />
                    <SPLIT distance="400" swimtime="00:08:02.53" />
                    <SPLIT distance="450" swimtime="00:09:05.44" />
                    <SPLIT distance="500" swimtime="00:10:09.24" />
                    <SPLIT distance="550" swimtime="00:11:11.08" />
                    <SPLIT distance="600" swimtime="00:12:14.36" />
                    <SPLIT distance="650" swimtime="00:13:19.09" />
                    <SPLIT distance="700" swimtime="00:14:24.97" />
                    <SPLIT distance="750" swimtime="00:15:31.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="130" reactiontime="+66" swimtime="00:04:34.06" resultid="21616" heatid="24338" lane="3" entrytime="00:04:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.83" />
                    <SPLIT distance="100" swimtime="00:02:12.78" />
                    <SPLIT distance="150" swimtime="00:03:22.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="128" reactiontime="+42" swimtime="00:02:07.22" resultid="21617" heatid="24377" lane="0" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="120" reactiontime="+56" swimtime="00:03:48.91" resultid="21618" heatid="24411" lane="9" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:53.20" />
                    <SPLIT distance="100" swimtime="00:01:51.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="62" reactiontime="+98" swimtime="00:02:19.90" resultid="21619" heatid="24434" lane="4" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="166" reactiontime="+81" swimtime="00:00:53.48" resultid="21620" heatid="24455" lane="4" entrytime="00:00:53.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-04-20" firstname="Wojciech" gender="M" lastname="Kosiak" nation="POL" athleteid="21635">
              <RESULTS>
                <RESULT eventid="1079" points="137" reactiontime="+119" swimtime="00:00:40.53" resultid="21636" heatid="24284" lane="7" entrytime="00:00:42.00" />
                <RESULT eventid="1273" points="123" reactiontime="+98" swimtime="00:01:34.17" resultid="21637" heatid="24355" lane="6" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="58" reactiontime="+92" swimtime="00:00:57.38" resultid="21638" heatid="24390" lane="6" entrytime="00:00:56.00" />
                <RESULT eventid="1508" points="97" reactiontime="+90" swimtime="00:03:41.29" resultid="21639" heatid="24416" lane="5" entrytime="00:03:46.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:49.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-16" firstname="Stanisław" gender="M" lastname="Twardysko" nation="POL" athleteid="21621">
              <RESULTS>
                <RESULT eventid="1079" points="209" reactiontime="+91" swimtime="00:00:35.23" resultid="21622" heatid="24285" lane="5" entrytime="00:00:36.53" />
                <RESULT eventid="1205" points="177" swimtime="00:00:42.72" resultid="21623" heatid="24331" lane="7" entrytime="00:00:43.70" />
                <RESULT eventid="1273" points="198" reactiontime="+62" swimtime="00:01:20.38" resultid="21624" heatid="24356" lane="3" entrytime="00:01:23.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="129" reactiontime="+64" swimtime="00:00:43.97" resultid="21625" heatid="24390" lane="5" entrytime="00:00:55.00" />
                <RESULT eventid="1508" points="169" reactiontime="+95" swimtime="00:03:04.28" resultid="21626" heatid="24418" lane="2" entrytime="00:03:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.42" />
                    <SPLIT distance="100" swimtime="00:01:27.91" />
                    <SPLIT distance="150" swimtime="00:02:17.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="172" reactiontime="+55" swimtime="00:06:35.05" resultid="21627" heatid="24477" lane="9" entrytime="00:06:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.91" />
                    <SPLIT distance="100" swimtime="00:01:30.62" />
                    <SPLIT distance="150" swimtime="00:04:04.91" />
                    <SPLIT distance="200" swimtime="00:03:12.78" />
                    <SPLIT distance="250" swimtime="00:05:47.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-06-24" firstname="Joanna" gender="F" lastname="Zagała" nation="POL" athleteid="21604">
              <RESULTS>
                <RESULT eventid="1062" points="228" reactiontime="+76" swimtime="00:00:38.74" resultid="21605" heatid="24277" lane="9" entrytime="00:00:44.00" />
                <RESULT eventid="1147" points="175" reactiontime="+95" swimtime="00:14:25.38" resultid="21606" heatid="24310" lane="5" entrytime="00:16:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.76" />
                    <SPLIT distance="100" swimtime="00:01:41.73" />
                    <SPLIT distance="150" swimtime="00:02:36.23" />
                    <SPLIT distance="200" swimtime="00:03:31.55" />
                    <SPLIT distance="250" swimtime="00:04:26.23" />
                    <SPLIT distance="350" swimtime="00:06:15.94" />
                    <SPLIT distance="450" swimtime="00:08:05.56" />
                    <SPLIT distance="550" swimtime="00:09:55.13" />
                    <SPLIT distance="650" swimtime="00:11:45.40" />
                    <SPLIT distance="750" swimtime="00:13:35.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="166" swimtime="00:00:49.20" resultid="21607" heatid="24324" lane="7" entrytime="00:00:59.00" />
                <RESULT eventid="1256" points="210" reactiontime="+76" swimtime="00:01:26.88" resultid="21608" heatid="24349" lane="2" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="147" reactiontime="+82" swimtime="00:02:01.49" resultid="21609" heatid="24377" lane="8" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="182" reactiontime="+45" swimtime="00:03:19.19" resultid="21610" heatid="24411" lane="0" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.74" />
                    <SPLIT distance="100" swimtime="00:01:41.04" />
                    <SPLIT distance="150" swimtime="00:02:32.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="187" reactiontime="+48" swimtime="00:00:51.37" resultid="21611" heatid="24455" lane="2" entrytime="00:01:00.00" />
                <RESULT eventid="1721" points="174" reactiontime="+88" swimtime="00:07:03.35" resultid="21612" heatid="24471" lane="8" entrytime="00:07:11.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.44" />
                    <SPLIT distance="150" swimtime="00:04:25.06" />
                    <SPLIT distance="350" swimtime="00:06:13.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-10-14" firstname="Teresa" gender="F" lastname="Żylińska" nation="POL" athleteid="21628">
              <RESULTS>
                <RESULT eventid="1062" points="95" reactiontime="+109" swimtime="00:00:51.83" resultid="21629" heatid="24276" lane="3" entrytime="00:00:53.00" />
                <RESULT eventid="1187" points="105" swimtime="00:00:57.35" resultid="21630" heatid="24324" lane="0" entrytime="00:01:02.00" />
                <RESULT eventid="1256" points="74" swimtime="00:02:02.96" resultid="21631" heatid="24348" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="84" reactiontime="+67" swimtime="00:02:12.30" resultid="21632" heatid="24400" lane="7" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="80" swimtime="00:04:21.54" resultid="21633" heatid="24410" lane="7" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.21" />
                    <SPLIT distance="100" swimtime="00:02:05.08" />
                    <SPLIT distance="150" swimtime="00:03:14.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="84" swimtime="00:04:42.73" resultid="21634" heatid="24443" lane="6" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.16" />
                    <SPLIT distance="100" swimtime="00:02:16.93" />
                    <SPLIT distance="150" swimtime="00:03:32.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" reactiontime="+80" swimtime="00:02:40.62" resultid="21640" heatid="24308" lane="6" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.81" />
                    <SPLIT distance="100" swimtime="00:01:26.45" />
                    <SPLIT distance="150" swimtime="00:02:01.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21613" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="21635" number="2" />
                    <RELAYPOSITION athleteid="21621" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="21604" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SSO GUB" nation="POL" region="LBS" clubid="22260" name="Sso Gubin">
          <CONTACT city="Poznań" email="jacek.thiem@gmail.com" name="Thiem Jacek" phone="502 499 565" state="LBS" street="Osiedle Dębina 19 m 34" zip="61-450" />
          <ATHLETES>
            <ATHLETE birthdate="1987-02-05" firstname="Paweł" gender="M" lastname="Krupiński" nation="POL" athleteid="22261">
              <RESULTS>
                <RESULT eventid="1113" points="124" reactiontime="+115" swimtime="00:03:48.24" resultid="22262" heatid="24302" lane="3" entrytime="00:03:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.86" />
                    <SPLIT distance="100" swimtime="00:01:53.12" />
                    <SPLIT distance="150" swimtime="00:02:52.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="149" reactiontime="+76" swimtime="00:03:58.75" resultid="22263" heatid="24343" lane="9" entrytime="00:03:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.44" />
                    <SPLIT distance="100" swimtime="00:01:53.57" />
                    <SPLIT distance="150" swimtime="00:02:57.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="133" reactiontime="+86" swimtime="00:00:43.62" resultid="22264" heatid="24391" lane="6" entrytime="00:00:43.00" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="22265" heatid="24461" lane="0" entrytime="00:00:46.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="22873" name="Start Poznań">
          <CONTACT city="Poznań" email="robert.beym@gmail.com" name="Beym Robert" phone="512111513" street="os. Stefana Batorego 8/67" zip="60-687" />
          <ATHLETES>
            <ATHLETE birthdate="1967-05-14" firstname="Piotr" gender="M" lastname="Monczak" nation="POL" athleteid="22874">
              <RESULTS>
                <RESULT eventid="1079" points="434" reactiontime="+83" swimtime="00:00:27.61" resultid="22875" heatid="24293" lane="3" entrytime="00:00:27.00" />
                <RESULT eventid="1113" points="400" reactiontime="+65" swimtime="00:02:34.60" resultid="22876" heatid="24306" lane="7" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                    <SPLIT distance="100" swimtime="00:01:12.94" />
                    <SPLIT distance="150" swimtime="00:01:59.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="485" swimtime="00:00:59.70" resultid="22877" heatid="24363" lane="8" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="22878" heatid="24395" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1508" points="446" swimtime="00:02:13.49" resultid="22879" heatid="24423" lane="3" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                    <SPLIT distance="100" swimtime="00:01:05.51" />
                    <SPLIT distance="150" swimtime="00:01:39.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="444" swimtime="00:04:48.38" resultid="22880" heatid="24481" lane="5" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.37" />
                    <SPLIT distance="100" swimtime="00:01:09.79" />
                    <SPLIT distance="150" swimtime="00:01:46.63" />
                    <SPLIT distance="200" swimtime="00:02:23.63" />
                    <SPLIT distance="250" swimtime="00:02:59.85" />
                    <SPLIT distance="300" swimtime="00:03:36.26" />
                    <SPLIT distance="350" swimtime="00:04:12.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="STEEF" nation="POL" region="DOL" clubid="21513" name="Steef">
          <CONTACT email="ste1@wp.pl" name="Stefan Skrzypek" phone="500388374" state="DOL" street="Edyty Stein 6" zip="50-322" />
          <ATHLETES>
            <ATHLETE birthdate="1957-06-08" firstname="Wiesław" gender="M" lastname="Ciekliński" nation="POL" athleteid="21527">
              <RESULTS>
                <RESULT eventid="14207" points="201" reactiontime="+104" swimtime="00:24:45.13" resultid="21528" heatid="24321" lane="2" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:16.22" />
                    <SPLIT distance="100" swimtime="00:03:06.30" />
                    <SPLIT distance="150" swimtime="00:03:55.44" />
                    <SPLIT distance="200" swimtime="00:04:44.28" />
                    <SPLIT distance="250" swimtime="00:08:52.27" />
                    <SPLIT distance="300" swimtime="00:14:46.27" />
                    <SPLIT distance="350" swimtime="00:10:34.38" />
                    <SPLIT distance="400" swimtime="00:18:07.26" />
                    <SPLIT distance="450" swimtime="00:13:55.10" />
                    <SPLIT distance="550" swimtime="00:18:57.27" />
                    <SPLIT distance="1150" swimtime="00:20:37.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="225" reactiontime="+79" swimtime="00:01:17.05" resultid="21529" heatid="24358" lane="9" entrytime="00:01:13.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="195" reactiontime="+66" swimtime="00:02:55.69" resultid="21530" heatid="24419" lane="8" entrytime="00:02:51.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.36" />
                    <SPLIT distance="150" swimtime="00:02:11.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="206" reactiontime="+69" swimtime="00:06:12.57" resultid="21531" heatid="24478" lane="8" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.86" />
                    <SPLIT distance="150" swimtime="00:02:13.50" />
                    <SPLIT distance="200" swimtime="00:03:03.38" />
                    <SPLIT distance="250" swimtime="00:03:53.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-09-02" firstname="Stefan" gender="M" lastname="Skrzypek" nation="POL" athleteid="21521">
              <RESULTS>
                <RESULT eventid="14207" points="139" reactiontime="+123" swimtime="00:27:58.20" resultid="21522" heatid="24321" lane="0" entrytime="00:26:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.97" />
                    <SPLIT distance="100" swimtime="00:01:40.32" />
                    <SPLIT distance="150" swimtime="00:02:33.20" />
                    <SPLIT distance="200" swimtime="00:03:28.17" />
                    <SPLIT distance="250" swimtime="00:04:22.11" />
                    <SPLIT distance="300" swimtime="00:05:17.27" />
                    <SPLIT distance="350" swimtime="00:06:10.50" />
                    <SPLIT distance="400" swimtime="00:07:05.80" />
                    <SPLIT distance="450" swimtime="00:08:00.80" />
                    <SPLIT distance="500" swimtime="00:08:56.85" />
                    <SPLIT distance="550" swimtime="00:09:51.70" />
                    <SPLIT distance="600" swimtime="00:10:46.89" />
                    <SPLIT distance="650" swimtime="00:11:43.11" />
                    <SPLIT distance="700" swimtime="00:12:40.77" />
                    <SPLIT distance="750" swimtime="00:13:39.48" />
                    <SPLIT distance="800" swimtime="00:14:36.87" />
                    <SPLIT distance="850" swimtime="00:15:35.55" />
                    <SPLIT distance="900" swimtime="00:16:34.29" />
                    <SPLIT distance="950" swimtime="00:17:30.72" />
                    <SPLIT distance="1000" swimtime="00:18:28.75" />
                    <SPLIT distance="1050" swimtime="00:19:24.43" />
                    <SPLIT distance="1100" swimtime="00:20:20.98" />
                    <SPLIT distance="1150" swimtime="00:21:17.68" />
                    <SPLIT distance="1200" swimtime="00:22:16.74" />
                    <SPLIT distance="1250" swimtime="00:23:14.42" />
                    <SPLIT distance="1300" swimtime="00:24:13.15" />
                    <SPLIT distance="1350" swimtime="00:25:11.44" />
                    <SPLIT distance="1400" swimtime="00:26:09.37" />
                    <SPLIT distance="1450" swimtime="00:27:05.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="21523" heatid="24391" lane="3" entrytime="00:00:42.00" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="21524" heatid="24418" lane="7" entrytime="00:03:04.21" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="21525" heatid="24438" lane="5" entrytime="00:01:35.00" />
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="21526" heatid="24478" lane="0" entrytime="00:06:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-03-19" firstname="Ewa" gender="F" lastname="Szała" nation="POL" athleteid="21514">
              <RESULTS>
                <RESULT eventid="1096" points="298" reactiontime="+104" swimtime="00:03:08.73" resultid="21515" heatid="24298" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.80" />
                    <SPLIT distance="100" swimtime="00:01:32.31" />
                    <SPLIT distance="150" swimtime="00:02:25.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="265" reactiontime="+104" swimtime="00:23:52.90" resultid="21516" heatid="24319" lane="8" entrytime="00:25:52.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.16" />
                    <SPLIT distance="100" swimtime="00:01:29.27" />
                    <SPLIT distance="150" swimtime="00:02:17.15" />
                    <SPLIT distance="200" swimtime="00:03:04.71" />
                    <SPLIT distance="250" swimtime="00:03:51.66" />
                    <SPLIT distance="300" swimtime="00:04:38.62" />
                    <SPLIT distance="350" swimtime="00:05:26.64" />
                    <SPLIT distance="400" swimtime="00:06:12.95" />
                    <SPLIT distance="450" swimtime="00:07:00.50" />
                    <SPLIT distance="500" swimtime="00:09:26.67" />
                    <SPLIT distance="550" swimtime="00:08:37.89" />
                    <SPLIT distance="600" swimtime="00:12:39.98" />
                    <SPLIT distance="650" swimtime="00:10:15.28" />
                    <SPLIT distance="700" swimtime="00:14:16.59" />
                    <SPLIT distance="750" swimtime="00:11:52.05" />
                    <SPLIT distance="800" swimtime="00:15:54.24" />
                    <SPLIT distance="850" swimtime="00:13:27.36" />
                    <SPLIT distance="900" swimtime="00:17:29.79" />
                    <SPLIT distance="950" swimtime="00:15:05.65" />
                    <SPLIT distance="1050" swimtime="00:16:41.78" />
                    <SPLIT distance="1150" swimtime="00:18:17.86" />
                    <SPLIT distance="1250" swimtime="00:19:54.52" />
                    <SPLIT distance="1350" swimtime="00:21:29.90" />
                    <SPLIT distance="1450" swimtime="00:23:06.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="299" reactiontime="+85" swimtime="00:01:26.68" resultid="21517" heatid="24401" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="292" reactiontime="+76" swimtime="00:06:41.47" resultid="21518" heatid="24429" lane="7" entrytime="00:07:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.80" />
                    <SPLIT distance="100" swimtime="00:01:37.91" />
                    <SPLIT distance="150" swimtime="00:02:28.23" />
                    <SPLIT distance="200" swimtime="00:03:18.15" />
                    <SPLIT distance="250" swimtime="00:04:14.88" />
                    <SPLIT distance="300" swimtime="00:05:13.02" />
                    <SPLIT distance="350" swimtime="00:05:58.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="288" reactiontime="+89" swimtime="00:03:07.79" resultid="21519" heatid="24444" lane="7" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.53" />
                    <SPLIT distance="100" swimtime="00:01:32.19" />
                    <SPLIT distance="150" swimtime="00:02:19.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="259" reactiontime="+106" swimtime="00:06:10.50" resultid="21520" heatid="24471" lane="4" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.50" />
                    <SPLIT distance="100" swimtime="00:01:29.69" />
                    <SPLIT distance="150" swimtime="00:02:17.12" />
                    <SPLIT distance="200" swimtime="00:03:05.22" />
                    <SPLIT distance="250" swimtime="00:03:51.85" />
                    <SPLIT distance="300" swimtime="00:04:38.74" />
                    <SPLIT distance="350" swimtime="00:05:25.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="20896" name="Swim Academy Krakow">
          <CONTACT email="lukasz.giminski@gmail.com" internet="www.swimacademy.pl" name="Łukasz Gimiński" phone="721404110" />
          <ATHLETES>
            <ATHLETE birthdate="1978-04-10" firstname="Alina" gender="F" lastname="Handzlik" nation="POL" athleteid="20897">
              <RESULTS>
                <RESULT eventid="1147" points="240" reactiontime="+118" swimtime="00:12:59.74" resultid="20898" heatid="24311" lane="8" entrytime="00:13:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.85" />
                    <SPLIT distance="100" swimtime="00:03:14.25" />
                    <SPLIT distance="150" swimtime="00:02:24.09" />
                    <SPLIT distance="250" swimtime="00:04:05.16" />
                    <SPLIT distance="350" swimtime="00:05:45.22" />
                    <SPLIT distance="400" swimtime="00:06:34.88" />
                    <SPLIT distance="450" swimtime="00:07:24.08" />
                    <SPLIT distance="500" swimtime="00:08:13.89" />
                    <SPLIT distance="550" swimtime="00:09:02.58" />
                    <SPLIT distance="600" swimtime="00:11:27.82" />
                    <SPLIT distance="650" swimtime="00:10:39.66" />
                    <SPLIT distance="750" swimtime="00:12:16.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="23011" name="Swim Club Masters Ślęza">
          <CONTACT name="Bloch" />
          <ATHLETES>
            <ATHLETE birthdate="1972-03-11" firstname="Dorota" gender="F" lastname="Batóg" nation="POL" athleteid="23350">
              <RESULTS>
                <RESULT eventid="1062" points="345" reactiontime="+90" swimtime="00:00:33.73" resultid="23351" heatid="24279" lane="8" entrytime="00:00:33.30" />
                <RESULT eventid="1187" points="298" swimtime="00:00:40.47" resultid="23352" heatid="24325" lane="3" entrytime="00:00:41.16" />
                <RESULT eventid="1256" points="276" reactiontime="+97" swimtime="00:01:19.37" resultid="23353" heatid="24351" lane="3" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="257" reactiontime="+55" swimtime="00:00:38.38" resultid="23354" heatid="24388" lane="0" entrytime="00:00:37.20" />
                <RESULT eventid="1457" points="204" reactiontime="+108" swimtime="00:01:38.45" resultid="23355" heatid="24401" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-12-15" firstname="Marta" gender="F" lastname="Burandt" nation="POL" athleteid="23362">
              <RESULTS>
                <RESULT eventid="1165" points="202" reactiontime="+95" swimtime="00:26:06.32" resultid="23363" heatid="24319" lane="7" entrytime="00:25:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.58" />
                    <SPLIT distance="100" swimtime="00:01:25.04" />
                    <SPLIT distance="150" swimtime="00:02:13.57" />
                    <SPLIT distance="200" swimtime="00:03:03.48" />
                    <SPLIT distance="250" swimtime="00:03:53.80" />
                    <SPLIT distance="300" swimtime="00:04:45.50" />
                    <SPLIT distance="350" swimtime="00:05:38.71" />
                    <SPLIT distance="400" swimtime="00:06:32.53" />
                    <SPLIT distance="450" swimtime="00:07:26.76" />
                    <SPLIT distance="500" swimtime="00:08:20.78" />
                    <SPLIT distance="550" swimtime="00:09:14.66" />
                    <SPLIT distance="600" swimtime="00:10:09.49" />
                    <SPLIT distance="650" swimtime="00:11:03.29" />
                    <SPLIT distance="700" swimtime="00:11:57.36" />
                    <SPLIT distance="750" swimtime="00:12:50.79" />
                    <SPLIT distance="800" swimtime="00:13:45.26" />
                    <SPLIT distance="850" swimtime="00:14:38.08" />
                    <SPLIT distance="900" swimtime="00:15:31.75" />
                    <SPLIT distance="950" swimtime="00:16:24.63" />
                    <SPLIT distance="1000" swimtime="00:17:17.16" />
                    <SPLIT distance="1050" swimtime="00:18:09.85" />
                    <SPLIT distance="1100" swimtime="00:19:02.82" />
                    <SPLIT distance="1150" swimtime="00:19:55.78" />
                    <SPLIT distance="1200" swimtime="00:20:48.39" />
                    <SPLIT distance="1250" swimtime="00:21:41.63" />
                    <SPLIT distance="1300" swimtime="00:22:35.06" />
                    <SPLIT distance="1350" swimtime="00:23:28.84" />
                    <SPLIT distance="1400" swimtime="00:24:22.30" />
                    <SPLIT distance="1450" swimtime="00:25:15.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="248" reactiontime="+103" swimtime="00:02:59.63" resultid="23364" heatid="24412" lane="3" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                    <SPLIT distance="100" swimtime="00:01:23.40" />
                    <SPLIT distance="150" swimtime="00:02:11.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-05-11" firstname="Joanna" gender="F" lastname="Krowicka" nation="POL" athleteid="23370">
              <RESULTS>
                <RESULT eventid="1222" points="217" reactiontime="+45" swimtime="00:03:51.23" resultid="23371" heatid="24339" lane="1" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.76" />
                    <SPLIT distance="100" swimtime="00:01:48.98" />
                    <SPLIT distance="150" swimtime="00:02:50.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="177" reactiontime="+55" swimtime="00:01:32.03" resultid="23372" heatid="24349" lane="1" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="213" reactiontime="+75" swimtime="00:01:47.36" resultid="23373" heatid="24377" lane="3" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="118" reactiontime="+89" swimtime="00:00:49.72" resultid="23374" heatid="24387" lane="8" entrytime="00:00:45.00" />
                <RESULT eventid="1664" status="DNS" swimtime="00:00:00.00" resultid="23375" heatid="24456" lane="1" entrytime="00:00:49.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-05-16" firstname="Mariusz" gender="M" lastname="Maciaszek" nation="POL" athleteid="23356">
              <RESULTS>
                <RESULT eventid="1079" points="469" reactiontime="+73" swimtime="00:00:26.90" resultid="23357" heatid="24293" lane="6" entrytime="00:00:27.01" />
                <RESULT eventid="1273" points="442" swimtime="00:01:01.54" resultid="23358" heatid="24362" lane="2" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="444" swimtime="00:00:29.18" resultid="23359" heatid="24396" lane="1" entrytime="00:00:29.23" />
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="23360" heatid="24440" lane="3" entrytime="00:01:10.00" />
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="23361" heatid="24464" lane="0" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-03-05" firstname="Dariusz" gender="M" lastname="Michalczuk" nation="POL" athleteid="23365">
              <RESULTS>
                <RESULT eventid="1079" points="235" reactiontime="+108" swimtime="00:00:33.87" resultid="23366" heatid="24288" lane="0" entrytime="00:00:32.00" />
                <RESULT eventid="14189" reactiontime="+106" status="OTL" swimtime="00:13:47.27" resultid="23367" heatid="24316" lane="3" entrytime="00:11:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.44" />
                    <SPLIT distance="100" swimtime="00:01:30.30" />
                    <SPLIT distance="150" swimtime="00:02:20.07" />
                    <SPLIT distance="200" swimtime="00:03:10.77" />
                    <SPLIT distance="250" swimtime="00:04:03.50" />
                    <SPLIT distance="300" swimtime="00:04:56.35" />
                    <SPLIT distance="350" swimtime="00:05:49.34" />
                    <SPLIT distance="400" swimtime="00:06:43.60" />
                    <SPLIT distance="450" swimtime="00:07:37.40" />
                    <SPLIT distance="500" swimtime="00:08:31.06" />
                    <SPLIT distance="550" swimtime="00:09:25.64" />
                    <SPLIT distance="600" swimtime="00:10:18.57" />
                    <SPLIT distance="700" swimtime="00:12:06.32" />
                    <SPLIT distance="750" swimtime="00:12:58.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="151" swimtime="00:00:44.98" resultid="23368" heatid="24332" lane="6" entrytime="00:00:39.50" />
                <RESULT eventid="1273" points="247" swimtime="00:01:14.71" resultid="23369" heatid="24357" lane="5" entrytime="00:01:14.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1698" status="DNS" swimtime="00:00:00.00" resultid="23376" heatid="24467" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="23350" number="1" />
                    <RELAYPOSITION athleteid="23362" number="2" />
                    <RELAYPOSITION athleteid="23356" number="3" />
                    <RELAYPOSITION athleteid="23365" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1130" reactiontime="+95" swimtime="00:02:06.69" resultid="23377" heatid="24308" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.48" />
                    <SPLIT distance="100" swimtime="00:01:08.13" />
                    <SPLIT distance="150" swimtime="00:01:34.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="23350" number="1" reactiontime="+95" />
                    <RELAYPOSITION athleteid="23362" number="2" />
                    <RELAYPOSITION athleteid="23356" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="23365" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="20466" name="Swim Tri Rzeszów">
          <CONTACT city="RZESZÓW" name="SWIM TRI RZESZÓW" street="POPIEŁUSZKI 26 C" zip="35-328" />
          <ATHLETES>
            <ATHLETE birthdate="1963-11-15" firstname="Mariusz" gender="M" lastname="Faff" nation="POL" athleteid="20467">
              <RESULTS>
                <RESULT eventid="1079" points="368" reactiontime="+100" swimtime="00:00:29.17" resultid="20468" heatid="24291" lane="6" entrytime="00:00:29.00" entrycourse="LCM" />
                <RESULT eventid="1113" points="260" reactiontime="+91" swimtime="00:02:58.54" resultid="20469" heatid="24304" lane="1" entrytime="00:03:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                    <SPLIT distance="100" swimtime="00:01:23.78" />
                    <SPLIT distance="150" swimtime="00:02:21.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="288" swimtime="00:00:36.33" resultid="20470" heatid="24333" lane="8" entrytime="00:00:36.32" entrycourse="LCM" />
                <RESULT eventid="1273" points="353" reactiontime="+88" swimtime="00:01:06.32" resultid="20471" heatid="24360" lane="4" entrytime="00:01:05.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="339" swimtime="00:00:31.92" resultid="20472" heatid="24394" lane="3" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="1508" points="295" reactiontime="+41" swimtime="00:02:33.06" resultid="20473" heatid="24421" lane="8" entrytime="00:02:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                    <SPLIT distance="100" swimtime="00:01:12.70" />
                    <SPLIT distance="150" swimtime="00:01:53.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="298" reactiontime="+75" swimtime="00:05:29.35" resultid="20474" heatid="24479" lane="4" entrytime="00:05:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.84" />
                    <SPLIT distance="100" swimtime="00:01:16.47" />
                    <SPLIT distance="150" swimtime="00:01:59.01" />
                    <SPLIT distance="200" swimtime="00:02:41.37" />
                    <SPLIT distance="250" swimtime="00:03:24.68" />
                    <SPLIT distance="300" swimtime="00:04:07.16" />
                    <SPLIT distance="350" swimtime="00:04:49.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="ZAC" clubid="20621" name="Swimming Masters Team Szczecin">
          <CONTACT city="Mierzyn" email="marekzet74@gmail.com" name="Zienkiewicz" phone="+48500641651" state="ZACHO" street="teresy 58" zip="72-006" />
          <ATHLETES>
            <ATHLETE birthdate="1987-08-03" firstname="Edyta" gender="F" lastname="Adamiak" nation="POL" athleteid="20637">
              <RESULTS>
                <RESULT eventid="1062" points="177" reactiontime="+102" swimtime="00:00:42.14" resultid="20638" heatid="24276" lane="5" entrytime="00:00:48.00" />
                <RESULT eventid="1147" reactiontime="+102" status="OTL" swimtime="00:15:31.95" resultid="20639" heatid="24310" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.14" />
                    <SPLIT distance="100" swimtime="00:01:42.21" />
                    <SPLIT distance="150" swimtime="00:02:40.91" />
                    <SPLIT distance="200" swimtime="00:03:40.43" />
                    <SPLIT distance="250" swimtime="00:04:39.53" />
                    <SPLIT distance="300" swimtime="00:05:38.79" />
                    <SPLIT distance="350" swimtime="00:06:38.75" />
                    <SPLIT distance="400" swimtime="00:07:39.39" />
                    <SPLIT distance="450" swimtime="00:08:39.29" />
                    <SPLIT distance="500" swimtime="00:09:39.53" />
                    <SPLIT distance="550" swimtime="00:10:39.05" />
                    <SPLIT distance="600" swimtime="00:11:39.04" />
                    <SPLIT distance="650" swimtime="00:12:38.36" />
                    <SPLIT distance="700" swimtime="00:13:37.44" />
                    <SPLIT distance="750" swimtime="00:14:36.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="140" reactiontime="+65" swimtime="00:01:39.48" resultid="20640" heatid="24349" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="157" reactiontime="+62" swimtime="00:03:29.09" resultid="20641" heatid="24411" lane="6" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.95" />
                    <SPLIT distance="100" swimtime="00:01:40.95" />
                    <SPLIT distance="150" swimtime="00:02:36.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="179" reactiontime="+50" swimtime="00:00:52.10" resultid="20642" heatid="24456" lane="0" entrytime="00:00:50.00" />
                <RESULT eventid="1721" points="145" reactiontime="+98" swimtime="00:07:30.09" resultid="20643" heatid="24470" lane="4" entrytime="00:07:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.35" />
                    <SPLIT distance="100" swimtime="00:01:46.21" />
                    <SPLIT distance="150" swimtime="00:02:43.72" />
                    <SPLIT distance="200" swimtime="00:03:41.68" />
                    <SPLIT distance="250" swimtime="00:04:40.64" />
                    <SPLIT distance="300" swimtime="00:05:38.66" />
                    <SPLIT distance="350" swimtime="00:06:36.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-03-27" firstname="Marek" gender="M" lastname="Piotrowski" nation="POL" athleteid="20630">
              <RESULTS>
                <RESULT eventid="1079" points="320" reactiontime="+84" swimtime="00:00:30.55" resultid="20631" heatid="24289" lane="0" entrytime="00:00:31.00" />
                <RESULT eventid="1205" points="165" swimtime="00:00:43.67" resultid="20632" heatid="24328" lane="7" />
                <RESULT eventid="1273" points="323" swimtime="00:01:08.30" resultid="20633" heatid="24359" lane="8" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="233" swimtime="00:00:36.16" resultid="20634" heatid="24392" lane="5" entrytime="00:00:37.00" />
                <RESULT eventid="1508" points="243" swimtime="00:02:43.28" resultid="20635" heatid="24419" lane="6" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                    <SPLIT distance="100" swimtime="00:01:15.60" />
                    <SPLIT distance="150" swimtime="00:01:58.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="224" swimtime="00:06:01.96" resultid="20636" heatid="24478" lane="6" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.07" />
                    <SPLIT distance="100" swimtime="00:01:21.08" />
                    <SPLIT distance="150" swimtime="00:02:06.11" />
                    <SPLIT distance="200" swimtime="00:02:52.47" />
                    <SPLIT distance="250" swimtime="00:03:40.22" />
                    <SPLIT distance="300" swimtime="00:04:28.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-05-09" firstname="Łukasz" gender="M" lastname="Rożek" nation="POL" athleteid="20622">
              <RESULTS>
                <RESULT eventid="1079" points="257" reactiontime="+82" swimtime="00:00:32.87" resultid="20623" heatid="24287" lane="9" entrytime="00:00:34.00" />
                <RESULT eventid="14189" points="166" reactiontime="+86" swimtime="00:13:41.14" resultid="20624" heatid="24313" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.99" />
                    <SPLIT distance="100" swimtime="00:01:25.19" />
                    <SPLIT distance="150" swimtime="00:02:14.78" />
                    <SPLIT distance="200" swimtime="00:03:04.59" />
                    <SPLIT distance="250" swimtime="00:03:56.74" />
                    <SPLIT distance="300" swimtime="00:06:35.84" />
                    <SPLIT distance="350" swimtime="00:05:42.88" />
                    <SPLIT distance="450" swimtime="00:07:29.56" />
                    <SPLIT distance="500" swimtime="00:08:22.78" />
                    <SPLIT distance="550" swimtime="00:09:15.51" />
                    <SPLIT distance="600" swimtime="00:10:09.34" />
                    <SPLIT distance="650" swimtime="00:11:02.77" />
                    <SPLIT distance="700" swimtime="00:11:56.67" />
                    <SPLIT distance="750" swimtime="00:12:50.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="223" swimtime="00:01:17.30" resultid="20625" heatid="24357" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="172" swimtime="00:00:39.99" resultid="20626" heatid="24391" lane="1" entrytime="00:00:45.15" />
                <RESULT eventid="1508" points="189" reactiontime="+43" swimtime="00:02:57.63" resultid="20627" heatid="24418" lane="8" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                    <SPLIT distance="100" swimtime="00:01:23.36" />
                    <SPLIT distance="150" swimtime="00:02:10.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="155" swimtime="00:00:48.28" resultid="20628" heatid="24460" lane="3" entrytime="00:00:49.57" />
                <RESULT eventid="1744" points="184" reactiontime="+50" swimtime="00:06:26.82" resultid="20629" heatid="24476" lane="2" entrytime="00:07:01.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.53" />
                    <SPLIT distance="100" swimtime="00:01:28.37" />
                    <SPLIT distance="150" swimtime="00:02:16.90" />
                    <SPLIT distance="200" swimtime="00:03:07.12" />
                    <SPLIT distance="250" swimtime="00:03:57.08" />
                    <SPLIT distance="300" swimtime="00:04:48.22" />
                    <SPLIT distance="350" swimtime="00:05:38.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-12-12" firstname="Dominika" gender="F" lastname="Zielińska" nation="POL" athleteid="20644">
              <RESULTS>
                <RESULT eventid="1096" points="374" reactiontime="+76" swimtime="00:02:55.00" resultid="20645" heatid="24299" lane="7" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                    <SPLIT distance="100" swimtime="00:01:19.09" />
                    <SPLIT distance="150" swimtime="00:02:12.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="373" swimtime="00:00:37.59" resultid="20646" heatid="24326" lane="0" entrytime="00:00:40.00" />
                <RESULT eventid="1256" points="410" swimtime="00:01:09.56" resultid="20647" heatid="24352" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="372" reactiontime="+77" swimtime="00:01:20.58" resultid="20648" heatid="24402" lane="0" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="379" reactiontime="+72" swimtime="00:02:36.09" resultid="20649" heatid="24413" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.29" />
                    <SPLIT distance="100" swimtime="00:01:15.04" />
                    <SPLIT distance="150" swimtime="00:01:55.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="372" reactiontime="+64" swimtime="00:02:52.46" resultid="20650" heatid="24445" lane="8" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.84" />
                    <SPLIT distance="100" swimtime="00:01:24.24" />
                    <SPLIT distance="150" swimtime="00:02:08.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="337" reactiontime="+69" swimtime="00:05:39.57" resultid="20651" heatid="24472" lane="6" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                    <SPLIT distance="100" swimtime="00:01:17.65" />
                    <SPLIT distance="150" swimtime="00:02:00.41" />
                    <SPLIT distance="200" swimtime="00:02:44.11" />
                    <SPLIT distance="250" swimtime="00:03:27.58" />
                    <SPLIT distance="300" swimtime="00:04:12.60" />
                    <SPLIT distance="350" swimtime="00:04:56.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-11-04" firstname="Kamil" gender="M" lastname="Zieliński" nation="POL" athleteid="20652">
              <RESULTS>
                <RESULT eventid="1079" points="256" reactiontime="+85" swimtime="00:00:32.93" resultid="20653" heatid="24284" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1205" points="214" swimtime="00:00:40.12" resultid="20654" heatid="24330" lane="2" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" reactiontime="+86" swimtime="00:02:17.02" resultid="20655" heatid="24309" lane="0" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.16" />
                    <SPLIT distance="100" swimtime="00:01:02.38" />
                    <SPLIT distance="150" swimtime="00:01:44.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="20630" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="20644" number="2" />
                    <RELAYPOSITION athleteid="20637" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="20622" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" reactiontime="+78" swimtime="00:02:40.94" resultid="20656" heatid="24467" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.62" />
                    <SPLIT distance="150" swimtime="00:02:06.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="20652" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="20637" number="2" />
                    <RELAYPOSITION athleteid="20644" number="3" reactiontime="+9" />
                    <RELAYPOSITION athleteid="20622" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="21246" name="T.P.Masters Opole">
          <CONTACT city="OPOLE" name="KRASNODĘBSKI" />
          <ATHLETES>
            <ATHLETE birthdate="1990-01-01" firstname="Agnieszka" gender="F" lastname="Bartnikowska" nation="POL" athleteid="21260">
              <RESULTS>
                <RESULT eventid="1062" points="526" reactiontime="+82" swimtime="00:00:29.31" resultid="21261" heatid="24280" lane="3" entrytime="00:00:30.22" />
                <RESULT eventid="1096" points="492" reactiontime="+81" swimtime="00:02:39.72" resultid="21262" heatid="24299" lane="6" entrytime="00:02:41.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.71" />
                    <SPLIT distance="100" swimtime="00:01:13.56" />
                    <SPLIT distance="150" swimtime="00:02:02.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-01" firstname="Zbigniew" gender="M" lastname="Januszkiewicz" nation="POL" athleteid="21254">
              <RESULTS>
                <RESULT eventid="1079" points="399" reactiontime="+90" swimtime="00:00:28.39" resultid="21255" heatid="24291" lane="0" entrytime="00:00:29.13" />
                <RESULT eventid="1113" points="384" reactiontime="+84" swimtime="00:02:36.73" resultid="21256" heatid="24305" lane="3" entrytime="00:02:39.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                    <SPLIT distance="100" swimtime="00:01:11.35" />
                    <SPLIT distance="150" swimtime="00:02:00.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="393" reactiontime="+72" swimtime="00:00:32.74" resultid="21257" heatid="24335" lane="0" entrytime="00:00:31.56" />
                <RESULT eventid="1474" points="415" swimtime="00:01:09.48" resultid="21258" heatid="24407" lane="5" entrytime="00:01:08.88" />
                <RESULT eventid="1647" points="415" reactiontime="+73" swimtime="00:02:30.00" resultid="21259" heatid="24452" lane="1" entrytime="00:02:26.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.40" />
                    <SPLIT distance="100" swimtime="00:01:12.94" />
                    <SPLIT distance="150" swimtime="00:01:51.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Minkiewicz" gender="M" lastname="Jerzy" nation="POL" athleteid="21263">
              <RESULTS>
                <RESULT eventid="1079" points="260" reactiontime="+92" swimtime="00:00:32.74" resultid="21264" heatid="24288" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="1273" points="250" reactiontime="+48" swimtime="00:01:14.38" resultid="21265" heatid="24358" lane="1" entrytime="00:01:12.00" />
                <RESULT eventid="1440" points="210" reactiontime="+60" swimtime="00:00:37.41" resultid="21266" heatid="24393" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="1613" points="125" swimtime="00:01:39.62" resultid="21267" heatid="24439" lane="9" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Zbigniew" gender="M" lastname="Krasnodębski" nation="POL" athleteid="21268">
              <RESULTS>
                <RESULT eventid="1681" points="218" reactiontime="+52" swimtime="00:00:43.06" resultid="21269" heatid="24461" lane="3" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Tomasz" gender="M" lastname="Samsel" nation="POL" athleteid="21247">
              <RESULTS>
                <RESULT eventid="1079" points="524" reactiontime="+69" swimtime="00:00:25.92" resultid="21248" heatid="24296" lane="9" entrytime="00:00:25.60" />
                <RESULT eventid="1113" points="443" reactiontime="+78" swimtime="00:02:29.44" resultid="21249" heatid="24306" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                    <SPLIT distance="100" swimtime="00:01:11.73" />
                    <SPLIT distance="150" swimtime="00:01:56.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="385" reactiontime="+83" swimtime="00:00:32.97" resultid="21250" heatid="24334" lane="1" entrytime="00:00:33.30" />
                <RESULT eventid="1273" points="519" reactiontime="+70" swimtime="00:00:58.36" resultid="21251" heatid="24365" lane="8" entrytime="00:00:56.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="362" reactiontime="+70" swimtime="00:01:12.71" resultid="21252" heatid="24406" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="443" swimtime="00:02:13.75" resultid="21253" heatid="24422" lane="2" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                    <SPLIT distance="100" swimtime="00:01:05.69" />
                    <SPLIT distance="150" swimtime="00:01:40.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="ZAC" clubid="21818" name="TKKF Koszalin Masters">
          <CONTACT email="rpieslak@wp.pl" name="Pieślak Roman" phone="600227112" />
          <ATHLETES>
            <ATHLETE birthdate="1960-08-26" firstname="Dorota" gender="F" lastname="Gudaniec" nation="POL" athleteid="21861">
              <RESULTS>
                <RESULT eventid="1165" points="221" reactiontime="+73" swimtime="00:25:20.63" resultid="21862" heatid="24319" lane="2" entrytime="00:25:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.45" />
                    <SPLIT distance="100" swimtime="00:01:32.58" />
                    <SPLIT distance="150" swimtime="00:02:22.97" />
                    <SPLIT distance="200" swimtime="00:03:13.63" />
                    <SPLIT distance="250" swimtime="00:04:05.12" />
                    <SPLIT distance="300" swimtime="00:04:56.22" />
                    <SPLIT distance="350" swimtime="00:05:46.59" />
                    <SPLIT distance="400" swimtime="00:06:38.24" />
                    <SPLIT distance="450" swimtime="00:07:29.68" />
                    <SPLIT distance="500" swimtime="00:08:20.56" />
                    <SPLIT distance="550" swimtime="00:09:11.41" />
                    <SPLIT distance="600" swimtime="00:10:02.50" />
                    <SPLIT distance="650" swimtime="00:10:53.52" />
                    <SPLIT distance="700" swimtime="00:11:43.94" />
                    <SPLIT distance="750" swimtime="00:12:35.25" />
                    <SPLIT distance="800" swimtime="00:13:26.69" />
                    <SPLIT distance="850" swimtime="00:14:18.04" />
                    <SPLIT distance="900" swimtime="00:15:08.91" />
                    <SPLIT distance="950" swimtime="00:15:59.86" />
                    <SPLIT distance="1000" swimtime="00:16:51.44" />
                    <SPLIT distance="1050" swimtime="00:17:42.84" />
                    <SPLIT distance="1100" swimtime="00:18:33.56" />
                    <SPLIT distance="1150" swimtime="00:19:24.60" />
                    <SPLIT distance="1200" swimtime="00:20:15.76" />
                    <SPLIT distance="1250" swimtime="00:21:07.12" />
                    <SPLIT distance="1300" swimtime="00:21:58.24" />
                    <SPLIT distance="1350" swimtime="00:22:49.18" />
                    <SPLIT distance="1400" swimtime="00:23:40.46" />
                    <SPLIT distance="1450" swimtime="00:24:31.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="180" swimtime="00:00:47.84" resultid="21863" heatid="24325" lane="6" entrytime="00:00:42.00" />
                <RESULT eventid="1222" points="191" reactiontime="+61" swimtime="00:04:01.38" resultid="21864" heatid="24339" lane="3" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.38" />
                    <SPLIT distance="100" swimtime="00:01:53.35" />
                    <SPLIT distance="150" swimtime="00:02:56.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="176" swimtime="00:01:43.35" resultid="21865" heatid="24400" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="205" reactiontime="+69" swimtime="00:07:31.30" resultid="21866" heatid="24429" lane="1" entrytime="00:07:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.87" />
                    <SPLIT distance="100" swimtime="00:01:49.00" />
                    <SPLIT distance="150" swimtime="00:04:47.95" />
                    <SPLIT distance="200" swimtime="00:03:45.25" />
                    <SPLIT distance="250" swimtime="00:06:42.39" />
                    <SPLIT distance="300" swimtime="00:05:51.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="169" reactiontime="+91" swimtime="00:03:43.97" resultid="21867" heatid="24444" lane="0" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.19" />
                    <SPLIT distance="150" swimtime="00:02:47.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="206" reactiontime="+96" swimtime="00:06:39.84" resultid="21868" heatid="24471" lane="3" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.84" />
                    <SPLIT distance="100" swimtime="00:01:35.08" />
                    <SPLIT distance="150" swimtime="00:02:26.22" />
                    <SPLIT distance="200" swimtime="00:03:17.64" />
                    <SPLIT distance="250" swimtime="00:04:08.27" />
                    <SPLIT distance="300" swimtime="00:05:00.18" />
                    <SPLIT distance="350" swimtime="00:05:50.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-07-15" firstname="Marian" gender="M" lastname="Lasowy" nation="POL" athleteid="21834">
              <RESULTS>
                <RESULT eventid="14207" points="159" reactiontime="+128" swimtime="00:26:46.31" resultid="21835" heatid="24320" lane="3" entrytime="00:27:16.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.30" />
                    <SPLIT distance="100" swimtime="00:01:38.50" />
                    <SPLIT distance="150" swimtime="00:02:32.04" />
                    <SPLIT distance="200" swimtime="00:03:25.48" />
                    <SPLIT distance="250" swimtime="00:04:20.14" />
                    <SPLIT distance="300" swimtime="00:05:13.75" />
                    <SPLIT distance="350" swimtime="00:06:08.23" />
                    <SPLIT distance="400" swimtime="00:07:02.08" />
                    <SPLIT distance="450" swimtime="00:07:55.97" />
                    <SPLIT distance="500" swimtime="00:08:49.87" />
                    <SPLIT distance="550" swimtime="00:09:43.85" />
                    <SPLIT distance="600" swimtime="00:10:37.59" />
                    <SPLIT distance="650" swimtime="00:11:31.75" />
                    <SPLIT distance="700" swimtime="00:12:26.17" />
                    <SPLIT distance="750" swimtime="00:13:20.48" />
                    <SPLIT distance="800" swimtime="00:14:14.65" />
                    <SPLIT distance="850" swimtime="00:15:08.61" />
                    <SPLIT distance="900" swimtime="00:16:02.66" />
                    <SPLIT distance="950" swimtime="00:16:56.84" />
                    <SPLIT distance="1000" swimtime="00:17:50.93" />
                    <SPLIT distance="1050" swimtime="00:18:45.28" />
                    <SPLIT distance="1100" swimtime="00:19:39.27" />
                    <SPLIT distance="1150" swimtime="00:20:33.59" />
                    <SPLIT distance="1200" swimtime="00:21:27.47" />
                    <SPLIT distance="1250" swimtime="00:22:21.26" />
                    <SPLIT distance="1300" swimtime="00:23:14.99" />
                    <SPLIT distance="1350" swimtime="00:24:09.43" />
                    <SPLIT distance="1400" swimtime="00:25:03.84" />
                    <SPLIT distance="1450" swimtime="00:25:58.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="96" reactiontime="+74" swimtime="00:04:04.00" resultid="21836" heatid="24448" lane="9" entrytime="00:04:00.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.39" />
                    <SPLIT distance="100" swimtime="00:04:03.94" />
                    <SPLIT distance="150" swimtime="00:03:03.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="143" reactiontime="+112" swimtime="00:07:00.53" resultid="21837" heatid="24476" lane="3" entrytime="00:06:51.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.46" />
                    <SPLIT distance="100" swimtime="00:01:37.26" />
                    <SPLIT distance="150" swimtime="00:02:32.29" />
                    <SPLIT distance="200" swimtime="00:03:26.81" />
                    <SPLIT distance="250" swimtime="00:04:21.61" />
                    <SPLIT distance="300" swimtime="00:05:15.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-02-24" firstname="Wioletta" gender="F" lastname="Pawliczek" nation="POL" athleteid="21819">
              <RESULTS>
                <RESULT eventid="1062" points="335" reactiontime="+83" swimtime="00:00:34.07" resultid="21820" heatid="24278" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1187" points="311" swimtime="00:00:39.91" resultid="21821" heatid="24326" lane="9" entrytime="00:00:40.00" />
                <RESULT eventid="1256" points="303" reactiontime="+53" swimtime="00:01:16.97" resultid="21822" heatid="24351" lane="0" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="300" reactiontime="+82" swimtime="00:01:26.57" resultid="21823" heatid="24401" lane="1" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="267" reactiontime="+70" swimtime="00:03:12.64" resultid="21824" heatid="24444" lane="5" entrytime="00:03:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-05" firstname="Agnieszka" gender="F" lastname="Paziewska" nation="POL" athleteid="21838">
              <RESULTS>
                <RESULT eventid="1062" points="365" reactiontime="+89" swimtime="00:00:33.12" resultid="21839" heatid="24280" lane="9" entrytime="00:00:32.45" />
                <RESULT eventid="1388" points="201" reactiontime="+68" swimtime="00:01:49.34" resultid="21840" heatid="24378" lane="1" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="267" reactiontime="+64" swimtime="00:02:55.32" resultid="21841" heatid="24413" lane="0" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                    <SPLIT distance="100" swimtime="00:01:20.82" />
                    <SPLIT distance="150" swimtime="00:02:08.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-28" firstname="Roman" gender="M" lastname="Pieślak" nation="POL" athleteid="21847">
              <RESULTS>
                <RESULT eventid="1079" points="366" reactiontime="+79" swimtime="00:00:29.23" resultid="21848" heatid="24290" lane="6" entrytime="00:00:29.50" />
                <RESULT eventid="1239" points="330" swimtime="00:03:03.19" resultid="21849" heatid="24345" lane="7" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.32" />
                    <SPLIT distance="100" swimtime="00:01:28.10" />
                    <SPLIT distance="150" swimtime="00:02:15.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="346" swimtime="00:01:06.78" resultid="21850" heatid="24361" lane="9" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="333" reactiontime="+69" swimtime="00:01:22.35" resultid="21851" heatid="24384" lane="8" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="301" swimtime="00:02:32.16" resultid="21852" heatid="24421" lane="6" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                    <SPLIT distance="100" swimtime="00:01:13.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="368" swimtime="00:00:36.21" resultid="21853" heatid="24464" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="1744" points="294" swimtime="00:05:30.77" resultid="21854" heatid="24479" lane="5" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.23" />
                    <SPLIT distance="200" swimtime="00:02:42.45" />
                    <SPLIT distance="300" swimtime="00:04:09.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-02-20" firstname="Artur" gender="M" lastname="Rutkowski" nation="POL" athleteid="21869">
              <RESULTS>
                <RESULT eventid="1113" points="277" reactiontime="+96" swimtime="00:02:54.73" resultid="21870" heatid="24304" lane="6" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                    <SPLIT distance="100" swimtime="00:01:24.58" />
                    <SPLIT distance="150" swimtime="00:02:15.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14189" points="265" reactiontime="+101" swimtime="00:11:43.02" resultid="21871" heatid="24315" lane="2" entrytime="00:12:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.90" />
                    <SPLIT distance="100" swimtime="00:01:21.22" />
                    <SPLIT distance="150" swimtime="00:02:04.68" />
                    <SPLIT distance="200" swimtime="00:02:48.66" />
                    <SPLIT distance="250" swimtime="00:03:32.92" />
                    <SPLIT distance="300" swimtime="00:04:17.49" />
                    <SPLIT distance="350" swimtime="00:05:02.72" />
                    <SPLIT distance="400" swimtime="00:05:47.93" />
                    <SPLIT distance="450" swimtime="00:06:32.97" />
                    <SPLIT distance="500" swimtime="00:07:17.83" />
                    <SPLIT distance="550" swimtime="00:08:03.78" />
                    <SPLIT distance="600" swimtime="00:08:49.04" />
                    <SPLIT distance="650" swimtime="00:09:35.11" />
                    <SPLIT distance="700" swimtime="00:10:19.76" />
                    <SPLIT distance="750" swimtime="00:11:03.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="220" reactiontime="+70" swimtime="00:03:04.71" resultid="21872" heatid="24370" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.87" />
                    <SPLIT distance="100" swimtime="00:01:28.27" />
                    <SPLIT distance="150" swimtime="00:02:18.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="346" reactiontime="+42" swimtime="00:00:31.70" resultid="21873" heatid="24394" lane="8" entrytime="00:00:32.50" />
                <RESULT eventid="1578" status="DNS" swimtime="00:00:00.00" resultid="21874" heatid="24432" lane="8" entrytime="00:06:15.00" />
                <RESULT eventid="1613" points="257" reactiontime="+55" swimtime="00:01:18.33" resultid="21875" heatid="24439" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-07-05" firstname="Krzysztof" gender="M" lastname="Stefański" nation="POL" athleteid="21876">
              <RESULTS>
                <RESULT eventid="1079" points="375" reactiontime="+86" swimtime="00:00:28.99" resultid="21877" heatid="24286" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="21878" heatid="24304" lane="8" entrytime="00:03:00.00" />
                <RESULT eventid="1273" points="341" reactiontime="+84" swimtime="00:01:07.11" resultid="21879" heatid="24360" lane="2" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="285" reactiontime="+77" swimtime="00:00:33.82" resultid="21880" heatid="24393" lane="3" entrytime="00:00:34.00" />
                <RESULT eventid="1681" points="226" reactiontime="+86" swimtime="00:00:42.55" resultid="21881" heatid="24463" lane="2" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-02-25" firstname="Tomasz" gender="M" lastname="Szymanowski" nation="POL" athleteid="21855">
              <RESULTS>
                <RESULT eventid="1079" points="381" reactiontime="+86" swimtime="00:00:28.83" resultid="21856" heatid="24291" lane="5" entrytime="00:00:28.80" />
                <RESULT eventid="14189" points="260" reactiontime="+103" swimtime="00:11:48.05" resultid="21857" heatid="24316" lane="9" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.77" />
                    <SPLIT distance="100" swimtime="00:01:19.86" />
                    <SPLIT distance="150" swimtime="00:02:03.02" />
                    <SPLIT distance="200" swimtime="00:02:47.42" />
                    <SPLIT distance="250" swimtime="00:03:32.22" />
                    <SPLIT distance="300" swimtime="00:04:16.93" />
                    <SPLIT distance="350" swimtime="00:05:01.98" />
                    <SPLIT distance="400" swimtime="00:05:47.61" />
                    <SPLIT distance="450" swimtime="00:06:32.69" />
                    <SPLIT distance="500" swimtime="00:07:18.74" />
                    <SPLIT distance="550" swimtime="00:08:04.06" />
                    <SPLIT distance="600" swimtime="00:08:50.35" />
                    <SPLIT distance="650" swimtime="00:09:36.63" />
                    <SPLIT distance="700" swimtime="00:10:22.18" />
                    <SPLIT distance="750" swimtime="00:11:07.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="354" swimtime="00:00:33.90" resultid="21858" heatid="24333" lane="4" entrytime="00:00:34.00" />
                <RESULT eventid="1474" points="320" swimtime="00:01:15.75" resultid="21859" heatid="24406" lane="4" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="286" reactiontime="+99" swimtime="00:02:49.72" resultid="21860" heatid="24450" lane="7" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.35" />
                    <SPLIT distance="100" swimtime="00:01:24.17" />
                    <SPLIT distance="150" swimtime="00:02:07.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-11-16" firstname="Dawid" gender="M" lastname="Wróblewski" nation="POL" athleteid="21882">
              <RESULTS>
                <RESULT eventid="1079" points="569" reactiontime="+82" swimtime="00:00:25.22" resultid="21883" heatid="24295" lane="0" entrytime="00:00:26.15" />
                <RESULT eventid="1113" points="466" reactiontime="+75" swimtime="00:02:27.03" resultid="21884" heatid="24306" lane="8" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.18" />
                    <SPLIT distance="100" swimtime="00:01:11.92" />
                    <SPLIT distance="150" swimtime="00:01:52.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="506" swimtime="00:02:38.91" resultid="21885" heatid="24345" lane="5" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="561" swimtime="00:00:26.99" resultid="21886" heatid="24397" lane="6" entrytime="00:00:27.30" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="21887" heatid="24423" lane="8" entrytime="00:02:13.00" />
                <RESULT eventid="1613" points="557" swimtime="00:01:00.54" resultid="21888" heatid="24441" lane="3" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="21889" heatid="24481" lane="8" entrytime="00:05:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-04-14" firstname="Wiesław" gender="M" lastname="Załuski" nation="POL" athleteid="21842">
              <RESULTS>
                <RESULT eventid="1113" points="235" reactiontime="+102" swimtime="00:03:04.62" resultid="21843" heatid="24303" lane="2" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                    <SPLIT distance="100" swimtime="00:01:25.45" />
                    <SPLIT distance="150" swimtime="00:02:21.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="267" swimtime="00:00:37.27" resultid="21844" heatid="24332" lane="4" entrytime="00:00:37.50" />
                <RESULT eventid="1440" points="257" reactiontime="+66" swimtime="00:00:35.01" resultid="21845" heatid="24392" lane="8" entrytime="00:00:38.50" />
                <RESULT eventid="1613" points="181" reactiontime="+66" swimtime="00:01:28.05" resultid="21846" heatid="24439" lane="8" entrytime="00:01:32.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-08-22" firstname="Grzegorz" gender="M" lastname="Ćwikła" nation="POL" athleteid="21825">
              <RESULTS>
                <RESULT eventid="1079" points="317" reactiontime="+88" swimtime="00:00:30.66" resultid="21826" heatid="24292" lane="1" entrytime="00:00:28.42" />
                <RESULT eventid="14207" points="247" reactiontime="+93" swimtime="00:23:08.19" resultid="21827" heatid="24322" lane="0" entrytime="00:21:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.94" />
                    <SPLIT distance="100" swimtime="00:01:23.23" />
                    <SPLIT distance="150" swimtime="00:02:09.15" />
                    <SPLIT distance="200" swimtime="00:02:55.47" />
                    <SPLIT distance="250" swimtime="00:03:41.64" />
                    <SPLIT distance="300" swimtime="00:04:28.20" />
                    <SPLIT distance="350" swimtime="00:05:14.40" />
                    <SPLIT distance="400" swimtime="00:06:00.45" />
                    <SPLIT distance="450" swimtime="00:06:46.54" />
                    <SPLIT distance="500" swimtime="00:07:32.87" />
                    <SPLIT distance="550" swimtime="00:08:19.62" />
                    <SPLIT distance="600" swimtime="00:09:06.27" />
                    <SPLIT distance="650" swimtime="00:09:53.30" />
                    <SPLIT distance="700" swimtime="00:10:40.06" />
                    <SPLIT distance="750" swimtime="00:11:26.79" />
                    <SPLIT distance="800" swimtime="00:12:13.97" />
                    <SPLIT distance="850" swimtime="00:13:00.75" />
                    <SPLIT distance="900" swimtime="00:13:47.96" />
                    <SPLIT distance="950" swimtime="00:14:34.71" />
                    <SPLIT distance="1000" swimtime="00:15:22.04" />
                    <SPLIT distance="1050" swimtime="00:16:09.11" />
                    <SPLIT distance="1100" swimtime="00:16:56.70" />
                    <SPLIT distance="1150" swimtime="00:17:44.01" />
                    <SPLIT distance="1200" swimtime="00:18:31.71" />
                    <SPLIT distance="1250" swimtime="00:19:19.09" />
                    <SPLIT distance="1300" swimtime="00:20:06.68" />
                    <SPLIT distance="1350" swimtime="00:20:54.01" />
                    <SPLIT distance="1400" swimtime="00:21:40.96" />
                    <SPLIT distance="1450" swimtime="00:22:26.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="344" swimtime="00:00:34.23" resultid="21828" heatid="24334" lane="8" entrytime="00:00:33.54" />
                <RESULT eventid="1273" points="350" reactiontime="+77" swimtime="00:01:06.56" resultid="21829" heatid="24361" lane="3" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="301" reactiontime="+62" swimtime="00:01:17.29" resultid="21830" heatid="24407" lane="7" entrytime="00:01:13.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="296" reactiontime="+78" swimtime="00:02:33.02" resultid="21831" heatid="24421" lane="3" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                    <SPLIT distance="100" swimtime="00:01:14.76" />
                    <SPLIT distance="150" swimtime="00:01:54.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="236" swimtime="00:03:01.00" resultid="21832" heatid="24450" lane="6" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.18" />
                    <SPLIT distance="100" swimtime="00:01:29.31" />
                    <SPLIT distance="150" swimtime="00:02:16.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="273" swimtime="00:05:39.02" resultid="21833" heatid="24480" lane="0" entrytime="00:05:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                    <SPLIT distance="100" swimtime="00:01:17.27" />
                    <SPLIT distance="150" swimtime="00:01:59.67" />
                    <SPLIT distance="200" swimtime="00:02:43.82" />
                    <SPLIT distance="250" swimtime="00:03:27.35" />
                    <SPLIT distance="300" swimtime="00:04:12.75" />
                    <SPLIT distance="350" swimtime="00:04:57.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" name="TKKF Koszalin Masters - kat. C" number="2">
              <RESULTS>
                <RESULT comment="S1 - Pływak utracił kontakt stopami z platformą startową słupka zanim poprzedzający go pływak dotknął ściany (przedwczesna zmiana sztafetowa). (Time: 16:02), Na 3 zmianie" eventid="1381" reactiontime="+68" status="DSQ" swimtime="00:02:06.07" resultid="21892" heatid="24374" lane="1" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.61" />
                    <SPLIT distance="100" swimtime="00:01:10.91" />
                    <SPLIT distance="150" swimtime="00:01:37.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21825" number="1" reactiontime="+68" status="DSQ" />
                    <RELAYPOSITION athleteid="21847" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="21882" number="3" reactiontime="-7" status="DSQ" />
                    <RELAYPOSITION athleteid="21876" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" name="TKKF Koszalin Masters - kat. D" number="3">
              <RESULTS>
                <RESULT eventid="1548" points="361" reactiontime="+42" swimtime="00:01:59.13" resultid="21890" heatid="24427" lane="1" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.57" />
                    <SPLIT distance="100" swimtime="00:01:00.77" />
                    <SPLIT distance="150" swimtime="00:01:31.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21855" number="1" reactiontime="+42" />
                    <RELAYPOSITION athleteid="21842" number="2" />
                    <RELAYPOSITION athleteid="21869" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="21876" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="TKKF Koszalin Masters - kat. C" number="1">
              <RESULTS>
                <RESULT eventid="1130" reactiontime="+83" swimtime="00:02:01.23" resultid="21891" heatid="24309" lane="1" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.98" />
                    <SPLIT distance="100" swimtime="00:00:59.34" />
                    <SPLIT distance="150" swimtime="00:01:32.63" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21882" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="21838" number="2" />
                    <RELAYPOSITION athleteid="21819" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="21876" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" name="TKKF Koszalin Masters - kat. C" number="4">
              <RESULTS>
                <RESULT eventid="1698" reactiontime="+69" swimtime="00:02:20.98" resultid="21893" heatid="24468" lane="8" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.06" />
                    <SPLIT distance="100" swimtime="00:01:15.67" />
                    <SPLIT distance="150" swimtime="00:01:42.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21819" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="21847" number="2" />
                    <RELAYPOSITION athleteid="21882" number="3" />
                    <RELAYPOSITION athleteid="21861" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="505815" nation="POL" region="WIE" clubid="21769" name="Tm Barracuda Kalisz">
          <CONTACT city="KALISZ" email="GALCZYNSKIWOJ@OP.PL" name="GAŁCZYŃSKI WOJCIECH" phone="790690666" state="WLKP" zip="62-800" />
          <ATHLETES>
            <ATHLETE birthdate="1984-02-23" firstname="Justyna" gender="F" lastname="Dominiak" nation="POL" athleteid="22910">
              <RESULTS>
                <RESULT eventid="1165" reactiontime="+87" status="OTL" swimtime="00:25:15.25" resultid="22911" heatid="24319" lane="6" entrytime="00:22:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.60" />
                    <SPLIT distance="100" swimtime="00:01:24.78" />
                    <SPLIT distance="150" swimtime="00:02:12.84" />
                    <SPLIT distance="200" swimtime="00:03:02.45" />
                    <SPLIT distance="250" swimtime="00:03:52.97" />
                    <SPLIT distance="300" swimtime="00:04:43.23" />
                    <SPLIT distance="350" swimtime="00:05:33.43" />
                    <SPLIT distance="400" swimtime="00:06:24.92" />
                    <SPLIT distance="450" swimtime="00:07:16.85" />
                    <SPLIT distance="500" swimtime="00:08:07.66" />
                    <SPLIT distance="550" swimtime="00:08:58.50" />
                    <SPLIT distance="600" swimtime="00:09:49.52" />
                    <SPLIT distance="650" swimtime="00:10:40.75" />
                    <SPLIT distance="700" swimtime="00:11:31.58" />
                    <SPLIT distance="750" swimtime="00:12:23.22" />
                    <SPLIT distance="800" swimtime="00:13:13.98" />
                    <SPLIT distance="850" swimtime="00:14:05.99" />
                    <SPLIT distance="900" swimtime="00:14:57.53" />
                    <SPLIT distance="950" swimtime="00:15:49.37" />
                    <SPLIT distance="1000" swimtime="00:16:40.76" />
                    <SPLIT distance="1050" swimtime="00:17:33.07" />
                    <SPLIT distance="1100" swimtime="00:18:24.53" />
                    <SPLIT distance="1150" swimtime="00:19:15.98" />
                    <SPLIT distance="1200" swimtime="00:20:07.42" />
                    <SPLIT distance="1250" swimtime="00:20:59.19" />
                    <SPLIT distance="1300" swimtime="00:21:50.47" />
                    <SPLIT distance="1350" swimtime="00:22:42.30" />
                    <SPLIT distance="1400" swimtime="00:23:32.82" />
                    <SPLIT distance="1450" swimtime="00:24:24.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="238" reactiontime="+49" swimtime="00:03:44.45" resultid="22912" heatid="24340" lane="0" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.25" />
                    <SPLIT distance="100" swimtime="00:01:44.35" />
                    <SPLIT distance="150" swimtime="00:02:43.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" status="DNS" swimtime="00:00:00.00" resultid="22913" heatid="24350" lane="6" entrytime="00:01:22.00" />
                <RESULT eventid="1388" points="248" reactiontime="+83" swimtime="00:01:42.04" resultid="22914" heatid="24377" lane="5" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="250" reactiontime="+82" swimtime="00:02:59.11" resultid="22915" heatid="24412" lane="5" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-04-07" firstname="Arkadiusz" gender="M" lastname="Figiel" nation="POL" athleteid="22892">
              <RESULTS>
                <RESULT eventid="1079" points="147" reactiontime="+105" swimtime="00:00:39.55" resultid="22893" heatid="24282" lane="5" />
                <RESULT eventid="1113" points="66" reactiontime="+100" swimtime="00:04:41.13" resultid="22894" heatid="24301" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.12" />
                    <SPLIT distance="100" swimtime="00:02:26.56" />
                    <SPLIT distance="150" swimtime="00:03:42.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="79" swimtime="00:00:55.93" resultid="22895" heatid="24328" lane="5" />
                <RESULT comment="K6 - Pływak wykonał nierównoczesne ruchy ramion. (Time: 10:08)" eventid="1239" reactiontime="+61" status="DSQ" swimtime="00:04:23.43" resultid="22896" heatid="24341" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.25" />
                    <SPLIT distance="100" swimtime="00:02:03.52" />
                    <SPLIT distance="150" swimtime="00:03:13.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="118" reactiontime="+83" swimtime="00:01:56.41" resultid="22897" heatid="24381" lane="8" entrytime="00:01:55.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="78" swimtime="00:03:58.65" resultid="22898" heatid="24416" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.81" />
                    <SPLIT distance="100" swimtime="00:01:51.17" />
                    <SPLIT distance="150" swimtime="00:02:59.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="142" reactiontime="+76" swimtime="00:00:49.67" resultid="23858" heatid="24459" lane="2" />
                <RESULT eventid="1744" points="82" reactiontime="+50" swimtime="00:08:25.05" resultid="23859" heatid="24474" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:53.47" />
                    <SPLIT distance="200" swimtime="00:04:08.67" />
                    <SPLIT distance="300" swimtime="00:06:22.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-10-29" firstname="Katarzyna" gender="F" lastname="Figiel" nation="POL" athleteid="22899">
              <RESULTS>
                <RESULT eventid="1062" points="69" swimtime="00:00:57.44" resultid="22900" heatid="24275" lane="6" />
                <RESULT eventid="1222" points="112" swimtime="00:04:48.11" resultid="22901" heatid="24337" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.73" />
                    <SPLIT distance="100" swimtime="00:02:21.36" />
                    <SPLIT distance="150" swimtime="00:03:35.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="45" swimtime="00:02:25.13" resultid="22902" heatid="24348" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="97" swimtime="00:02:19.14" resultid="22903" heatid="24375" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="86" swimtime="00:01:06.51" resultid="22904" heatid="24454" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-11-02" firstname="Anna" gender="F" lastname="Gałczyńska" nation="POL" athleteid="22905">
              <RESULTS>
                <RESULT eventid="1187" points="52" swimtime="00:01:12.41" resultid="22906" heatid="24323" lane="2" />
                <RESULT eventid="1388" points="88" reactiontime="+74" swimtime="00:02:23.94" resultid="22907" heatid="24376" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="43" reactiontime="+129" swimtime="00:02:44.76" resultid="22908" heatid="24399" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="76" reactiontime="+74" swimtime="00:01:09.40" resultid="22909" heatid="24454" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-09-30" firstname="Magdalena" gender="F" lastname="Kolera" nation="POL" athleteid="22881">
              <RESULTS>
                <RESULT eventid="1062" points="246" reactiontime="+106" swimtime="00:00:37.75" resultid="22882" heatid="24277" lane="5" entrytime="00:00:38.20" />
                <RESULT eventid="1187" points="236" swimtime="00:00:43.73" resultid="22883" heatid="24325" lane="7" entrytime="00:00:44.00" />
                <RESULT eventid="1457" points="208" reactiontime="+89" swimtime="00:01:37.87" resultid="22884" heatid="24400" lane="5" entrytime="00:01:36.00" />
                <RESULT eventid="1630" points="190" reactiontime="+139" swimtime="00:03:35.68" resultid="22885" heatid="24443" lane="4" entrytime="00:03:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.72" />
                    <SPLIT distance="100" swimtime="00:01:47.35" />
                    <SPLIT distance="150" swimtime="00:02:43.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="22886" heatid="24470" lane="5" entrytime="00:08:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-04-12" firstname="Karolina" gender="F" lastname="Radomska" nation="POL" athleteid="22922">
              <RESULTS>
                <RESULT eventid="1062" points="268" reactiontime="+125" swimtime="00:00:36.69" resultid="22923" heatid="24275" lane="5" />
                <RESULT eventid="1256" points="232" reactiontime="+87" swimtime="00:01:24.09" resultid="22924" heatid="24347" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="194" reactiontime="+89" swimtime="00:03:15.12" resultid="22925" heatid="24409" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.65" />
                    <SPLIT distance="100" swimtime="00:01:32.48" />
                    <SPLIT distance="150" swimtime="00:02:25.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="174" reactiontime="+104" swimtime="00:07:02.79" resultid="22926" heatid="24469" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.44" />
                    <SPLIT distance="100" swimtime="00:01:35.12" />
                    <SPLIT distance="150" swimtime="00:02:29.04" />
                    <SPLIT distance="200" swimtime="00:03:23.08" />
                    <SPLIT distance="250" swimtime="00:04:18.48" />
                    <SPLIT distance="300" swimtime="00:05:14.63" />
                    <SPLIT distance="350" swimtime="00:06:11.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-06-27" firstname="Małgorzata" gender="F" lastname="Rembowska-Świeboda" nation="POL" athleteid="22887">
              <RESULTS>
                <RESULT eventid="1062" points="375" reactiontime="+79" swimtime="00:00:32.81" resultid="22888" heatid="24279" lane="5" entrytime="00:00:32.50" />
                <RESULT eventid="1187" points="357" swimtime="00:00:38.11" resultid="22889" heatid="24326" lane="3" entrytime="00:00:38.00" />
                <RESULT eventid="1256" points="332" reactiontime="+63" swimtime="00:01:14.65" resultid="22890" heatid="24351" lane="7" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="342" swimtime="00:01:22.88" resultid="22891" heatid="24402" lane="9" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-11" firstname="Patrycja" gender="F" lastname="Rupa" nation="POL" athleteid="22916">
              <RESULTS>
                <RESULT eventid="1062" points="416" reactiontime="+81" swimtime="00:00:31.69" resultid="22917" heatid="24275" lane="3" />
                <RESULT eventid="1147" status="DNS" swimtime="00:00:00.00" resultid="22918" heatid="24311" lane="4" entrytime="00:12:00.00" />
                <RESULT eventid="1187" points="467" swimtime="00:00:34.86" resultid="22919" heatid="24327" lane="6" entrytime="00:00:33.55" />
                <RESULT eventid="1457" points="453" swimtime="00:01:15.49" resultid="22920" heatid="24402" lane="6" entrytime="00:01:12.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="396" reactiontime="+67" swimtime="00:02:48.82" resultid="22921" heatid="24445" lane="2" entrytime="00:02:42.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.61" />
                    <SPLIT distance="100" swimtime="00:01:22.04" />
                    <SPLIT distance="150" swimtime="00:02:05.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1525" points="318" reactiontime="+78" swimtime="00:02:21.25" resultid="22927" heatid="24425" lane="2" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.37" />
                    <SPLIT distance="100" swimtime="00:01:12.10" />
                    <SPLIT distance="150" swimtime="00:01:49.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22910" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="22922" number="2" />
                    <RELAYPOSITION athleteid="22881" number="3" reactiontime="+14" />
                    <RELAYPOSITION athleteid="22887" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1358" points="163" reactiontime="+114" swimtime="00:03:14.38" resultid="22928" heatid="24372" lane="2" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.89" />
                    <SPLIT distance="150" swimtime="00:02:40.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22905" number="1" reactiontime="+114" />
                    <RELAYPOSITION athleteid="22910" number="2" />
                    <RELAYPOSITION athleteid="22887" number="3" />
                    <RELAYPOSITION athleteid="22922" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="TMT" nation="POL" region="KUJ" clubid="20479" name="Toruń Multisport Team">
          <CONTACT city="Toruń" email="g.arentewicz@onet.pl" name="Arentewicz" phone="535763476" state="KUJ-P" street="Rydygiera 42A/19" zip="87-100" />
          <ATHLETES>
            <ATHLETE birthdate="1949-08-24" firstname="Jan" gender="M" lastname="Bantkowski" nation="POL" athleteid="20512">
              <RESULTS>
                <RESULT eventid="1113" points="41" reactiontime="+126" swimtime="00:05:28.37" resultid="20513" heatid="24301" lane="8" entrytime="00:04:58.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:04:29.39" />
                    <SPLIT distance="100" swimtime="00:02:54.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14189" reactiontime="+143" status="OTL" swimtime="00:21:02.27" resultid="20514" heatid="24314" lane="0" entrytime="00:18:20.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.50" />
                    <SPLIT distance="100" swimtime="00:02:36.34" />
                    <SPLIT distance="150" swimtime="00:03:57.84" />
                    <SPLIT distance="200" swimtime="00:05:20.64" />
                    <SPLIT distance="250" swimtime="00:06:41.71" />
                    <SPLIT distance="300" swimtime="00:08:01.91" />
                    <SPLIT distance="350" swimtime="00:09:22.26" />
                    <SPLIT distance="400" swimtime="00:10:43.21" />
                    <SPLIT distance="450" swimtime="00:12:03.84" />
                    <SPLIT distance="500" swimtime="00:13:24.21" />
                    <SPLIT distance="550" swimtime="00:14:45.16" />
                    <SPLIT distance="650" swimtime="00:17:29.57" />
                    <SPLIT distance="700" swimtime="00:18:49.60" />
                    <SPLIT distance="750" swimtime="00:20:02.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="34" swimtime="00:01:13.99" resultid="20515" heatid="24329" lane="1" entrytime="00:01:01.78" />
                <RESULT eventid="1341" points="23" reactiontime="+104" swimtime="00:06:27.05" resultid="20516" heatid="24368" lane="3" entrytime="00:05:45.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:27.46" />
                    <SPLIT distance="100" swimtime="00:03:09.82" />
                    <SPLIT distance="150" swimtime="00:04:52.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="52" reactiontime="+86" swimtime="00:04:32.81" resultid="20517" heatid="24416" lane="6" entrytime="00:03:59.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.97" />
                    <SPLIT distance="100" swimtime="00:02:15.25" />
                    <SPLIT distance="150" swimtime="00:03:28.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="40" reactiontime="+94" swimtime="00:11:48.95" resultid="20518" heatid="24430" lane="8" entrytime="00:10:48.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.09" />
                    <SPLIT distance="100" swimtime="00:06:17.06" />
                    <SPLIT distance="150" swimtime="00:04:41.15" />
                    <SPLIT distance="250" swimtime="00:07:56.18" />
                    <SPLIT distance="300" swimtime="00:09:35.24" />
                    <SPLIT distance="350" swimtime="00:10:46.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="26" reactiontime="+94" swimtime="00:02:48.12" resultid="20519" heatid="24437" lane="6" entrytime="00:02:34.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="46" reactiontime="+95" swimtime="00:10:13.36" resultid="20520" heatid="24475" lane="8" entrytime="00:08:59.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.70" />
                    <SPLIT distance="150" swimtime="00:03:53.40" />
                    <SPLIT distance="250" swimtime="00:06:34.13" />
                    <SPLIT distance="350" swimtime="00:09:11.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-28" firstname="Marek" gender="M" lastname="Brożyna" nation="POL" athleteid="20504">
              <RESULTS>
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="20505" heatid="24305" lane="6" entrytime="00:02:41.53" />
                <RESULT eventid="1205" points="338" swimtime="00:00:34.43" resultid="20506" heatid="24334" lane="0" entrytime="00:00:33.78" />
                <RESULT eventid="1273" points="386" reactiontime="+80" swimtime="00:01:04.38" resultid="20507" heatid="24360" lane="3" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="371" reactiontime="+74" swimtime="00:01:12.11" resultid="20508" heatid="24407" lane="2" entrytime="00:01:12.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="334" swimtime="00:05:51.13" resultid="20509" heatid="24432" lane="3" entrytime="00:05:44.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.03" />
                    <SPLIT distance="100" swimtime="00:01:19.56" />
                    <SPLIT distance="150" swimtime="00:02:04.11" />
                    <SPLIT distance="200" swimtime="00:02:47.30" />
                    <SPLIT distance="250" swimtime="00:03:39.14" />
                    <SPLIT distance="300" swimtime="00:04:31.45" />
                    <SPLIT distance="350" swimtime="00:05:10.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="367" swimtime="00:02:36.27" resultid="20510" heatid="24451" lane="8" entrytime="00:02:37.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                    <SPLIT distance="100" swimtime="00:01:15.12" />
                    <SPLIT distance="150" swimtime="00:01:56.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="344" reactiontime="+43" swimtime="00:05:14.06" resultid="20511" heatid="24480" lane="2" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                    <SPLIT distance="100" swimtime="00:01:11.99" />
                    <SPLIT distance="150" swimtime="00:01:51.95" />
                    <SPLIT distance="200" swimtime="00:02:32.66" />
                    <SPLIT distance="250" swimtime="00:03:13.33" />
                    <SPLIT distance="300" swimtime="00:03:54.77" />
                    <SPLIT distance="350" swimtime="00:04:35.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-10-28" firstname="Andrzej" gender="M" lastname="Gołembiewski" nation="POL" athleteid="20497">
              <RESULTS>
                <RESULT eventid="14189" points="389" reactiontime="+84" swimtime="00:10:18.89" resultid="20498" heatid="24317" lane="2" entrytime="00:10:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:10.15" />
                    <SPLIT distance="150" swimtime="00:01:48.46" />
                    <SPLIT distance="200" swimtime="00:02:27.28" />
                    <SPLIT distance="250" swimtime="00:03:06.32" />
                    <SPLIT distance="300" swimtime="00:03:45.72" />
                    <SPLIT distance="350" swimtime="00:04:25.41" />
                    <SPLIT distance="400" swimtime="00:05:05.26" />
                    <SPLIT distance="450" swimtime="00:05:45.39" />
                    <SPLIT distance="500" swimtime="00:06:25.39" />
                    <SPLIT distance="550" swimtime="00:07:05.04" />
                    <SPLIT distance="600" swimtime="00:07:44.70" />
                    <SPLIT distance="650" swimtime="00:08:24.28" />
                    <SPLIT distance="700" swimtime="00:09:03.57" />
                    <SPLIT distance="750" swimtime="00:09:42.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="439" reactiontime="+43" swimtime="00:02:46.64" resultid="20499" heatid="24346" lane="1" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.85" />
                    <SPLIT distance="100" swimtime="00:01:22.19" />
                    <SPLIT distance="150" swimtime="00:02:05.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="489" reactiontime="+76" swimtime="00:01:12.44" resultid="20500" heatid="24385" lane="8" entrytime="00:01:10.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="20501" heatid="24423" lane="2" entrytime="00:02:11.00" />
                <RESULT eventid="1681" points="499" swimtime="00:00:32.71" resultid="20502" heatid="24466" lane="9" entrytime="00:00:32.00" />
                <RESULT eventid="1744" points="435" reactiontime="+71" swimtime="00:04:50.33" resultid="20503" heatid="24482" lane="8" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                    <SPLIT distance="100" swimtime="00:01:06.22" />
                    <SPLIT distance="150" swimtime="00:01:41.91" />
                    <SPLIT distance="200" swimtime="00:02:18.78" />
                    <SPLIT distance="250" swimtime="00:02:56.03" />
                    <SPLIT distance="300" swimtime="00:03:34.58" />
                    <SPLIT distance="350" swimtime="00:04:13.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-04-23" firstname="Krzysztof" gender="M" lastname="Lietz" nation="POL" athleteid="20489">
              <RESULTS>
                <RESULT eventid="1079" points="242" reactiontime="+88" swimtime="00:00:33.55" resultid="20490" heatid="24287" lane="1" entrytime="00:00:33.20" />
                <RESULT eventid="14189" points="185" reactiontime="+88" swimtime="00:13:12.13" resultid="20491" heatid="24315" lane="1" entrytime="00:12:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.11" />
                    <SPLIT distance="100" swimtime="00:01:31.24" />
                    <SPLIT distance="250" swimtime="00:04:01.83" />
                    <SPLIT distance="300" swimtime="00:04:51.54" />
                    <SPLIT distance="350" swimtime="00:05:42.65" />
                    <SPLIT distance="400" swimtime="00:06:33.33" />
                    <SPLIT distance="450" swimtime="00:07:24.47" />
                    <SPLIT distance="500" swimtime="00:08:14.17" />
                    <SPLIT distance="550" swimtime="00:09:05.55" />
                    <SPLIT distance="600" swimtime="00:09:55.69" />
                    <SPLIT distance="650" swimtime="00:10:47.60" />
                    <SPLIT distance="700" swimtime="00:11:37.45" />
                    <SPLIT distance="750" swimtime="00:12:27.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="229" reactiontime="+71" swimtime="00:01:16.61" resultid="20492" heatid="24357" lane="3" entrytime="00:01:14.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="204" swimtime="00:00:37.77" resultid="20493" heatid="24392" lane="7" entrytime="00:00:37.50" />
                <RESULT eventid="1508" points="191" reactiontime="+84" swimtime="00:02:56.98" resultid="20494" heatid="24418" lane="4" entrytime="00:02:57.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.89" />
                    <SPLIT distance="100" swimtime="00:01:29.35" />
                    <SPLIT distance="150" swimtime="00:02:15.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="20495" heatid="24439" lane="1" entrytime="00:01:32.00" />
                <RESULT eventid="1744" points="189" reactiontime="+78" swimtime="00:06:22.84" resultid="20496" heatid="24477" lane="4" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.93" />
                    <SPLIT distance="100" swimtime="00:01:33.18" />
                    <SPLIT distance="150" swimtime="00:02:23.43" />
                    <SPLIT distance="200" swimtime="00:03:12.67" />
                    <SPLIT distance="250" swimtime="00:04:02.91" />
                    <SPLIT distance="300" swimtime="00:04:51.01" />
                    <SPLIT distance="350" swimtime="00:05:38.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-06-29" firstname="Lucyna" gender="F" lastname="Serożyńska" nation="POL" athleteid="20480">
              <RESULTS>
                <RESULT eventid="1062" points="72" reactiontime="+145" swimtime="00:00:56.70" resultid="20481" heatid="24276" lane="7" entrytime="00:01:01.00" />
                <RESULT eventid="1147" points="91" reactiontime="+112" swimtime="00:17:56.60" resultid="20482" heatid="24310" lane="2" entrytime="00:18:29.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:58.65" />
                    <SPLIT distance="150" swimtime="00:03:05.53" />
                    <SPLIT distance="250" swimtime="00:07:41.78" />
                    <SPLIT distance="300" swimtime="00:06:32.37" />
                    <SPLIT distance="350" swimtime="00:10:03.52" />
                    <SPLIT distance="400" swimtime="00:08:53.96" />
                    <SPLIT distance="450" swimtime="00:12:21.51" />
                    <SPLIT distance="500" swimtime="00:11:14.08" />
                    <SPLIT distance="550" swimtime="00:14:39.36" />
                    <SPLIT distance="600" swimtime="00:13:29.26" />
                    <SPLIT distance="650" swimtime="00:16:52.94" />
                    <SPLIT distance="700" swimtime="00:15:45.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="78" swimtime="00:01:03.20" resultid="20483" heatid="24324" lane="9" entrytime="00:01:03.00" />
                <RESULT eventid="1256" points="95" reactiontime="+87" swimtime="00:01:53.10" resultid="20484" heatid="24348" lane="6" entrytime="00:02:02.00" />
                <RESULT eventid="1457" points="85" reactiontime="+95" swimtime="00:02:11.91" resultid="20485" heatid="24400" lane="1" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="20486" heatid="24410" lane="1" entrytime="00:04:25.00" />
                <RESULT eventid="1630" points="88" reactiontime="+80" swimtime="00:04:38.46" resultid="20487" heatid="24443" lane="2" entrytime="00:04:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.68" />
                    <SPLIT distance="100" swimtime="00:02:16.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="88" reactiontime="+120" swimtime="00:08:51.24" resultid="20488" heatid="24470" lane="8" entrytime="00:09:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:03:12.48" />
                    <SPLIT distance="250" swimtime="00:05:31.63" />
                    <SPLIT distance="300" swimtime="00:06:39.63" />
                    <SPLIT distance="350" swimtime="00:07:46.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="OLPOZ" nation="POL" region="WIE" clubid="21456" name="TS Olimpia Poznań">
          <CONTACT name="Pietraszewski" phone="501 648 415" />
          <ATHLETES>
            <ATHLETE birthdate="1944-01-01" firstname="Jacek" gender="M" lastname="Lesiński" nation="POL" athleteid="21457">
              <RESULTS>
                <RESULT eventid="1079" points="133" reactiontime="+112" swimtime="00:00:40.89" resultid="21458" heatid="24284" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="1113" points="113" reactiontime="+110" swimtime="00:03:55.30" resultid="21459" heatid="24302" lane="6" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.78" />
                    <SPLIT distance="100" swimtime="00:01:55.27" />
                    <SPLIT distance="150" swimtime="00:03:01.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="135" swimtime="00:00:46.73" resultid="21460" heatid="24330" lane="3" entrytime="00:00:46.00" />
                <RESULT eventid="1273" points="130" reactiontime="+107" swimtime="00:01:32.59" resultid="21461" heatid="24355" lane="4" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="112" reactiontime="+84" swimtime="00:01:47.40" resultid="21463" heatid="24404" lane="1" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="112" swimtime="00:03:51.80" resultid="21464" heatid="24448" lane="1" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.60" />
                    <SPLIT distance="100" swimtime="00:03:55.19" />
                    <SPLIT distance="150" swimtime="00:02:52.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-01-01" firstname="Jacek" gender="M" lastname="Matyszczak" nation="POL" athleteid="21474">
              <RESULTS>
                <RESULT eventid="1079" points="378" reactiontime="+88" swimtime="00:00:28.91" resultid="21475" heatid="24291" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="14189" points="202" reactiontime="+104" swimtime="00:12:50.26" resultid="21476" heatid="24315" lane="3" entrytime="00:12:15.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.17" />
                    <SPLIT distance="200" swimtime="00:02:48.44" />
                    <SPLIT distance="250" swimtime="00:03:33.79" />
                    <SPLIT distance="300" swimtime="00:04:19.12" />
                    <SPLIT distance="350" swimtime="00:05:04.67" />
                    <SPLIT distance="400" swimtime="00:05:51.84" />
                    <SPLIT distance="450" swimtime="00:06:39.09" />
                    <SPLIT distance="500" swimtime="00:07:26.57" />
                    <SPLIT distance="550" swimtime="00:08:23.60" />
                    <SPLIT distance="600" swimtime="00:09:18.93" />
                    <SPLIT distance="650" swimtime="00:10:16.95" />
                    <SPLIT distance="700" swimtime="00:11:18.85" />
                    <SPLIT distance="750" swimtime="00:12:05.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="220" swimtime="00:00:39.75" resultid="21477" heatid="24332" lane="3" entrytime="00:00:38.50" />
                <RESULT eventid="1273" points="347" swimtime="00:01:06.72" resultid="21478" heatid="24360" lane="7" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="21479" heatid="24393" lane="4" entrytime="00:00:34.00" />
                <RESULT eventid="1508" points="274" swimtime="00:02:36.89" resultid="21480" heatid="24421" lane="9" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                    <SPLIT distance="100" swimtime="00:01:13.01" />
                    <SPLIT distance="150" swimtime="00:01:54.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="166" reactiontime="+89" swimtime="00:03:23.60" resultid="21481" heatid="24449" lane="0" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.03" />
                    <SPLIT distance="100" swimtime="00:01:40.06" />
                    <SPLIT distance="150" swimtime="00:02:33.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="244" reactiontime="+101" swimtime="00:05:51.94" resultid="21482" heatid="24479" lane="3" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                    <SPLIT distance="100" swimtime="00:01:19.47" />
                    <SPLIT distance="300" swimtime="00:04:22.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Zbigniew" gender="M" lastname="Pietraszewski" nation="POL" athleteid="21466">
              <RESULTS>
                <RESULT eventid="1113" points="194" reactiontime="+104" swimtime="00:03:16.90" resultid="21467" heatid="24303" lane="3" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.25" />
                    <SPLIT distance="100" swimtime="00:01:36.29" />
                    <SPLIT distance="150" swimtime="00:02:31.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14189" points="190" reactiontime="+99" swimtime="00:13:06.19" resultid="21468" heatid="24315" lane="8" entrytime="00:13:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.69" />
                    <SPLIT distance="100" swimtime="00:01:31.66" />
                    <SPLIT distance="150" swimtime="00:02:22.17" />
                    <SPLIT distance="200" swimtime="00:03:12.81" />
                    <SPLIT distance="250" swimtime="00:04:03.79" />
                    <SPLIT distance="300" swimtime="00:04:54.66" />
                    <SPLIT distance="350" swimtime="00:05:45.81" />
                    <SPLIT distance="400" swimtime="00:06:36.64" />
                    <SPLIT distance="450" swimtime="00:07:26.91" />
                    <SPLIT distance="500" swimtime="00:08:17.10" />
                    <SPLIT distance="550" swimtime="00:09:06.30" />
                    <SPLIT distance="600" swimtime="00:09:55.60" />
                    <SPLIT distance="650" swimtime="00:10:44.67" />
                    <SPLIT distance="700" swimtime="00:11:34.05" />
                    <SPLIT distance="750" swimtime="00:12:22.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="170" swimtime="00:00:43.26" resultid="21469" heatid="24331" lane="4" entrytime="00:00:41.00" />
                <RESULT eventid="1474" points="179" reactiontime="+87" swimtime="00:01:31.95" resultid="21470" heatid="24405" lane="2" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="193" reactiontime="+70" swimtime="00:07:01.41" resultid="21471" heatid="24431" lane="4" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.83" />
                    <SPLIT distance="100" swimtime="00:01:50.67" />
                    <SPLIT distance="150" swimtime="00:02:42.76" />
                    <SPLIT distance="200" swimtime="00:03:34.34" />
                    <SPLIT distance="250" swimtime="00:04:31.55" />
                    <SPLIT distance="300" swimtime="00:05:28.42" />
                    <SPLIT distance="350" swimtime="00:06:15.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="196" reactiontime="+89" swimtime="00:03:12.56" resultid="21472" heatid="24449" lane="3" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.37" />
                    <SPLIT distance="100" swimtime="00:01:35.53" />
                    <SPLIT distance="150" swimtime="00:02:24.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="21473" heatid="24478" lane="9" entrytime="00:06:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Maria" gender="F" lastname="Łutowicz" nation="POL" athleteid="21483">
              <RESULTS>
                <RESULT eventid="1062" points="199" reactiontime="+96" swimtime="00:00:40.52" resultid="21484" heatid="24277" lane="8" entrytime="00:00:43.00" />
                <RESULT eventid="1187" points="108" swimtime="00:00:56.79" resultid="21485" heatid="24324" lane="3" entrytime="00:00:53.00" />
                <RESULT eventid="1256" points="154" reactiontime="+78" swimtime="00:01:36.43" resultid="21486" heatid="24349" lane="6" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="98" reactiontime="+99" swimtime="00:00:52.96" resultid="21487" heatid="24386" lane="3" entrytime="00:00:54.00" />
                <RESULT eventid="1491" points="131" reactiontime="+77" swimtime="00:03:41.99" resultid="21488" heatid="24411" lane="1" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.48" />
                    <SPLIT distance="100" swimtime="00:01:49.31" />
                    <SPLIT distance="150" swimtime="00:02:47.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="109" reactiontime="+80" swimtime="00:04:19.31" resultid="21489" heatid="24443" lane="3" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.46" />
                    <SPLIT distance="100" swimtime="00:02:10.89" />
                    <SPLIT distance="150" swimtime="00:03:15.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="145" reactiontime="+83" swimtime="00:07:29.19" resultid="21490" heatid="24471" lane="1" entrytime="00:07:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.01" />
                    <SPLIT distance="100" swimtime="00:01:49.20" />
                    <SPLIT distance="150" swimtime="00:02:48.61" />
                    <SPLIT distance="200" swimtime="00:03:46.13" />
                    <SPLIT distance="250" swimtime="00:04:43.84" />
                    <SPLIT distance="300" swimtime="00:05:41.19" />
                    <SPLIT distance="350" swimtime="00:06:37.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01414" nation="POL" region="WA" clubid="20657" name="UKS Delfin Legionowo">
          <CONTACT city="LEGIONOWO" email="delfin-trener@wp.pl" internet="www.delfinlegionowo.pl" name="RAFAŁ PERL" phone="0-601 436 700" state="MAZ" street="KRÓLOWEJ JADWIGI 11" zip="05-120" />
          <ATHLETES>
            <ATHLETE birthdate="1996-06-07" firstname="Michał" gender="M" lastname="Perl" nation="POL" license="101414700068" athleteid="21424">
              <RESULTS>
                <RESULT eventid="14189" reactiontime="+79" status="OTL" swimtime="00:11:23.02" resultid="21425" heatid="24317" lane="8" entrytime="00:10:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                    <SPLIT distance="100" swimtime="00:01:12.26" />
                    <SPLIT distance="150" swimtime="00:01:51.90" />
                    <SPLIT distance="250" swimtime="00:03:16.41" />
                    <SPLIT distance="450" swimtime="00:06:12.13" />
                    <SPLIT distance="650" swimtime="00:09:11.26" />
                    <SPLIT distance="750" swimtime="00:10:41.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="470" reactiontime="+82" swimtime="00:02:42.87" resultid="21426" heatid="24346" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.12" />
                    <SPLIT distance="100" swimtime="00:01:16.86" />
                    <SPLIT distance="150" swimtime="00:01:59.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1079" points="640" reactiontime="+73" swimtime="00:00:24.26" resultid="21427" heatid="24296" lane="4" entrytime="00:00:23.00" />
                <RESULT eventid="1273" points="567" swimtime="00:00:56.66" resultid="21428" heatid="24365" lane="5" entrytime="00:00:54.00" />
                <RESULT eventid="1406" points="531" swimtime="00:01:10.48" resultid="21429" heatid="24385" lane="5" entrytime="00:01:06.00" />
                <RESULT eventid="1440" points="554" swimtime="00:00:27.10" resultid="21430" heatid="24398" lane="2" entrytime="00:00:26.00" />
                <RESULT eventid="1681" points="660" swimtime="00:00:29.79" resultid="21431" heatid="24466" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="1744" points="270" reactiontime="+69" swimtime="00:05:40.29" resultid="21432" heatid="24480" lane="7" entrytime="00:05:14.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.29" />
                    <SPLIT distance="100" swimtime="00:01:15.39" />
                    <SPLIT distance="150" swimtime="00:01:57.44" />
                    <SPLIT distance="200" swimtime="00:02:40.63" />
                    <SPLIT distance="250" swimtime="00:03:25.03" />
                    <SPLIT distance="300" swimtime="00:04:10.71" />
                    <SPLIT distance="350" swimtime="00:04:56.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-05-19" firstname="Dawid" gender="M" lastname="Szulich" nation="POL" license="101414700035" athleteid="21433">
              <RESULTS>
                <RESULT eventid="1681" points="672" reactiontime="+68" swimtime="00:00:29.62" resultid="21434" heatid="24466" lane="3" entrytime="00:00:29.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-31" firstname="Joanna" gender="F" lastname="Żbikowska" nation="POL" athleteid="21440">
              <RESULTS>
                <RESULT eventid="1062" points="476" reactiontime="+73" swimtime="00:00:30.31" resultid="21441" heatid="24280" lane="7" entrytime="00:00:31.00" />
                <RESULT eventid="1096" points="348" reactiontime="+79" swimtime="00:02:59.26" resultid="21442" heatid="24299" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.76" />
                    <SPLIT distance="100" swimtime="00:01:23.45" />
                    <SPLIT distance="150" swimtime="00:02:12.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="421" swimtime="00:01:08.95" resultid="21443" heatid="24351" lane="5" entrytime="00:01:15.00" />
                <RESULT eventid="1388" points="404" reactiontime="+70" swimtime="00:01:26.69" resultid="21444" heatid="24379" lane="7" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="384" swimtime="00:00:33.61" resultid="21445" heatid="24388" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1664" points="453" swimtime="00:00:38.28" resultid="21446" heatid="24458" lane="3" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-06-23" firstname="Krzysztof" gender="M" lastname="Żbikowski" nation="POL" athleteid="21435">
              <RESULTS>
                <RESULT eventid="1079" points="425" reactiontime="+75" swimtime="00:00:27.80" resultid="21436" heatid="24295" lane="1" entrytime="00:00:26.00" />
                <RESULT eventid="1273" points="441" swimtime="00:01:01.60" resultid="21437" heatid="24365" lane="9" entrytime="00:00:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="560" swimtime="00:01:09.26" resultid="21438" heatid="24385" lane="2" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="587" swimtime="00:00:30.99" resultid="21439" heatid="24466" lane="1" entrytime="00:00:30.15" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00408" nation="POL" region="RZ" clubid="21397" name="UKS Delfin Masters Tarnobrzeg">
          <CONTACT city="TARNOBRZEG" email="piotr.michalik@i-bs.pl" name="MICHALIK ANGELIKA" state="PODKA" street="SKALNA GÓRA 8/21" street2="TARNOBRZEG" zip="39-400" />
          <ATHLETES>
            <ATHLETE birthdate="1971-01-14" firstname="Piotr" gender="M" lastname="Darowski" nation="POL" athleteid="21414">
              <RESULTS>
                <RESULT eventid="1113" points="416" reactiontime="+75" swimtime="00:02:32.70" resultid="21415" heatid="24305" lane="4" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                    <SPLIT distance="100" swimtime="00:01:13.24" />
                    <SPLIT distance="150" swimtime="00:01:57.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="431" swimtime="00:02:47.69" resultid="21416" heatid="24346" lane="9" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                    <SPLIT distance="100" swimtime="00:01:19.40" />
                    <SPLIT distance="150" swimtime="00:02:03.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="414" swimtime="00:01:16.56" resultid="21417" heatid="24384" lane="2" entrytime="00:01:19.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="359" swimtime="00:05:43.00" resultid="21418" heatid="24432" lane="1" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.53" />
                    <SPLIT distance="100" swimtime="00:01:16.79" />
                    <SPLIT distance="150" swimtime="00:02:04.24" />
                    <SPLIT distance="200" swimtime="00:02:51.32" />
                    <SPLIT distance="250" swimtime="00:03:38.99" />
                    <SPLIT distance="300" swimtime="00:04:25.29" />
                    <SPLIT distance="350" swimtime="00:05:05.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="419" swimtime="00:00:34.66" resultid="21419" heatid="24465" lane="1" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-03-14" firstname="Maciej" gender="M" lastname="Kunicki" nation="POL" athleteid="20288">
              <RESULTS>
                <RESULT eventid="1113" points="271" reactiontime="+94" swimtime="00:02:55.98" resultid="20289" heatid="24304" lane="3" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                    <SPLIT distance="100" swimtime="00:01:23.58" />
                    <SPLIT distance="150" swimtime="00:02:18.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="210" reactiontime="+44" swimtime="00:03:07.41" resultid="20290" heatid="24370" lane="6" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.18" />
                    <SPLIT distance="100" swimtime="00:01:28.59" />
                    <SPLIT distance="150" swimtime="00:02:18.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="309" reactiontime="+54" swimtime="00:00:32.92" resultid="20291" heatid="24394" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="1613" points="244" reactiontime="+45" swimtime="00:01:19.69" resultid="20292" heatid="24439" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-12" firstname="Maciej" gender="M" lastname="Płaneta" nation="POL" athleteid="21398">
              <RESULTS>
                <RESULT eventid="1079" points="303" reactiontime="+89" swimtime="00:00:31.10" resultid="21399" heatid="24289" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="14207" points="267" reactiontime="+81" swimtime="00:22:32.36" resultid="21400" heatid="24321" lane="6" entrytime="00:23:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                    <SPLIT distance="100" swimtime="00:01:21.26" />
                    <SPLIT distance="150" swimtime="00:02:04.75" />
                    <SPLIT distance="200" swimtime="00:02:49.66" />
                    <SPLIT distance="250" swimtime="00:03:35.65" />
                    <SPLIT distance="300" swimtime="00:04:21.51" />
                    <SPLIT distance="350" swimtime="00:05:07.48" />
                    <SPLIT distance="400" swimtime="00:05:52.56" />
                    <SPLIT distance="450" swimtime="00:06:38.67" />
                    <SPLIT distance="500" swimtime="00:07:24.23" />
                    <SPLIT distance="550" swimtime="00:08:09.92" />
                    <SPLIT distance="600" swimtime="00:08:55.38" />
                    <SPLIT distance="650" swimtime="00:09:41.47" />
                    <SPLIT distance="700" swimtime="00:10:26.97" />
                    <SPLIT distance="750" swimtime="00:11:12.44" />
                    <SPLIT distance="800" swimtime="00:11:58.08" />
                    <SPLIT distance="850" swimtime="00:12:43.61" />
                    <SPLIT distance="900" swimtime="00:13:28.89" />
                    <SPLIT distance="950" swimtime="00:14:15.08" />
                    <SPLIT distance="1000" swimtime="00:15:00.60" />
                    <SPLIT distance="1050" swimtime="00:15:46.25" />
                    <SPLIT distance="1100" swimtime="00:16:32.04" />
                    <SPLIT distance="1150" swimtime="00:17:17.30" />
                    <SPLIT distance="1200" swimtime="00:18:02.58" />
                    <SPLIT distance="1250" swimtime="00:18:48.44" />
                    <SPLIT distance="1300" swimtime="00:19:34.53" />
                    <SPLIT distance="1350" swimtime="00:20:20.57" />
                    <SPLIT distance="1400" swimtime="00:21:06.22" />
                    <SPLIT distance="1450" swimtime="00:21:50.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="328" swimtime="00:01:07.97" resultid="21401" heatid="24359" lane="2" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="180" reactiontime="+80" swimtime="00:03:17.41" resultid="21402" heatid="24370" lane="7" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.50" />
                    <SPLIT distance="100" swimtime="00:01:35.13" />
                    <SPLIT distance="150" swimtime="00:02:28.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="215" reactiontime="+77" swimtime="00:01:26.55" resultid="21403" heatid="24405" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="277" reactiontime="+53" swimtime="00:02:36.45" resultid="21404" heatid="24421" lane="0" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                    <SPLIT distance="100" swimtime="00:01:14.86" />
                    <SPLIT distance="150" swimtime="00:01:55.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="218" reactiontime="+78" swimtime="00:03:05.70" resultid="21405" heatid="24450" lane="8" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.83" />
                    <SPLIT distance="100" swimtime="00:01:32.11" />
                    <SPLIT distance="150" swimtime="00:02:20.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="21406" heatid="24480" lane="9" entrytime="00:05:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-03-14" firstname="Katarzyna" gender="F" lastname="Szwagiel" nation="POL" athleteid="21407">
              <RESULTS>
                <RESULT eventid="1096" points="331" reactiontime="+95" swimtime="00:03:02.19" resultid="21408" heatid="24298" lane="3" entrytime="00:03:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.07" />
                    <SPLIT distance="100" swimtime="00:01:28.96" />
                    <SPLIT distance="150" swimtime="00:02:19.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="289" reactiontime="+102" swimtime="00:12:12.61" resultid="21409" heatid="24311" lane="5" entrytime="00:12:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.98" />
                    <SPLIT distance="100" swimtime="00:01:21.62" />
                    <SPLIT distance="150" swimtime="00:02:06.99" />
                    <SPLIT distance="200" swimtime="00:02:53.12" />
                    <SPLIT distance="250" swimtime="00:03:40.33" />
                    <SPLIT distance="300" swimtime="00:04:27.26" />
                    <SPLIT distance="350" swimtime="00:05:13.92" />
                    <SPLIT distance="400" swimtime="00:06:00.62" />
                    <SPLIT distance="450" swimtime="00:06:47.18" />
                    <SPLIT distance="500" swimtime="00:07:33.68" />
                    <SPLIT distance="550" swimtime="00:08:20.80" />
                    <SPLIT distance="600" swimtime="00:09:06.86" />
                    <SPLIT distance="650" swimtime="00:09:53.65" />
                    <SPLIT distance="700" swimtime="00:10:40.25" />
                    <SPLIT distance="750" swimtime="00:11:26.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="353" reactiontime="+52" swimtime="00:02:39.75" resultid="21410" heatid="24413" lane="7" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.32" />
                    <SPLIT distance="100" swimtime="00:01:16.02" />
                    <SPLIT distance="150" swimtime="00:01:58.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1555" points="305" reactiontime="+99" swimtime="00:06:35.70" resultid="21411" heatid="24429" lane="2" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.91" />
                    <SPLIT distance="100" swimtime="00:01:34.30" />
                    <SPLIT distance="150" swimtime="00:02:26.67" />
                    <SPLIT distance="200" swimtime="00:03:18.25" />
                    <SPLIT distance="250" swimtime="00:04:11.87" />
                    <SPLIT distance="300" swimtime="00:05:06.56" />
                    <SPLIT distance="350" swimtime="00:05:52.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1595" points="236" swimtime="00:01:29.71" resultid="21412" heatid="24436" lane="9" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="310" reactiontime="+85" swimtime="00:05:49.36" resultid="21413" heatid="24472" lane="8" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                    <SPLIT distance="100" swimtime="00:01:21.85" />
                    <SPLIT distance="150" swimtime="00:02:05.36" />
                    <SPLIT distance="200" swimtime="00:02:49.69" />
                    <SPLIT distance="250" swimtime="00:03:34.09" />
                    <SPLIT distance="350" swimtime="00:05:04.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-12-29" firstname="Tomasz" gender="M" lastname="Szwagiel" nation="POL" athleteid="21420">
              <RESULTS>
                <RESULT eventid="1079" points="316" reactiontime="+83" swimtime="00:00:30.67" resultid="21421" heatid="24289" lane="3" entrytime="00:00:30.28" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="322" reactiontime="+102" swimtime="00:02:16.22" resultid="21422" heatid="24374" lane="0" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.01" />
                    <SPLIT distance="100" swimtime="00:01:11.99" />
                    <SPLIT distance="150" swimtime="00:01:45.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21398" number="1" reactiontime="+102" />
                    <RELAYPOSITION athleteid="21414" number="2" />
                    <RELAYPOSITION athleteid="20288" number="3" reactiontime="+11" />
                    <RELAYPOSITION athleteid="21420" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="338" swimtime="00:02:01.72" resultid="21423" heatid="24427" lane="0" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.67" />
                    <SPLIT distance="100" swimtime="00:01:00.66" />
                    <SPLIT distance="150" swimtime="00:01:31.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21414" number="1" />
                    <RELAYPOSITION athleteid="20288" number="2" />
                    <RELAYPOSITION athleteid="21420" number="3" />
                    <RELAYPOSITION athleteid="21398" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00501" nation="POL" region="DOL" clubid="20382" name="UKS Energetyk Zgorzelec">
          <CONTACT city="Zgorzelec" email="biuro@plywanie-zgorzelec.pl" internet="www.plywanie-zgorzelec.pl" name="Kondracki Łukasz" phone="693852488" state="DOL" street="Maratońska" street2="2" zip="59-900" />
          <ATHLETES>
            <ATHLETE birthdate="1948-11-29" firstname="Andrzej" gender="M" lastname="Daszyński" nation="POL" athleteid="20383">
              <RESULTS>
                <RESULT eventid="1113" points="81" reactiontime="+102" swimtime="00:04:23.18" resultid="20384" heatid="24301" lane="4" entrytime="00:04:15.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.75" />
                    <SPLIT distance="100" swimtime="00:02:11.83" />
                    <SPLIT distance="150" swimtime="00:03:26.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14189" points="78" reactiontime="+106" swimtime="00:17:33.74" resultid="20385" heatid="24314" lane="1" entrytime="00:16:46.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.56" />
                    <SPLIT distance="100" swimtime="00:02:04.22" />
                    <SPLIT distance="150" swimtime="00:03:10.60" />
                    <SPLIT distance="200" swimtime="00:04:17.35" />
                    <SPLIT distance="250" swimtime="00:05:24.81" />
                    <SPLIT distance="300" swimtime="00:06:31.07" />
                    <SPLIT distance="350" swimtime="00:07:38.30" />
                    <SPLIT distance="400" swimtime="00:08:45.53" />
                    <SPLIT distance="450" swimtime="00:09:52.89" />
                    <SPLIT distance="500" swimtime="00:10:58.62" />
                    <SPLIT distance="550" swimtime="00:12:06.23" />
                    <SPLIT distance="600" swimtime="00:13:13.85" />
                    <SPLIT distance="650" swimtime="00:14:20.88" />
                    <SPLIT distance="700" swimtime="00:15:27.64" />
                    <SPLIT distance="750" swimtime="00:16:32.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="83" swimtime="00:04:49.48" resultid="20386" heatid="24342" lane="0" entrytime="00:04:55.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.13" />
                    <SPLIT distance="100" swimtime="00:02:22.97" />
                    <SPLIT distance="150" swimtime="00:03:37.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="43" reactiontime="+92" swimtime="00:05:16.07" resultid="20387" heatid="24368" lane="4" entrytime="00:04:41.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.99" />
                    <SPLIT distance="100" swimtime="00:02:31.93" />
                    <SPLIT distance="150" swimtime="00:03:58.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="80" reactiontime="+78" swimtime="00:02:00.18" resultid="20388" heatid="24403" lane="5" entrytime="00:01:55.84" />
                <RESULT eventid="1578" points="79" reactiontime="+65" swimtime="00:09:27.97" resultid="20389" heatid="24430" lane="3" entrytime="00:09:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.10" />
                    <SPLIT distance="100" swimtime="00:02:28.05" />
                    <SPLIT distance="150" swimtime="00:03:42.13" />
                    <SPLIT distance="200" swimtime="00:04:53.05" />
                    <SPLIT distance="250" swimtime="00:06:07.93" />
                    <SPLIT distance="300" swimtime="00:07:27.11" />
                    <SPLIT distance="350" swimtime="00:08:25.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="43" reactiontime="+79" swimtime="00:02:21.95" resultid="20390" heatid="24437" lane="3" entrytime="00:02:12.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="76" swimtime="00:08:37.70" resultid="20391" heatid="24475" lane="6" entrytime="00:08:20.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.15" />
                    <SPLIT distance="100" swimtime="00:02:04.88" />
                    <SPLIT distance="150" swimtime="00:03:12.53" />
                    <SPLIT distance="200" swimtime="00:04:19.81" />
                    <SPLIT distance="250" swimtime="00:05:25.36" />
                    <SPLIT distance="300" swimtime="00:06:32.27" />
                    <SPLIT distance="350" swimtime="00:07:36.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="107414" nation="POL" region="OL" clubid="20475" name="UKS Manta Warszawa Włochy">
          <CONTACT name="Barański" phone="510835478" />
          <ATHLETES>
            <ATHLETE birthdate="1993-12-20" firstname="Arkadiusz" gender="M" lastname="Aptewicz" nation="POL" license="507414700150" athleteid="20476">
              <RESULTS>
                <RESULT eventid="1613" points="502" reactiontime="+46" swimtime="00:01:02.68" resultid="20477" heatid="24442" lane="1" entrytime="00:01:01.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="599" swimtime="00:04:20.97" resultid="20478" heatid="24482" lane="5" entrytime="00:04:16.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.11" />
                    <SPLIT distance="200" swimtime="00:02:07.40" />
                    <SPLIT distance="300" swimtime="00:03:14.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02201" nation="POL" region="DOL" clubid="20778" name="UKS Shark Rudna">
          <CONTACT name="SZAJNICKI" />
          <ATHLETES>
            <ATHLETE birthdate="1995-02-19" firstname="Katarzyna" gender="F" lastname="Kita" nation="POL" athleteid="20779">
              <RESULTS>
                <RESULT eventid="1062" points="587" reactiontime="+74" swimtime="00:00:28.26" resultid="20780" heatid="24281" lane="4" entrytime="00:00:27.09" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAŁ" nation="POL" region="MAL" clubid="19770" name="UKS Sp 8 Chrzanów">
          <CONTACT city="CHRZANÓW" email="abalp@poczta.onet.pl" name="ZABRZAŃSKI" phone="692076808" state="MAŁ" street="NIEPODLEGŁOŚCI 7 / 46" zip="32 500" />
          <ATHLETES>
            <ATHLETE birthdate="1954-05-12" firstname="Alfred" gender="M" lastname="Zabrzański" nation="POL" athleteid="19771">
              <RESULTS>
                <RESULT eventid="1079" points="268" reactiontime="+88" swimtime="00:00:32.43" resultid="19772" heatid="24287" lane="5" entrytime="00:00:32.50" />
                <RESULT eventid="14189" status="DNS" swimtime="00:00:00.00" resultid="19773" heatid="24315" lane="9" entrytime="00:13:39.00" />
                <RESULT eventid="1205" points="173" swimtime="00:00:43.05" resultid="19774" heatid="24331" lane="6" entrytime="00:00:43.00" />
                <RESULT eventid="1273" points="230" reactiontime="+43" swimtime="00:01:16.53" resultid="19775" heatid="24358" lane="0" entrytime="00:01:13.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="19776" heatid="24418" lane="3" entrytime="00:02:58.60" />
                <RESULT eventid="1681" points="146" reactiontime="+42" swimtime="00:00:49.27" resultid="19777" heatid="24461" lane="5" entrytime="00:00:44.00" />
                <RESULT eventid="1744" points="144" reactiontime="+77" swimtime="00:06:59.82" resultid="19778" heatid="24477" lane="1" entrytime="00:06:38.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.83" />
                    <SPLIT distance="100" swimtime="00:01:31.50" />
                    <SPLIT distance="150" swimtime="00:02:24.87" />
                    <SPLIT distance="200" swimtime="00:03:18.73" />
                    <SPLIT distance="250" swimtime="00:04:14.67" />
                    <SPLIT distance="300" swimtime="00:05:10.07" />
                    <SPLIT distance="350" swimtime="00:06:06.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="LBL" clubid="19760" name="UKS Trójka Puławy">
          <CONTACT name="Gogacz" phone="506694816" />
          <ATHLETES>
            <ATHLETE birthdate="1976-10-28" firstname="Sebastian" gender="M" lastname="Gogacz" nation="POL" license="501203700057" athleteid="19761">
              <RESULTS>
                <RESULT eventid="1113" points="374" reactiontime="+85" swimtime="00:02:38.14" resultid="19762" heatid="24305" lane="7" entrytime="00:02:43.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                    <SPLIT distance="100" swimtime="00:01:17.13" />
                    <SPLIT distance="150" swimtime="00:02:02.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14189" points="350" reactiontime="+89" swimtime="00:10:41.20" resultid="19763" heatid="24317" lane="7" entrytime="00:10:22.31">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.10" />
                    <SPLIT distance="200" swimtime="00:02:33.41" />
                    <SPLIT distance="300" swimtime="00:03:53.35" />
                    <SPLIT distance="400" swimtime="00:05:14.77" />
                    <SPLIT distance="500" swimtime="00:06:35.52" />
                    <SPLIT distance="600" swimtime="00:07:57.15" />
                    <SPLIT distance="750" swimtime="00:10:02.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="324" reactiontime="+53" swimtime="00:02:42.27" resultid="19764" heatid="24371" lane="0" entrytime="00:02:34.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                    <SPLIT distance="100" swimtime="00:01:17.39" />
                    <SPLIT distance="150" swimtime="00:01:59.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="354" reactiontime="+49" swimtime="00:05:44.59" resultid="19765" heatid="24432" lane="5" entrytime="00:05:42.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.38" />
                    <SPLIT distance="100" swimtime="00:01:14.32" />
                    <SPLIT distance="150" swimtime="00:02:01.65" />
                    <SPLIT distance="200" swimtime="00:02:47.63" />
                    <SPLIT distance="250" swimtime="00:03:35.73" />
                    <SPLIT distance="300" swimtime="00:04:25.18" />
                    <SPLIT distance="350" swimtime="00:05:05.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="343" reactiontime="+51" swimtime="00:03:00.84" resultid="23413" heatid="24345" lane="8" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.80" />
                    <SPLIT distance="100" swimtime="00:01:28.19" />
                    <SPLIT distance="150" swimtime="00:02:15.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WODKAT" nation="POL" region="KA" clubid="21968" name="UKS Wodnik 29 Katowice">
          <CONTACT name="Skoczylas" />
          <ATHLETES>
            <ATHLETE birthdate="1937-11-14" firstname="Aleksander" gender="M" lastname="Aleksandrowicz" nation="POL" athleteid="21987">
              <RESULTS>
                <RESULT eventid="1079" points="78" reactiontime="+108" swimtime="00:00:48.76" resultid="21988" heatid="24283" lane="6" entrytime="00:00:51.00" />
                <RESULT eventid="1205" points="63" swimtime="00:01:00.17" resultid="21989" heatid="24329" lane="8" entrytime="00:01:04.00" />
                <RESULT eventid="1474" points="56" reactiontime="+61" swimtime="00:02:14.82" resultid="21990" heatid="24403" lane="6" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="56" reactiontime="+84" swimtime="00:04:51.40" resultid="21991" heatid="24447" lane="1" entrytime="00:04:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.77" />
                    <SPLIT distance="100" swimtime="00:02:22.99" />
                    <SPLIT distance="150" swimtime="00:03:40.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="48" reactiontime="+103" swimtime="00:01:11.10" resultid="21992" heatid="24459" lane="4" entrytime="00:01:11.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-04-21" firstname="Agnieszka" gender="F" lastname="Koenig" nation="POL" athleteid="21993">
              <RESULTS>
                <RESULT eventid="1222" points="91" swimtime="00:05:08.17" resultid="21994" heatid="24338" lane="1" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.28" />
                    <SPLIT distance="100" swimtime="00:02:26.99" />
                    <SPLIT distance="150" swimtime="00:03:46.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="93" swimtime="00:02:21.54" resultid="21995" heatid="24376" lane="2" entrytime="00:02:25.00" />
                <RESULT eventid="1664" points="86" swimtime="00:01:06.39" resultid="21996" heatid="24455" lane="9" entrytime="00:01:08.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-19" firstname="Krzysztof" gender="M" lastname="Kulczyk" nation="POL" athleteid="21969">
              <RESULTS>
                <RESULT eventid="1079" points="233" reactiontime="+92" swimtime="00:00:33.98" resultid="21970" heatid="24286" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1113" points="141" reactiontime="+98" swimtime="00:03:38.75" resultid="21971" heatid="24302" lane="5" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                    <SPLIT distance="100" swimtime="00:01:38.99" />
                    <SPLIT distance="150" swimtime="00:02:49.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="163" swimtime="00:00:43.86" resultid="21972" heatid="24330" lane="4" entrytime="00:00:45.00" />
                <RESULT eventid="1341" points="93" reactiontime="+53" swimtime="00:04:05.48" resultid="21973" heatid="24369" lane="6" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.70" />
                    <SPLIT distance="100" swimtime="00:01:54.85" />
                    <SPLIT distance="150" swimtime="00:03:00.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="253" reactiontime="+84" swimtime="00:00:35.18" resultid="21974" heatid="24392" lane="3" entrytime="00:00:37.00" />
                <RESULT eventid="1474" points="144" reactiontime="+81" swimtime="00:01:38.89" resultid="21975" heatid="24404" lane="6" entrytime="00:01:40.00" />
                <RESULT eventid="1613" points="119" reactiontime="+96" swimtime="00:01:41.17" resultid="21976" heatid="24438" lane="7" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="128" reactiontime="+82" swimtime="00:03:42.06" resultid="21977" heatid="24448" lane="8" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.55" />
                    <SPLIT distance="100" swimtime="00:01:49.95" />
                    <SPLIT distance="150" swimtime="00:02:49.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-28" firstname="Jerzy" gender="M" lastname="Mroziński" nation="POL" athleteid="21997">
              <RESULTS>
                <RESULT eventid="1239" points="289" reactiontime="+44" swimtime="00:03:11.58" resultid="21998" heatid="24344" lane="5" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="297" swimtime="00:01:25.53" resultid="21999" heatid="24383" lane="5" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="382" reactiontime="+45" swimtime="00:00:35.74" resultid="22000" heatid="24464" lane="6" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-04-22" firstname="Tomasz" gender="M" lastname="Skoczylas" nation="POL" athleteid="21978">
              <RESULTS>
                <RESULT eventid="1079" points="348" reactiontime="+104" swimtime="00:00:29.70" resultid="21979" heatid="24290" lane="3" entrytime="00:00:29.50" />
                <RESULT eventid="14189" points="302" reactiontime="+97" swimtime="00:11:13.57" resultid="21980" heatid="24316" lane="5" entrytime="00:10:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.70" />
                    <SPLIT distance="100" swimtime="00:01:13.20" />
                    <SPLIT distance="150" swimtime="00:01:54.30" />
                    <SPLIT distance="200" swimtime="00:02:37.28" />
                    <SPLIT distance="250" swimtime="00:03:19.33" />
                    <SPLIT distance="300" swimtime="00:04:02.42" />
                    <SPLIT distance="350" swimtime="00:04:45.26" />
                    <SPLIT distance="400" swimtime="00:05:28.58" />
                    <SPLIT distance="450" swimtime="00:06:11.94" />
                    <SPLIT distance="500" swimtime="00:06:55.78" />
                    <SPLIT distance="550" swimtime="00:07:39.20" />
                    <SPLIT distance="600" swimtime="00:08:22.55" />
                    <SPLIT distance="650" swimtime="00:09:05.79" />
                    <SPLIT distance="700" swimtime="00:09:49.00" />
                    <SPLIT distance="750" swimtime="00:10:31.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="362" swimtime="00:01:05.82" resultid="21981" heatid="24360" lane="8" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="195" reactiontime="+51" swimtime="00:03:12.26" resultid="21982" heatid="24370" lane="1" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.74" />
                    <SPLIT distance="100" swimtime="00:01:26.86" />
                    <SPLIT distance="150" swimtime="00:02:18.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="230" swimtime="00:01:24.57" resultid="21983" heatid="24406" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="298" reactiontime="+92" swimtime="00:02:32.69" resultid="21984" heatid="24421" lane="7" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                    <SPLIT distance="100" swimtime="00:01:14.32" />
                    <SPLIT distance="150" swimtime="00:01:55.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="235" swimtime="00:01:20.62" resultid="21985" heatid="24439" lane="5" entrytime="00:01:20.00" />
                <RESULT eventid="1647" points="241" reactiontime="+95" swimtime="00:02:59.72" resultid="21986" heatid="24450" lane="0" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.38" />
                    <SPLIT distance="100" swimtime="00:01:27.60" />
                    <SPLIT distance="150" swimtime="00:02:14.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-03-01" firstname="Jan" gender="M" lastname="Wilczek" nation="POL" athleteid="22001">
              <RESULTS>
                <RESULT eventid="1079" points="332" reactiontime="+108" swimtime="00:00:30.17" resultid="22002" heatid="24290" lane="2" entrytime="00:00:29.50" />
                <RESULT eventid="1341" points="170" reactiontime="+101" swimtime="00:03:21.06" resultid="22003" heatid="24370" lane="8" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.59" />
                    <SPLIT distance="100" swimtime="00:01:39.43" />
                    <SPLIT distance="150" swimtime="00:02:33.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="313" reactiontime="+70" swimtime="00:00:32.79" resultid="22004" heatid="24394" lane="1" entrytime="00:00:32.10" />
                <RESULT eventid="1613" points="239" reactiontime="+68" swimtime="00:01:20.21" resultid="22005" heatid="24440" lane="0" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1548" points="311" swimtime="00:02:05.14" resultid="22006" heatid="24426" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.74" />
                    <SPLIT distance="100" swimtime="00:01:01.49" />
                    <SPLIT distance="150" swimtime="00:01:35.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21978" number="1" />
                    <RELAYPOSITION athleteid="21997" number="2" />
                    <RELAYPOSITION athleteid="21969" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="22001" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="01006" nation="POL" region="06" clubid="19836" name="Unia Oświęcim Masters">
          <ATHLETES>
            <ATHLETE birthdate="1952-07-01" firstname="Barbara" gender="F" lastname="Lipniarska-Skubis" nation="POL" license="501006600377" athleteid="19837">
              <RESULTS>
                <RESULT eventid="1187" points="90" swimtime="00:01:00.26" resultid="19838" heatid="24324" lane="2" entrytime="00:00:58.00" />
                <RESULT eventid="1256" points="91" swimtime="00:01:54.77" resultid="19839" heatid="24348" lane="4" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="95" swimtime="00:02:20.18" resultid="19840" heatid="24376" lane="3" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="83" swimtime="00:04:18.71" resultid="19841" heatid="24410" lane="2" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.02" />
                    <SPLIT distance="100" swimtime="00:02:02.91" />
                    <SPLIT distance="150" swimtime="00:03:10.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="101" swimtime="00:01:03.09" resultid="19842" heatid="24455" lane="6" entrytime="00:00:59.00" />
                <RESULT eventid="1721" points="86" swimtime="00:08:55.03" resultid="19843" heatid="24470" lane="6" entrytime="00:08:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.96" />
                    <SPLIT distance="100" swimtime="00:02:04.38" />
                    <SPLIT distance="150" swimtime="00:03:11.71" />
                    <SPLIT distance="200" swimtime="00:04:20.86" />
                    <SPLIT distance="250" swimtime="00:05:30.95" />
                    <SPLIT distance="300" swimtime="00:06:40.38" />
                    <SPLIT distance="350" swimtime="00:07:49.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="21092" name="USKS Ostrołęka">
          <CONTACT name="USKS OSTROŁĘKA" />
          <ATHLETES>
            <ATHLETE birthdate="1990-12-06" firstname="Adam" gender="M" lastname="Janczewski" nation="POL" athleteid="21093">
              <RESULTS>
                <RESULT eventid="1113" points="460" reactiontime="+91" swimtime="00:02:27.64" resultid="21094" heatid="24306" lane="4" entrytime="00:02:26.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.04" />
                    <SPLIT distance="100" swimtime="00:01:10.70" />
                    <SPLIT distance="150" swimtime="00:01:54.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14189" reactiontime="+94" status="OTL" swimtime="00:10:47.13" resultid="21095" heatid="24317" lane="9" entrytime="00:10:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="100" swimtime="00:01:12.80" />
                    <SPLIT distance="150" swimtime="00:01:52.95" />
                    <SPLIT distance="200" swimtime="00:02:34.28" />
                    <SPLIT distance="250" swimtime="00:03:16.39" />
                    <SPLIT distance="300" swimtime="00:03:59.44" />
                    <SPLIT distance="350" swimtime="00:04:41.46" />
                    <SPLIT distance="400" swimtime="00:05:23.17" />
                    <SPLIT distance="450" swimtime="00:06:05.20" />
                    <SPLIT distance="500" swimtime="00:06:46.84" />
                    <SPLIT distance="550" swimtime="00:07:28.17" />
                    <SPLIT distance="600" swimtime="00:08:09.40" />
                    <SPLIT distance="750" swimtime="00:10:09.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="555" reactiontime="+43" swimtime="00:00:57.06" resultid="21096" heatid="24365" lane="1" entrytime="00:00:56.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="031/05" nation="POL" region="LOD" clubid="21103" name="UTW&quot;Masters&quot;ZGIERZ">
          <CONTACT city="ZGIERZ" email="roman.wiczel@gmail.com" name="WICZEL" phone="691-928-922" state="ŁODZK" street="ŁĘCZYCKA 24" zip="95-100" />
          <ATHLETES>
            <ATHLETE birthdate="1973-03-18" firstname="Daria" gender="F" lastname="Fajkowska" nation="POL" license="503105600018" athleteid="21170">
              <RESULTS>
                <RESULT eventid="1062" points="476" reactiontime="+88" swimtime="00:00:30.31" resultid="21171" heatid="24281" lane="0" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT eventid="1187" points="490" swimtime="00:00:34.32" resultid="21172" heatid="24327" lane="5" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT eventid="1457" points="429" reactiontime="+75" swimtime="00:01:16.86" resultid="21173" heatid="24402" lane="7" entrytime="00:01:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="389" reactiontime="+82" swimtime="00:02:49.90" resultid="21174" heatid="24445" lane="1" entrytime="00:02:49.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.51" />
                    <SPLIT distance="100" swimtime="00:01:21.48" />
                    <SPLIT distance="150" swimtime="00:02:06.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-03-08" firstname="Katarzyna" gender="F" lastname="Izert" nation="POL" license="503105600" athleteid="21186">
              <RESULTS>
                <RESULT eventid="1062" points="322" reactiontime="+80" swimtime="00:00:34.50" resultid="21187" heatid="24278" lane="5" entrytime="00:00:34.00" entrycourse="LCM" />
                <RESULT eventid="1256" points="289" reactiontime="+64" swimtime="00:01:18.17" resultid="21188" heatid="24351" lane="2" entrytime="00:01:16.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="252" reactiontime="+77" swimtime="00:02:58.82" resultid="21189" heatid="24412" lane="8" entrytime="00:02:59.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                    <SPLIT distance="100" swimtime="00:01:22.66" />
                    <SPLIT distance="150" swimtime="00:02:10.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" status="DNS" swimtime="00:00:00.00" resultid="21190" heatid="24472" lane="0" entrytime="00:06:00.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-03-01" firstname="Waldemar" gender="M" lastname="Jagiełło" nation="POL" license="503105700036" athleteid="21163">
              <RESULTS>
                <RESULT eventid="1079" points="448" reactiontime="+80" swimtime="00:00:27.31" resultid="21164" heatid="24293" lane="2" entrytime="00:00:27.33" entrycourse="LCM" />
                <RESULT eventid="1113" points="360" reactiontime="+99" swimtime="00:02:40.11" resultid="21165" heatid="24305" lane="2" entrytime="00:02:41.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                    <SPLIT distance="100" swimtime="00:01:16.82" />
                    <SPLIT distance="150" swimtime="00:02:02.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="389" reactiontime="+42" swimtime="00:02:53.48" resultid="21166" heatid="24341" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                    <SPLIT distance="100" swimtime="00:01:17.67" />
                    <SPLIT distance="150" swimtime="00:02:04.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="420" swimtime="00:01:02.63" resultid="21167" heatid="24362" lane="0" entrytime="00:01:01.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="427" reactiontime="+72" swimtime="00:01:15.81" resultid="21168" heatid="24384" lane="4" entrytime="00:01:15.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="360" reactiontime="+70" swimtime="00:00:31.28" resultid="21169" heatid="24395" lane="7" entrytime="00:00:30.66" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-11-08" firstname="Piotr" gender="M" lastname="Kapczyński" nation="POL" license="503105700043" athleteid="21191">
              <RESULTS>
                <RESULT eventid="1079" points="328" reactiontime="+102" swimtime="00:00:30.31" resultid="21192" heatid="24288" lane="3" entrytime="00:00:31.50" entrycourse="LCM" />
                <RESULT eventid="1406" points="274" reactiontime="+63" swimtime="00:01:27.84" resultid="21193" heatid="24383" lane="2" entrytime="00:01:27.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="21194" heatid="24392" lane="4" entrytime="00:00:36.10" entrycourse="LCM" />
                <RESULT eventid="1681" points="310" reactiontime="+61" swimtime="00:00:38.32" resultid="21195" heatid="24463" lane="1" entrytime="00:00:38.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-02-25" firstname="Joanna" gender="F" lastname="Kańska-Papiernik" nation="POL" license="503105600058" athleteid="21175">
              <RESULTS>
                <RESULT eventid="1062" points="409" reactiontime="+76" swimtime="00:00:31.87" resultid="21176" heatid="24279" lane="7" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT eventid="1187" points="381" swimtime="00:00:37.30" resultid="21177" heatid="24326" lane="6" entrytime="00:00:38.00" entrycourse="LCM" />
                <RESULT eventid="1388" points="380" reactiontime="+70" swimtime="00:01:28.49" resultid="21178" heatid="24375" lane="5" />
                <RESULT eventid="1457" points="356" reactiontime="+81" swimtime="00:01:21.80" resultid="21179" heatid="24401" lane="4" entrytime="00:01:22.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="415" swimtime="00:00:39.41" resultid="21180" heatid="24458" lane="9" entrytime="00:00:40.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-12" firstname="Maja" gender="F" lastname="Klusek" nation="POL" license="503105600059" athleteid="21143">
              <RESULTS>
                <RESULT eventid="1096" points="298" reactiontime="+100" swimtime="00:03:08.69" resultid="21144" heatid="24298" lane="5" entrytime="00:03:04.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="209" reactiontime="+78" swimtime="00:03:24.95" resultid="21145" heatid="24367" lane="6" entrytime="00:03:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                    <SPLIT distance="100" swimtime="00:01:30.97" />
                    <SPLIT distance="150" swimtime="00:02:24.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="279" reactiontime="+96" swimtime="00:00:37.36" resultid="21146" heatid="24388" lane="8" entrytime="00:00:36.00" entrycourse="LCM" />
                <RESULT eventid="1595" points="220" reactiontime="+79" swimtime="00:01:31.86" resultid="21147" heatid="24436" lane="8" entrytime="00:01:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-03-17" firstname="Maria" gender="F" lastname="Krakowiak" nation="POL" license="503105600" athleteid="21200">
              <RESULTS>
                <RESULT eventid="1147" points="296" reactiontime="+95" swimtime="00:12:06.90" resultid="21201" heatid="24310" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.72" />
                    <SPLIT distance="100" swimtime="00:01:23.39" />
                    <SPLIT distance="150" swimtime="00:02:08.27" />
                    <SPLIT distance="200" swimtime="00:02:53.53" />
                    <SPLIT distance="250" swimtime="00:03:39.20" />
                    <SPLIT distance="300" swimtime="00:04:24.80" />
                    <SPLIT distance="350" swimtime="00:05:10.90" />
                    <SPLIT distance="400" swimtime="00:05:57.19" />
                    <SPLIT distance="450" swimtime="00:06:43.60" />
                    <SPLIT distance="500" swimtime="00:07:30.41" />
                    <SPLIT distance="550" swimtime="00:08:16.60" />
                    <SPLIT distance="600" swimtime="00:09:03.30" />
                    <SPLIT distance="650" swimtime="00:09:49.75" />
                    <SPLIT distance="700" swimtime="00:10:36.67" />
                    <SPLIT distance="750" swimtime="00:11:23.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="337" reactiontime="+47" swimtime="00:03:19.71" resultid="21202" heatid="24340" lane="7" entrytime="00:03:12.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.05" />
                    <SPLIT distance="100" swimtime="00:01:33.95" />
                    <SPLIT distance="150" swimtime="00:02:26.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="348" swimtime="00:01:31.13" resultid="21203" heatid="24379" lane="9" entrytime="00:01:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="21204" heatid="24412" lane="7" entrytime="00:02:58.00" entrycourse="LCM" />
                <RESULT eventid="1664" points="354" reactiontime="+42" swimtime="00:00:41.56" resultid="21205" heatid="24457" lane="5" entrytime="00:00:41.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-12-03" firstname="Zbigniew" gender="M" lastname="Maciejczyk" nation="POL" license="503105700026" athleteid="21132">
              <RESULTS>
                <RESULT eventid="1079" points="211" reactiontime="+93" swimtime="00:00:35.10" resultid="21133" heatid="24286" lane="6" entrytime="00:00:35.00" entrycourse="LCM" />
                <RESULT eventid="1113" points="126" reactiontime="+85" swimtime="00:03:46.84" resultid="21134" heatid="24302" lane="7" entrytime="00:03:59.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.35" />
                    <SPLIT distance="100" swimtime="00:01:58.44" />
                    <SPLIT distance="150" swimtime="00:03:05.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="195" swimtime="00:01:20.78" resultid="21135" heatid="24357" lane="7" entrytime="00:01:18.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="166" reactiontime="+48" swimtime="00:00:40.49" resultid="21136" heatid="24392" lane="9" entrytime="00:00:39.00" entrycourse="LCM" />
                <RESULT eventid="1613" points="95" reactiontime="+71" swimtime="00:01:49.11" resultid="21137" heatid="24438" lane="2" entrytime="00:01:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-04-11" firstname="Rafał" gender="M" lastname="Maciejewski" nation="POL" license="503105700" athleteid="21181">
              <RESULTS>
                <RESULT eventid="1079" points="230" reactiontime="+96" swimtime="00:00:34.12" resultid="21182" heatid="24287" lane="8" entrytime="00:00:33.50" entrycourse="LCM" />
                <RESULT eventid="1205" points="162" swimtime="00:00:43.97" resultid="21183" heatid="24332" lane="2" entrytime="00:00:40.00" entrycourse="LCM" />
                <RESULT eventid="1273" points="211" reactiontime="+52" swimtime="00:01:18.70" resultid="21184" heatid="24356" lane="5" entrytime="00:01:20.00" entrycourse="LCM" />
                <RESULT eventid="1681" points="223" reactiontime="+43" swimtime="00:00:42.75" resultid="21185" heatid="24461" lane="1" entrytime="00:00:45.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-03" firstname="Urszula" gender="F" lastname="Mróz" nation="POL" license="503105600030" athleteid="21111">
              <RESULTS>
                <RESULT eventid="1062" points="363" reactiontime="+100" swimtime="00:00:33.18" resultid="21112" heatid="24279" lane="0" entrytime="00:00:33.50" entrycourse="LCM" />
                <RESULT eventid="1187" points="286" swimtime="00:00:41.04" resultid="21113" heatid="24326" lane="8" entrytime="00:00:39.20" entrycourse="LCM" />
                <RESULT eventid="1256" points="301" reactiontime="+94" swimtime="00:01:17.10" resultid="21114" heatid="24351" lane="8" entrytime="00:01:17.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="336" reactiontime="+54" swimtime="00:00:35.13" resultid="21115" heatid="24388" lane="1" entrytime="00:00:35.50" entrycourse="LCM" />
                <RESULT eventid="1457" points="223" reactiontime="+88" swimtime="00:01:35.55" resultid="21116" heatid="24401" lane="2" entrytime="00:01:26.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="296" reactiontime="+72" swimtime="00:00:44.08" resultid="21117" heatid="24457" lane="6" entrytime="00:00:42.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-05-12" firstname="Tadeusz" gender="M" lastname="Obiedziński" nation="POL" license="503105700038" athleteid="23409">
              <RESULTS>
                <RESULT eventid="1239" points="153" reactiontime="+80" swimtime="00:03:56.33" resultid="23410" heatid="24343" lane="0" entrytime="00:03:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.65" />
                    <SPLIT distance="100" swimtime="00:01:52.27" />
                    <SPLIT distance="150" swimtime="00:02:55.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="193" reactiontime="+78" swimtime="00:01:38.67" resultid="23411" heatid="24382" lane="1" entrytime="00:01:38.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="238" swimtime="00:00:41.85" resultid="23412" heatid="24462" lane="9" entrytime="00:00:43.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-09" firstname="Włodzimierz" gender="M" lastname="Przytulski" nation="POL" license="503105700027" athleteid="21118">
              <RESULTS>
                <RESULT eventid="1113" status="DNS" swimtime="00:00:00.00" resultid="21119" heatid="24304" lane="2" entrytime="00:03:00.00" entrycourse="LCM" />
                <RESULT eventid="14189" points="230" reactiontime="+91" swimtime="00:12:17.03" resultid="21120" heatid="24316" lane="8" entrytime="00:12:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.92" />
                    <SPLIT distance="100" swimtime="00:01:20.50" />
                    <SPLIT distance="150" swimtime="00:02:04.75" />
                    <SPLIT distance="200" swimtime="00:02:51.61" />
                    <SPLIT distance="250" swimtime="00:03:38.13" />
                    <SPLIT distance="300" swimtime="00:04:25.98" />
                    <SPLIT distance="350" swimtime="00:05:12.97" />
                    <SPLIT distance="400" swimtime="00:06:00.54" />
                    <SPLIT distance="450" swimtime="00:06:48.27" />
                    <SPLIT distance="500" swimtime="00:07:35.86" />
                    <SPLIT distance="550" swimtime="00:08:23.74" />
                    <SPLIT distance="600" swimtime="00:09:11.96" />
                    <SPLIT distance="650" swimtime="00:09:59.80" />
                    <SPLIT distance="700" swimtime="00:10:46.83" />
                    <SPLIT distance="750" swimtime="00:11:34.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="245" swimtime="00:00:38.32" resultid="21121" heatid="24333" lane="9" entrytime="00:00:37.00" entrycourse="LCM" />
                <RESULT eventid="1273" points="289" reactiontime="+58" swimtime="00:01:10.90" resultid="21122" heatid="24359" lane="1" entrytime="00:01:09.00" entrycourse="LCM" />
                <RESULT eventid="1474" status="DNS" swimtime="00:00:00.00" resultid="21123" heatid="24405" lane="5" entrytime="00:01:24.00" entrycourse="LCM" />
                <RESULT eventid="1508" points="250" reactiontime="+64" swimtime="00:02:41.72" resultid="21124" heatid="24420" lane="2" entrytime="00:02:35.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                    <SPLIT distance="100" swimtime="00:01:16.43" />
                    <SPLIT distance="150" swimtime="00:01:59.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="21125" heatid="24449" lane="5" entrytime="00:03:05.00" entrycourse="LCM" />
                <RESULT eventid="1744" points="244" reactiontime="+62" swimtime="00:05:52.12" resultid="21126" heatid="24479" lane="9" entrytime="00:05:42.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:06.53" />
                    <SPLIT distance="100" swimtime="00:01:20.65" />
                    <SPLIT distance="200" swimtime="00:02:50.44" />
                    <SPLIT distance="250" swimtime="00:03:36.78" />
                    <SPLIT distance="300" swimtime="00:04:22.89" />
                    <SPLIT distance="350" swimtime="00:05:09.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1997-05-30" firstname="Adrianna" gender="F" lastname="Rzewuska" nation="POL" license="503105600" athleteid="21196">
              <RESULTS>
                <RESULT eventid="1062" points="367" reactiontime="+79" swimtime="00:00:33.05" resultid="21197" heatid="24281" lane="9" entrytime="00:00:30.15" entrycourse="LCM" />
                <RESULT eventid="1187" points="486" swimtime="00:00:34.41" resultid="21198" heatid="24327" lane="4" entrytime="00:00:32.30" entrycourse="LCM" />
                <RESULT eventid="1457" points="473" reactiontime="+80" swimtime="00:01:14.41" resultid="21199" heatid="24402" lane="4" entrytime="00:01:10.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-02-01" firstname="Andrzej" gender="M" lastname="Sypniewski" nation="POL" license="503105700060" athleteid="21148">
              <RESULTS>
                <RESULT eventid="1079" points="244" reactiontime="+80" swimtime="00:00:33.45" resultid="21149" heatid="24288" lane="8" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="1113" points="219" reactiontime="+78" swimtime="00:03:09.05" resultid="21150" heatid="24303" lane="6" entrytime="00:03:12.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.44" />
                    <SPLIT distance="100" swimtime="00:01:30.55" />
                    <SPLIT distance="150" swimtime="00:02:24.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="228" swimtime="00:00:39.25" resultid="21151" heatid="24332" lane="9" entrytime="00:00:41.00" entrycourse="LCM" />
                <RESULT eventid="1239" points="221" swimtime="00:03:29.26" resultid="21152" heatid="24343" lane="5" entrytime="00:03:27.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" status="DNS" swimtime="00:00:00.00" resultid="21153" heatid="24382" lane="6" entrytime="00:01:33.27" entrycourse="LCM" />
                <RESULT eventid="1474" points="217" swimtime="00:01:26.20" resultid="21154" heatid="24405" lane="8" entrytime="00:01:32.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNF" swimtime="00:00:00.00" resultid="21155" heatid="24439" lane="0" entrytime="00:01:33.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" status="DNS" swimtime="00:00:00.00" resultid="21156" heatid="24462" lane="3" entrytime="00:00:41.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-08-06" firstname="Robert" gender="M" lastname="Szalbierz" nation="POL" license="503105700056" athleteid="21138">
              <RESULTS>
                <RESULT eventid="1079" points="271" reactiontime="+92" swimtime="00:00:32.31" resultid="21139" heatid="24290" lane="8" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="21140" heatid="24358" lane="3" entrytime="00:01:10.00" entrycourse="LCM" />
                <RESULT eventid="1440" points="268" reactiontime="+46" swimtime="00:00:34.51" resultid="21141" heatid="24394" lane="9" entrytime="00:00:33.50" entrycourse="LCM" />
                <RESULT eventid="1508" status="DNS" swimtime="00:00:00.00" resultid="21142" heatid="24419" lane="9" entrytime="00:02:57.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-22" firstname="Roman" gender="M" lastname="Wiczel" nation="POL" license="503105700034" athleteid="21104">
              <RESULTS>
                <RESULT eventid="1205" points="160" swimtime="00:00:44.16" resultid="21105" heatid="24331" lane="1" entrytime="00:00:44.00" entrycourse="LCM" />
                <RESULT eventid="1239" points="187" reactiontime="+81" swimtime="00:03:41.18" resultid="21106" heatid="24343" lane="2" entrytime="00:03:33.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.47" />
                    <SPLIT distance="100" swimtime="00:01:49.57" />
                    <SPLIT distance="150" swimtime="00:02:47.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="192" reactiontime="+69" swimtime="00:01:38.82" resultid="21107" heatid="24382" lane="2" entrytime="00:01:35.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="147" swimtime="00:01:38.07" resultid="21108" heatid="24404" lane="4" entrytime="00:01:37.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="140" swimtime="00:03:35.40" resultid="21109" heatid="24448" lane="5" entrytime="00:03:30.00" entrycourse="LCM" />
                <RESULT eventid="1681" points="226" reactiontime="+53" swimtime="00:00:42.56" resultid="21110" heatid="24462" lane="1" entrytime="00:00:42.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-08-25" firstname="Michał" gender="M" lastname="Woźniak" nation="POL" license="503105700039" athleteid="21157">
              <RESULTS>
                <RESULT eventid="1205" points="471" swimtime="00:00:30.84" resultid="21158" heatid="24335" lane="6" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT eventid="1440" points="487" swimtime="00:00:28.29" resultid="21159" heatid="24390" lane="9" />
                <RESULT eventid="1474" points="443" reactiontime="+67" swimtime="00:01:08.01" resultid="21160" heatid="24408" lane="0" entrytime="00:01:07.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" points="426" reactiontime="+72" swimtime="00:01:06.16" resultid="21161" heatid="24437" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="380" reactiontime="+57" swimtime="00:02:34.51" resultid="21162" heatid="24452" lane="9" entrytime="00:02:28.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                    <SPLIT distance="150" swimtime="00:01:55.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-12" firstname="Małgorzata" gender="F" lastname="Ścibiorek" nation="POL" license="503105600028" athleteid="21127">
              <RESULTS>
                <RESULT eventid="1096" points="453" reactiontime="+86" swimtime="00:02:44.11" resultid="21128" heatid="24299" lane="1" entrytime="00:02:49.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                    <SPLIT distance="100" swimtime="00:01:16.40" />
                    <SPLIT distance="150" swimtime="00:02:04.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1324" points="330" reactiontime="+61" swimtime="00:02:56.20" resultid="21129" heatid="24367" lane="5" entrytime="00:02:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="441" swimtime="00:00:32.09" resultid="21130" heatid="24389" lane="7" entrytime="00:00:33.50" entrycourse="LCM" />
                <RESULT eventid="1595" points="414" reactiontime="+41" swimtime="00:01:14.40" resultid="21131" heatid="24436" lane="3" entrytime="00:01:10.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" status="DNS" swimtime="00:00:00.00" resultid="21206" heatid="24374" lane="8" entrytime="00:02:11.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21157" number="1" />
                    <RELAYPOSITION athleteid="21148" number="2" />
                    <RELAYPOSITION athleteid="21118" number="3" />
                    <RELAYPOSITION athleteid="21163" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" status="DNS" swimtime="00:00:00.00" resultid="21207" heatid="24427" lane="9" entrytime="00:02:03.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21163" number="1" />
                    <RELAYPOSITION athleteid="21148" number="2" />
                    <RELAYPOSITION athleteid="21118" number="3" />
                    <RELAYPOSITION athleteid="21157" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="212" swimtime="00:02:36.48" resultid="21208" heatid="24373" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21104" number="1" />
                    <RELAYPOSITION athleteid="21191" number="2" />
                    <RELAYPOSITION athleteid="21138" number="3" reactiontime="+23" />
                    <RELAYPOSITION athleteid="21132" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1548" points="227" reactiontime="+61" swimtime="00:02:19.01" resultid="21209" heatid="24426" lane="5" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21191" number="1" reactiontime="+61" />
                    <RELAYPOSITION athleteid="21104" number="2" />
                    <RELAYPOSITION athleteid="21132" number="3" reactiontime="+9" />
                    <RELAYPOSITION athleteid="21138" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1358" points="444" reactiontime="+123" swimtime="00:02:19.32" resultid="21210" heatid="24372" lane="4" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                    <SPLIT distance="100" swimtime="00:01:13.13" />
                    <SPLIT distance="150" swimtime="00:01:46.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21170" number="1" reactiontime="+123" />
                    <RELAYPOSITION athleteid="21175" number="2" />
                    <RELAYPOSITION athleteid="21127" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="21111" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1525" points="411" swimtime="00:02:09.67" resultid="21211" heatid="24425" lane="5" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21127" number="1" />
                    <RELAYPOSITION athleteid="21143" number="2" />
                    <RELAYPOSITION athleteid="21111" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="21170" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" reactiontime="+99" swimtime="00:02:05.62" resultid="21212" heatid="24309" lane="3" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.07" />
                    <SPLIT distance="100" swimtime="00:01:02.24" />
                    <SPLIT distance="150" swimtime="00:01:36.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21170" number="1" reactiontime="+99" />
                    <RELAYPOSITION athleteid="21127" number="2" />
                    <RELAYPOSITION athleteid="21181" number="3" reactiontime="+72" />
                    <RELAYPOSITION athleteid="21163" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" reactiontime="+75" swimtime="00:02:18.90" resultid="21213" heatid="24468" lane="2" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:47.58" />
                    <SPLIT distance="100" swimtime="00:01:12.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21170" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="21191" number="2" />
                    <RELAYPOSITION athleteid="21138" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="21175" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" reactiontime="+93" swimtime="00:02:06.56" resultid="21214" heatid="24308" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                    <SPLIT distance="100" swimtime="00:01:04.88" />
                    <SPLIT distance="150" swimtime="00:01:35.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21111" number="1" reactiontime="+93" />
                    <RELAYPOSITION athleteid="21175" number="2" />
                    <RELAYPOSITION athleteid="21191" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="21138" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1698" reactiontime="+82" swimtime="00:02:27.14" resultid="21215" heatid="24468" lane="1" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.39" />
                    <SPLIT distance="100" swimtime="00:01:22.34" />
                    <SPLIT distance="150" swimtime="00:01:57.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21111" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="21148" number="2" />
                    <RELAYPOSITION athleteid="21118" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="21127" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="04214" nation="POL" region="14" clubid="22096" name="Warsaw Masters Team">
          <CONTACT city="Warszawa" email="jarecka.skorykow@gmail.com" name="jarecka" phone="606286265" street="Żółkiewskiego 40/11" zip="04-305" />
          <ATHLETES>
            <ATHLETE birthdate="1977-08-13" firstname="Dymitr" gender="M" lastname="Bielski" nation="POL" athleteid="22387">
              <RESULTS>
                <RESULT eventid="1079" points="248" reactiontime="+97" swimtime="00:00:33.26" resultid="22388" heatid="24284" lane="6" entrytime="00:00:40.00" />
                <RESULT eventid="1113" points="222" reactiontime="+95" swimtime="00:03:08.03" resultid="22389" heatid="24303" lane="4" entrytime="00:03:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                    <SPLIT distance="100" swimtime="00:01:34.07" />
                    <SPLIT distance="150" swimtime="00:02:23.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="290" reactiontime="+57" swimtime="00:03:11.26" resultid="22390" heatid="24344" lane="6" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.98" />
                    <SPLIT distance="100" swimtime="00:01:29.61" />
                    <SPLIT distance="150" swimtime="00:02:19.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="213" reactiontime="+67" swimtime="00:02:50.66" resultid="22391" heatid="24419" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                    <SPLIT distance="100" swimtime="00:01:19.77" />
                    <SPLIT distance="150" swimtime="00:02:05.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-03-04" firstname="Stefan" gender="M" lastname="Borodziuk" nation="POL" athleteid="22422">
              <RESULTS>
                <RESULT eventid="1079" points="128" reactiontime="+82" swimtime="00:00:41.43" resultid="22423" heatid="24285" lane="9" entrytime="00:00:39.00" />
                <RESULT eventid="14189" points="71" reactiontime="+92" swimtime="00:18:08.15" resultid="22424" heatid="24314" lane="8" entrytime="00:16:55.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:54.26" />
                    <SPLIT distance="200" swimtime="00:04:09.90" />
                    <SPLIT distance="300" swimtime="00:06:30.10" />
                    <SPLIT distance="400" swimtime="00:08:52.46" />
                    <SPLIT distance="500" swimtime="00:11:16.49" />
                    <SPLIT distance="550" swimtime="00:12:26.01" />
                    <SPLIT distance="600" swimtime="00:13:36.80" />
                    <SPLIT distance="650" swimtime="00:14:47.37" />
                    <SPLIT distance="700" swimtime="00:15:58.21" />
                    <SPLIT distance="750" swimtime="00:17:04.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="102" swimtime="00:00:51.31" resultid="22425" heatid="24329" lane="4" entrytime="00:00:52.50" />
                <RESULT eventid="1273" points="117" reactiontime="+59" swimtime="00:01:35.65" resultid="22426" heatid="24356" lane="1" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="90" reactiontime="+71" swimtime="00:01:55.30" resultid="22427" heatid="24404" lane="9" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="92" reactiontime="+86" swimtime="00:03:45.89" resultid="22428" heatid="24416" lane="4" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.47" />
                    <SPLIT distance="100" swimtime="00:01:45.57" />
                    <SPLIT distance="150" swimtime="00:02:47.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="80" reactiontime="+80" swimtime="00:04:19.20" resultid="22429" heatid="24447" lane="2" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.90" />
                    <SPLIT distance="100" swimtime="00:02:04.00" />
                    <SPLIT distance="150" swimtime="00:03:14.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="82" reactiontime="+47" swimtime="00:08:25.64" resultid="22430" heatid="24475" lane="5" entrytime="00:07:50.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:48.87" />
                    <SPLIT distance="200" swimtime="00:04:00.68" />
                    <SPLIT distance="300" swimtime="00:06:16.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-20" firstname="Katarzyna" gender="F" lastname="Dziedzic" nation="POL" athleteid="22498">
              <RESULTS>
                <RESULT eventid="1096" points="355" reactiontime="+88" swimtime="00:02:57.97" resultid="22499" heatid="24299" lane="0" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.56" />
                    <SPLIT distance="100" swimtime="00:01:25.14" />
                    <SPLIT distance="150" swimtime="00:02:16.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="301" reactiontime="+89" swimtime="00:22:52.14" resultid="22500" heatid="24319" lane="3" entrytime="00:22:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.87" />
                    <SPLIT distance="100" swimtime="00:01:20.97" />
                    <SPLIT distance="150" swimtime="00:02:04.73" />
                    <SPLIT distance="200" swimtime="00:02:49.21" />
                    <SPLIT distance="250" swimtime="00:03:33.73" />
                    <SPLIT distance="300" swimtime="00:04:18.96" />
                    <SPLIT distance="350" swimtime="00:05:04.46" />
                    <SPLIT distance="400" swimtime="00:05:50.98" />
                    <SPLIT distance="450" swimtime="00:06:37.50" />
                    <SPLIT distance="500" swimtime="00:07:23.62" />
                    <SPLIT distance="550" swimtime="00:08:10.18" />
                    <SPLIT distance="600" swimtime="00:08:55.93" />
                    <SPLIT distance="650" swimtime="00:09:42.26" />
                    <SPLIT distance="700" swimtime="00:10:28.82" />
                    <SPLIT distance="750" swimtime="00:11:15.08" />
                    <SPLIT distance="800" swimtime="00:12:01.52" />
                    <SPLIT distance="850" swimtime="00:12:48.08" />
                    <SPLIT distance="900" swimtime="00:13:35.21" />
                    <SPLIT distance="950" swimtime="00:14:21.90" />
                    <SPLIT distance="1000" swimtime="00:15:08.66" />
                    <SPLIT distance="1050" swimtime="00:15:55.28" />
                    <SPLIT distance="1100" swimtime="00:16:41.61" />
                    <SPLIT distance="1150" swimtime="00:17:28.17" />
                    <SPLIT distance="1200" swimtime="00:18:14.66" />
                    <SPLIT distance="1250" swimtime="00:19:01.33" />
                    <SPLIT distance="1300" swimtime="00:19:48.29" />
                    <SPLIT distance="1350" swimtime="00:20:35.08" />
                    <SPLIT distance="1400" swimtime="00:21:22.11" />
                    <SPLIT distance="1450" swimtime="00:22:08.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="250" reactiontime="+79" swimtime="00:00:38.75" resultid="22501" heatid="24388" lane="4" entrytime="00:00:34.20" />
                <RESULT eventid="1555" points="317" reactiontime="+81" swimtime="00:06:30.35" resultid="22502" heatid="24429" lane="3" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.81" />
                    <SPLIT distance="100" swimtime="00:01:33.82" />
                    <SPLIT distance="150" swimtime="00:02:23.27" />
                    <SPLIT distance="200" swimtime="00:03:12.94" />
                    <SPLIT distance="250" swimtime="00:04:04.26" />
                    <SPLIT distance="300" swimtime="00:04:59.27" />
                    <SPLIT distance="350" swimtime="00:05:46.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="314" swimtime="00:03:02.43" resultid="22503" heatid="24444" lane="4" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.38" />
                    <SPLIT distance="100" swimtime="00:01:28.75" />
                    <SPLIT distance="150" swimtime="00:02:16.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-11-26" firstname="Ewa" gender="F" lastname="Galica" nation="POL" athleteid="22455">
              <RESULTS>
                <RESULT eventid="1062" points="376" reactiontime="+76" swimtime="00:00:32.78" resultid="22456" heatid="24280" lane="8" entrytime="00:00:31.50" />
                <RESULT eventid="1256" points="341" swimtime="00:01:13.97" resultid="22457" heatid="24352" lane="1" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="292" swimtime="00:00:36.80" resultid="22458" heatid="24389" lane="9" entrytime="00:00:34.00" />
                <RESULT eventid="1491" points="341" reactiontime="+49" swimtime="00:02:41.71" resultid="22459" heatid="24413" lane="9" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                    <SPLIT distance="100" swimtime="00:01:16.54" />
                    <SPLIT distance="150" swimtime="00:01:59.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="352" reactiontime="+61" swimtime="00:05:34.84" resultid="24645" heatid="24469" lane="2" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                    <SPLIT distance="100" swimtime="00:01:16.99" />
                    <SPLIT distance="150" swimtime="00:01:59.48" />
                    <SPLIT distance="200" swimtime="00:02:43.61" />
                    <SPLIT distance="250" swimtime="00:03:27.19" />
                    <SPLIT distance="300" swimtime="00:04:11.06" />
                    <SPLIT distance="350" swimtime="00:04:54.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-06-13" firstname="Marcin" gender="M" lastname="Giejsztowt" nation="POL" athleteid="22477">
              <RESULTS>
                <RESULT eventid="1273" points="418" swimtime="00:01:02.73" resultid="22478" heatid="24361" lane="6" entrytime="00:01:03.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="417" swimtime="00:02:16.51" resultid="22479" heatid="24422" lane="3" entrytime="00:02:17.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                    <SPLIT distance="100" swimtime="00:01:05.23" />
                    <SPLIT distance="150" swimtime="00:01:41.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="424" swimtime="00:04:52.71" resultid="22480" heatid="24481" lane="1" entrytime="00:04:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                    <SPLIT distance="100" swimtime="00:01:08.13" />
                    <SPLIT distance="150" swimtime="00:01:45.71" />
                    <SPLIT distance="200" swimtime="00:02:23.72" />
                    <SPLIT distance="250" swimtime="00:03:01.93" />
                    <SPLIT distance="300" swimtime="00:03:40.47" />
                    <SPLIT distance="350" swimtime="00:04:18.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-30" firstname="Monika" gender="F" lastname="Jarecka-Skorykow" nation="POL" athleteid="22375">
              <RESULTS>
                <RESULT eventid="1664" points="340" reactiontime="+75" swimtime="00:00:42.12" resultid="22376" heatid="24456" lane="6" entrytime="00:00:46.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-05-28" firstname="Konrad" gender="M" lastname="Karnaszewski" nation="POL" athleteid="22440">
              <RESULTS>
                <RESULT eventid="1079" points="647" reactiontime="+69" swimtime="00:00:24.17" resultid="22441" heatid="24296" lane="1" entrytime="00:00:24.99" />
                <RESULT eventid="1273" points="625" swimtime="00:00:54.86" resultid="22442" heatid="24365" lane="2" entrytime="00:00:55.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="558" reactiontime="+55" swimtime="00:00:27.05" resultid="22443" heatid="24397" lane="3" entrytime="00:00:27.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-09-27" firstname="Wojciech" gender="M" lastname="Kossowski" nation="POL" athleteid="22444">
              <RESULTS>
                <RESULT eventid="1113" points="146" reactiontime="+138" swimtime="00:03:36.23" resultid="22445" heatid="24303" lane="8" entrytime="00:03:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.70" />
                    <SPLIT distance="100" swimtime="00:01:51.44" />
                    <SPLIT distance="150" swimtime="00:02:48.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="204" reactiontime="+131" swimtime="00:03:35.01" resultid="22446" heatid="24343" lane="7" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.54" />
                    <SPLIT distance="100" swimtime="00:01:44.40" />
                    <SPLIT distance="150" swimtime="00:02:40.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="203" reactiontime="+127" swimtime="00:01:37.07" resultid="22447" heatid="24382" lane="3" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="139" reactiontime="+125" swimtime="00:07:50.16" resultid="22448" heatid="24431" lane="7" entrytime="00:07:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.15" />
                    <SPLIT distance="100" swimtime="00:01:59.63" />
                    <SPLIT distance="150" swimtime="00:03:05.83" />
                    <SPLIT distance="200" swimtime="00:04:11.50" />
                    <SPLIT distance="250" swimtime="00:05:11.71" />
                    <SPLIT distance="300" swimtime="00:06:11.51" />
                    <SPLIT distance="350" swimtime="00:07:03.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="227" reactiontime="+114" swimtime="00:00:42.49" resultid="22449" heatid="24462" lane="8" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-06-17" firstname="Leszek" gender="M" lastname="Madej" nation="POL" athleteid="22465">
              <RESULTS>
                <RESULT eventid="1079" points="410" reactiontime="+77" swimtime="00:00:28.14" resultid="22466" heatid="24293" lane="9" entrytime="00:00:27.93" />
                <RESULT eventid="1273" points="419" swimtime="00:01:02.67" resultid="22467" heatid="24361" lane="5" entrytime="00:01:03.31" />
                <RESULT eventid="1508" points="387" swimtime="00:02:19.92" resultid="22468" heatid="24422" lane="8" entrytime="00:02:19.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                    <SPLIT distance="100" swimtime="00:01:09.40" />
                    <SPLIT distance="150" swimtime="00:01:44.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="342" reactiontime="+79" swimtime="00:00:37.08" resultid="22469" heatid="24463" lane="4" entrytime="00:00:37.18" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-05-04" firstname="Ewa" gender="F" lastname="Matlak" nation="POL" athleteid="22493">
              <RESULTS>
                <RESULT eventid="1147" points="336" reactiontime="+76" swimtime="00:11:36.81" resultid="22494" heatid="24311" lane="6" entrytime="00:12:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.31" />
                    <SPLIT distance="100" swimtime="00:01:19.52" />
                    <SPLIT distance="150" swimtime="00:02:03.16" />
                    <SPLIT distance="200" swimtime="00:02:47.11" />
                    <SPLIT distance="250" swimtime="00:03:30.97" />
                    <SPLIT distance="300" swimtime="00:04:14.88" />
                    <SPLIT distance="350" swimtime="00:04:59.04" />
                    <SPLIT distance="400" swimtime="00:05:43.42" />
                    <SPLIT distance="450" swimtime="00:06:27.93" />
                    <SPLIT distance="500" swimtime="00:07:12.04" />
                    <SPLIT distance="550" swimtime="00:07:56.52" />
                    <SPLIT distance="600" swimtime="00:08:41.44" />
                    <SPLIT distance="650" swimtime="00:09:25.61" />
                    <SPLIT distance="700" swimtime="00:10:10.28" />
                    <SPLIT distance="750" swimtime="00:10:54.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="373" swimtime="00:00:33.91" resultid="22495" heatid="24388" lane="2" entrytime="00:00:35.33" />
                <RESULT eventid="1491" points="361" swimtime="00:02:38.62" resultid="22496" heatid="24413" lane="1" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                    <SPLIT distance="100" swimtime="00:01:14.82" />
                    <SPLIT distance="150" swimtime="00:01:57.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="355" swimtime="00:05:33.91" resultid="22497" heatid="24472" lane="5" entrytime="00:05:42.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.27" />
                    <SPLIT distance="200" swimtime="00:02:42.78" />
                    <SPLIT distance="300" swimtime="00:04:09.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-10-11" firstname="Grzegorz" gender="M" lastname="Matyszewski" nation="POL" athleteid="22399">
              <RESULTS>
                <RESULT eventid="1079" points="242" reactiontime="+73" swimtime="00:00:33.53" resultid="22400" heatid="24287" lane="7" entrytime="00:00:33.00" />
                <RESULT eventid="1113" points="184" reactiontime="+81" swimtime="00:03:20.31" resultid="22401" heatid="24303" lane="1" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.59" />
                    <SPLIT distance="100" swimtime="00:01:39.78" />
                    <SPLIT distance="150" swimtime="00:02:30.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="260" swimtime="00:03:18.45" resultid="22402" heatid="24344" lane="0" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.25" />
                    <SPLIT distance="100" swimtime="00:01:34.50" />
                    <SPLIT distance="150" swimtime="00:02:25.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="186" swimtime="00:01:22.04" resultid="22403" heatid="24357" lane="9" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="272" reactiontime="+77" swimtime="00:01:28.08" resultid="22404" heatid="24383" lane="7" entrytime="00:01:27.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="149" swimtime="00:03:12.02" resultid="22405" heatid="24418" lane="0" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.68" />
                    <SPLIT distance="100" swimtime="00:01:32.63" />
                    <SPLIT distance="150" swimtime="00:02:22.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="291" swimtime="00:00:39.13" resultid="22406" heatid="24463" lane="0" entrytime="00:00:38.60" />
                <RESULT eventid="1744" points="150" swimtime="00:06:53.42" resultid="22407" heatid="24476" lane="4" entrytime="00:06:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.99" />
                    <SPLIT distance="100" swimtime="00:01:33.66" />
                    <SPLIT distance="150" swimtime="00:02:25.69" />
                    <SPLIT distance="200" swimtime="00:03:17.27" />
                    <SPLIT distance="250" swimtime="00:04:12.01" />
                    <SPLIT distance="300" swimtime="00:05:06.24" />
                    <SPLIT distance="350" swimtime="00:06:01.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-12-17" firstname="Michał" gender="M" lastname="Nowak" nation="POL" athleteid="22431">
              <RESULTS>
                <RESULT eventid="1113" points="191" reactiontime="+85" swimtime="00:03:17.82" resultid="22432" heatid="24303" lane="7" entrytime="00:03:15.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.28" />
                    <SPLIT distance="100" swimtime="00:01:39.30" />
                    <SPLIT distance="150" swimtime="00:02:31.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="239" swimtime="00:03:24.03" resultid="22433" heatid="24344" lane="9" entrytime="00:03:20.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.27" />
                    <SPLIT distance="100" swimtime="00:01:37.37" />
                    <SPLIT distance="150" swimtime="00:02:29.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="265" swimtime="00:01:28.80" resultid="22434" heatid="24383" lane="9" entrytime="00:01:29.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="160" reactiontime="+72" swimtime="00:07:28.30" resultid="22435" heatid="24431" lane="6" entrytime="00:07:18.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.41" />
                    <SPLIT distance="100" swimtime="00:01:39.54" />
                    <SPLIT distance="200" swimtime="00:03:54.85" />
                    <SPLIT distance="250" swimtime="00:04:52.07" />
                    <SPLIT distance="300" swimtime="00:05:51.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="297" reactiontime="+80" swimtime="00:00:38.86" resultid="22436" heatid="24463" lane="7" entrytime="00:00:38.37" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-08-01" firstname="Joanna" gender="F" lastname="Olszewska" nation="POL" athleteid="22481">
              <RESULTS>
                <RESULT eventid="1222" points="306" swimtime="00:03:26.39" resultid="22482" heatid="24339" lane="5" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="323" swimtime="00:01:33.45" resultid="22483" heatid="24378" lane="5" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="231" reactiontime="+82" swimtime="00:03:03.91" resultid="22484" heatid="24411" lane="4" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.83" />
                    <SPLIT distance="100" swimtime="00:01:30.44" />
                    <SPLIT distance="150" swimtime="00:02:18.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="330" swimtime="00:00:42.51" resultid="22485" heatid="24457" lane="0" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-05-14" firstname="Bartosz" gender="M" lastname="Ostrowski" nation="POL" athleteid="22470">
              <RESULTS>
                <RESULT eventid="1079" points="403" reactiontime="+96" swimtime="00:00:28.29" resultid="22471" heatid="24290" lane="5" entrytime="00:00:29.50" />
                <RESULT eventid="1113" points="226" reactiontime="+85" swimtime="00:03:07.00" resultid="22472" heatid="24304" lane="4" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                    <SPLIT distance="100" swimtime="00:01:30.01" />
                    <SPLIT distance="150" swimtime="00:02:22.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="338" reactiontime="+63" swimtime="00:03:01.84" resultid="22473" heatid="24345" lane="4" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                    <SPLIT distance="100" swimtime="00:01:21.90" />
                    <SPLIT distance="150" swimtime="00:02:12.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="400" swimtime="00:01:17.47" resultid="22474" heatid="24384" lane="6" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="293" swimtime="00:02:33.52" resultid="22475" heatid="24420" lane="0" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.23" />
                    <SPLIT distance="100" swimtime="00:01:14.12" />
                    <SPLIT distance="150" swimtime="00:01:54.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="403" reactiontime="+71" swimtime="00:00:35.13" resultid="22476" heatid="24465" lane="3" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-02-17" firstname="Zbigniew" gender="M" lastname="Paluszak" nation="POL" athleteid="22381">
              <RESULTS>
                <RESULT eventid="1239" points="158" reactiontime="+65" swimtime="00:03:54.10" resultid="22382" heatid="24342" lane="3" entrytime="00:03:54.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.07" />
                    <SPLIT distance="100" swimtime="00:01:50.42" />
                    <SPLIT distance="150" swimtime="00:02:52.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="145" reactiontime="+46" swimtime="00:01:48.66" resultid="22383" heatid="24381" lane="6" entrytime="00:01:49.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="109" swimtime="00:03:33.46" resultid="22384" heatid="24417" lane="9" entrytime="00:03:41.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.65" />
                    <SPLIT distance="100" swimtime="00:01:41.58" />
                    <SPLIT distance="150" swimtime="00:02:38.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="155" reactiontime="+64" swimtime="00:00:48.25" resultid="22385" heatid="24460" lane="4" entrytime="00:00:49.13" />
                <RESULT eventid="1744" points="115" reactiontime="+78" swimtime="00:07:31.41" resultid="22386" heatid="24475" lane="4" entrytime="00:07:35.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.99" />
                    <SPLIT distance="100" swimtime="00:01:44.94" />
                    <SPLIT distance="150" swimtime="00:02:42.80" />
                    <SPLIT distance="200" swimtime="00:03:40.81" />
                    <SPLIT distance="250" swimtime="00:04:38.63" />
                    <SPLIT distance="300" swimtime="00:05:37.36" />
                    <SPLIT distance="350" swimtime="00:06:36.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-24" firstname="Jan" gender="M" lastname="Pfitzner" nation="POL" athleteid="22460">
              <RESULTS>
                <RESULT eventid="1079" points="448" reactiontime="+76" swimtime="00:00:27.32" resultid="22461" heatid="24294" lane="5" entrytime="00:00:26.50" />
                <RESULT eventid="1273" points="489" swimtime="00:00:59.53" resultid="22462" heatid="24364" lane="6" entrytime="00:00:57.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1508" points="490" swimtime="00:02:09.33" resultid="22463" heatid="24424" lane="8" entrytime="00:02:07.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.89" />
                    <SPLIT distance="100" swimtime="00:01:03.30" />
                    <SPLIT distance="150" swimtime="00:01:36.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="410" swimtime="00:04:56.12" resultid="22464" heatid="24482" lane="1" entrytime="00:04:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                    <SPLIT distance="100" swimtime="00:01:08.60" />
                    <SPLIT distance="150" swimtime="00:01:46.18" />
                    <SPLIT distance="200" swimtime="00:02:24.53" />
                    <SPLIT distance="250" swimtime="00:03:03.07" />
                    <SPLIT distance="300" swimtime="00:03:40.91" />
                    <SPLIT distance="350" swimtime="00:04:19.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-06-10" firstname="Łukasz" gender="M" lastname="Rybiński" nation="POL" athleteid="22377">
              <RESULTS>
                <RESULT eventid="1079" points="307" reactiontime="+93" swimtime="00:00:30.98" resultid="22378" heatid="24289" lane="9" entrytime="00:00:31.00" />
                <RESULT eventid="1273" points="287" reactiontime="+44" swimtime="00:01:11.10" resultid="22379" heatid="24358" lane="5" entrytime="00:01:10.00" />
                <RESULT eventid="1406" points="258" reactiontime="+41" swimtime="00:01:29.58" resultid="22380" heatid="24382" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-12-11" firstname="Igor" gender="M" lastname="Rębas" nation="POL" athleteid="22408">
              <RESULTS>
                <RESULT eventid="1273" points="616" swimtime="00:00:55.13" resultid="22409" heatid="24354" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="539" swimtime="00:00:27.36" resultid="22410" heatid="24390" lane="0" />
                <RESULT eventid="1508" points="472" swimtime="00:02:10.99" resultid="22411" heatid="24416" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.42" />
                    <SPLIT distance="100" swimtime="00:01:01.82" />
                    <SPLIT distance="150" swimtime="00:01:37.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1613" status="DNS" swimtime="00:00:00.00" resultid="22412" heatid="24437" lane="1" />
                <RESULT eventid="1744" points="195" reactiontime="+74" swimtime="00:06:18.93" resultid="22413" heatid="24474" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.98" />
                    <SPLIT distance="100" swimtime="00:01:16.62" />
                    <SPLIT distance="150" swimtime="00:02:05.84" />
                    <SPLIT distance="200" swimtime="00:02:56.05" />
                    <SPLIT distance="250" swimtime="00:03:45.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-10-03" firstname="Ryszard" gender="M" lastname="Sielski" nation="POL" athleteid="22414">
              <RESULTS>
                <RESULT eventid="1079" points="8" swimtime="00:01:44.49" resultid="22415" heatid="24283" lane="1" entrytime="00:01:10.00" />
                <RESULT eventid="1205" points="25" swimtime="00:01:21.98" resultid="22416" heatid="24328" lane="4" entrytime="00:01:25.00" />
                <RESULT eventid="1239" points="29" swimtime="00:06:51.35" resultid="22417" heatid="24342" lane="8" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:33.72" />
                    <SPLIT distance="100" swimtime="00:03:18.63" />
                    <SPLIT distance="150" swimtime="00:05:03.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="31" swimtime="00:03:01.63" resultid="22418" heatid="24380" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:32.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1474" points="21" reactiontime="+83" swimtime="00:03:07.16" resultid="22419" heatid="24403" lane="7" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:28.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="20" reactiontime="+123" swimtime="00:06:50.91" resultid="22420" heatid="24446" lane="4" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:36.00" />
                    <SPLIT distance="100" swimtime="00:03:21.73" />
                    <SPLIT distance="150" swimtime="00:05:05.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="36" swimtime="00:01:18.52" resultid="22421" heatid="24459" lane="5" entrytime="00:01:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-04-17" firstname="Andrzej" gender="M" lastname="Skorykow" nation="POL" athleteid="22373">
              <RESULTS>
                <RESULT eventid="1744" points="379" swimtime="00:05:04.03" resultid="22374" heatid="24481" lane="0" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.08" />
                    <SPLIT distance="100" swimtime="00:01:12.81" />
                    <SPLIT distance="150" swimtime="00:01:50.60" />
                    <SPLIT distance="200" swimtime="00:02:29.99" />
                    <SPLIT distance="250" swimtime="00:03:07.71" />
                    <SPLIT distance="300" swimtime="00:03:47.65" />
                    <SPLIT distance="350" swimtime="00:04:26.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-03" firstname="Robert" gender="M" lastname="Sutowski" nation="POL" athleteid="22392">
              <RESULTS>
                <RESULT eventid="1079" points="145" reactiontime="+95" swimtime="00:00:39.75" resultid="22393" heatid="24285" lane="8" entrytime="00:00:38.71" />
                <RESULT eventid="14189" points="166" reactiontime="+105" swimtime="00:13:41.06" resultid="22394" heatid="24314" lane="4" entrytime="00:13:40.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.43" />
                    <SPLIT distance="100" swimtime="00:01:36.07" />
                    <SPLIT distance="150" swimtime="00:02:28.82" />
                    <SPLIT distance="200" swimtime="00:03:20.79" />
                    <SPLIT distance="250" swimtime="00:04:13.08" />
                    <SPLIT distance="300" swimtime="00:05:04.74" />
                    <SPLIT distance="350" swimtime="00:05:56.17" />
                    <SPLIT distance="400" swimtime="00:06:47.85" />
                    <SPLIT distance="450" swimtime="00:09:25.21" />
                    <SPLIT distance="500" swimtime="00:08:33.27" />
                    <SPLIT distance="550" swimtime="00:11:09.43" />
                    <SPLIT distance="600" swimtime="00:10:16.62" />
                    <SPLIT distance="700" swimtime="00:12:00.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="165" reactiontime="+45" swimtime="00:01:25.49" resultid="22395" heatid="24356" lane="7" entrytime="00:01:26.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="92" reactiontime="+87" swimtime="00:00:49.21" resultid="22396" heatid="24390" lane="4" entrytime="00:00:49.63" />
                <RESULT eventid="1508" points="153" reactiontime="+87" swimtime="00:03:10.66" resultid="22397" heatid="24417" lane="4" entrytime="00:03:10.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.93" />
                    <SPLIT distance="100" swimtime="00:01:33.54" />
                    <SPLIT distance="150" swimtime="00:02:23.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" points="169" reactiontime="+43" swimtime="00:06:37.89" resultid="22398" heatid="24477" lane="7" entrytime="00:06:37.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:05:51.22" />
                    <SPLIT distance="100" swimtime="00:01:32.59" />
                    <SPLIT distance="200" swimtime="00:03:15.86" />
                    <SPLIT distance="300" swimtime="00:04:59.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-07-26" firstname="Anna" gender="F" lastname="Szemberg" nation="POL" athleteid="22437">
              <RESULTS>
                <RESULT eventid="1165" points="86" swimtime="00:34:39.12" resultid="22438" heatid="24318" lane="5" entrytime="00:34:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.53" />
                    <SPLIT distance="150" swimtime="00:03:21.79" />
                    <SPLIT distance="250" swimtime="00:05:40.88" />
                    <SPLIT distance="300" swimtime="00:06:50.18" />
                    <SPLIT distance="350" swimtime="00:07:58.81" />
                    <SPLIT distance="400" swimtime="00:09:08.23" />
                    <SPLIT distance="450" swimtime="00:10:17.62" />
                    <SPLIT distance="500" swimtime="00:16:03.76" />
                    <SPLIT distance="550" swimtime="00:12:36.82" />
                    <SPLIT distance="600" swimtime="00:18:23.70" />
                    <SPLIT distance="650" swimtime="00:14:55.21" />
                    <SPLIT distance="700" swimtime="00:20:43.76" />
                    <SPLIT distance="750" swimtime="00:17:13.82" />
                    <SPLIT distance="850" swimtime="00:19:34.60" />
                    <SPLIT distance="950" swimtime="00:21:53.50" />
                    <SPLIT distance="1050" swimtime="00:24:13.32" />
                    <SPLIT distance="1150" swimtime="00:26:33.40" />
                    <SPLIT distance="1200" swimtime="00:27:42.37" />
                    <SPLIT distance="1250" swimtime="00:28:53.16" />
                    <SPLIT distance="1300" swimtime="00:30:02.42" />
                    <SPLIT distance="1350" swimtime="00:31:13.46" />
                    <SPLIT distance="1400" swimtime="00:32:22.97" />
                    <SPLIT distance="1450" swimtime="00:33:32.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="88" swimtime="00:08:50.59" resultid="22439" heatid="24470" lane="7" entrytime="00:08:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:03:17.02" />
                    <SPLIT distance="100" swimtime="00:02:08.18" />
                    <SPLIT distance="200" swimtime="00:04:24.37" />
                    <SPLIT distance="250" swimtime="00:05:33.01" />
                    <SPLIT distance="350" swimtime="00:07:47.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-08-12" firstname="Jakub" gender="M" lastname="Szulc" nation="POL" athleteid="22486">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="22487" heatid="24290" lane="4" entrytime="00:00:29.50" />
                <RESULT eventid="14189" status="DNS" swimtime="00:00:00.00" resultid="22488" heatid="24316" lane="4" entrytime="00:10:55.00" />
                <RESULT eventid="1273" points="362" swimtime="00:01:05.81" resultid="22489" heatid="24360" lane="5" entrytime="00:01:05.00" />
                <RESULT eventid="1440" points="372" reactiontime="+58" swimtime="00:00:30.94" resultid="22490" heatid="24394" lane="7" entrytime="00:00:32.00" />
                <RESULT eventid="1508" points="358" swimtime="00:02:23.56" resultid="22491" heatid="24421" lane="5" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                    <SPLIT distance="100" swimtime="00:01:11.33" />
                    <SPLIT distance="150" swimtime="00:01:48.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1744" status="DNS" swimtime="00:00:00.00" resultid="22492" heatid="24480" lane="8" entrytime="00:05:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-10-04" firstname="Maciej" gender="M" lastname="Szymański" nation="POL" athleteid="22504">
              <RESULTS>
                <RESULT eventid="1079" points="541" reactiontime="+68" swimtime="00:00:25.65" resultid="22505" heatid="24296" lane="7" entrytime="00:00:24.98" />
                <RESULT eventid="1205" points="541" reactiontime="+78" swimtime="00:00:29.45" resultid="22506" heatid="24336" lane="1" entrytime="00:00:28.80" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="22507" heatid="24355" lane="9" />
                <RESULT eventid="1440" points="535" reactiontime="+63" swimtime="00:00:27.42" resultid="22508" heatid="24390" lane="7" />
                <RESULT eventid="1474" points="526" reactiontime="+75" swimtime="00:01:04.22" resultid="22509" heatid="24408" lane="6" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-08-30" firstname="Mirosław" gender="M" lastname="Warchoł" nation="POL" athleteid="22450">
              <RESULTS>
                <RESULT eventid="1079" points="363" reactiontime="+85" swimtime="00:00:29.29" resultid="22451" heatid="24290" lane="7" entrytime="00:00:29.88" />
                <RESULT eventid="1273" points="369" swimtime="00:01:05.36" resultid="22452" heatid="24359" lane="5" entrytime="00:01:07.69" />
                <RESULT eventid="1474" points="297" swimtime="00:01:17.63" resultid="22453" heatid="24406" lane="5" entrytime="00:01:17.88" />
                <RESULT eventid="1647" points="298" reactiontime="+83" swimtime="00:02:47.49" resultid="22454" heatid="24450" lane="2" entrytime="00:02:48.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.00" />
                    <SPLIT distance="100" swimtime="00:01:21.79" />
                    <SPLIT distance="150" swimtime="00:02:05.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1381" points="549" reactiontime="+110" swimtime="00:01:54.05" resultid="22510" heatid="24374" lane="4" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.75" />
                    <SPLIT distance="100" swimtime="00:01:03.77" />
                    <SPLIT distance="150" swimtime="00:01:30.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22504" number="1" reactiontime="+110" />
                    <RELAYPOSITION athleteid="22470" number="2" />
                    <RELAYPOSITION athleteid="22408" number="3" reactiontime="+17" />
                    <RELAYPOSITION athleteid="22440" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="3">
              <RESULTS>
                <RESULT comment="S1 - Pływak utracił kontakt stopami z platformą startową słupka zanim poprzedzający go pływak dotknął ściany (przedwczesna zmiana sztafetowa). (Time: 12:16), Na 3 zmianie" eventid="1381" reactiontime="+80" status="DSQ" swimtime="00:02:07.71" resultid="22512" heatid="24374" lane="7" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.78" />
                    <SPLIT distance="100" swimtime="00:01:08.93" />
                    <SPLIT distance="150" swimtime="00:01:39.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22460" number="1" reactiontime="+80" status="DSQ" />
                    <RELAYPOSITION athleteid="22387" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="22477" number="3" reactiontime="-23" status="DSQ" />
                    <RELAYPOSITION athleteid="22486" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1548" points="599" swimtime="00:01:40.63" resultid="22513" heatid="24427" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.00" />
                    <SPLIT distance="100" swimtime="00:00:51.16" />
                    <SPLIT distance="150" swimtime="00:01:16.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22440" number="1" />
                    <RELAYPOSITION athleteid="22460" number="2" />
                    <RELAYPOSITION athleteid="22504" number="3" reactiontime="+10" />
                    <RELAYPOSITION athleteid="22408" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1130" reactiontime="+74" swimtime="00:02:03.05" resultid="22511" heatid="24309" lane="6" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.54" />
                    <SPLIT distance="100" swimtime="00:01:00.81" />
                    <SPLIT distance="150" swimtime="00:01:32.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22504" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="22498" number="2" />
                    <RELAYPOSITION athleteid="22455" number="3" reactiontime="-68" />
                    <RELAYPOSITION athleteid="22450" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="5">
              <RESULTS>
                <RESULT eventid="1698" swimtime="00:02:20.44" resultid="22514" heatid="24468" lane="6" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.97" />
                    <SPLIT distance="100" swimtime="00:01:11.36" />
                    <SPLIT distance="150" swimtime="00:01:47.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="22373" number="1" />
                    <RELAYPOSITION athleteid="22470" number="2" />
                    <RELAYPOSITION athleteid="22498" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="22455" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="SLA" clubid="19851" name="Weteran  Zabrze">
          <CONTACT city="ZABRZE" email="weteranzabrze@op.pl" name="BOSOWSKI  WŁODZIMIERZ" street="ŚW.JANA  4A/4" zip="41-803" />
          <ATHLETES>
            <ATHLETE birthdate="1959-01-11" firstname="Jan" gender="M" lastname="Barucha" nation="POL" license="102611600021" athleteid="19857">
              <RESULTS>
                <RESULT eventid="1079" points="279" reactiontime="+75" swimtime="00:00:31.98" resultid="19858" heatid="24288" lane="7" entrytime="00:00:31.80" />
                <RESULT eventid="1205" points="195" swimtime="00:00:41.37" resultid="19859" heatid="24332" lane="0" entrytime="00:00:40.24" />
                <RESULT eventid="1273" points="249" swimtime="00:01:14.47" resultid="19860" heatid="24358" lane="7" entrytime="00:01:11.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="213" swimtime="00:00:37.29" resultid="19861" heatid="24393" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1474" points="194" swimtime="00:01:29.51" resultid="19862" heatid="24405" lane="3" entrytime="00:01:24.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" status="DNS" swimtime="00:00:00.00" resultid="19863" heatid="24449" lane="7" entrytime="00:03:12.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-12-02" firstname="Renata" gender="F" lastname="Bastek" nation="POL" license="102611600023" athleteid="19881">
              <RESULTS>
                <RESULT eventid="1062" points="223" reactiontime="+80" swimtime="00:00:38.99" resultid="19882" heatid="24277" lane="3" entrytime="00:00:39.00" />
                <RESULT eventid="1096" points="134" reactiontime="+76" swimtime="00:04:06.05" resultid="19883" heatid="24297" lane="3" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.05" />
                    <SPLIT distance="100" swimtime="00:01:59.87" />
                    <SPLIT distance="150" swimtime="00:03:14.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="184" swimtime="00:00:47.52" resultid="19884" heatid="24325" lane="0" entrytime="00:00:48.00" />
                <RESULT eventid="1256" points="183" reactiontime="+66" swimtime="00:01:31.05" resultid="19885" heatid="24349" lane="4" entrytime="00:01:30.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="161" reactiontime="+66" swimtime="00:03:27.62" resultid="19886" heatid="24411" lane="8" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.68" />
                    <SPLIT distance="100" swimtime="00:01:40.80" />
                    <SPLIT distance="150" swimtime="00:02:35.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-05-23" firstname="Janina" gender="F" lastname="Bosowska" nation="POL" license="102611600024" athleteid="19918">
              <RESULTS>
                <RESULT eventid="1388" points="101" reactiontime="+85" swimtime="00:02:17.26" resultid="19919" heatid="24376" lane="4" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="119" reactiontime="+78" swimtime="00:00:59.61" resultid="19920" heatid="24455" lane="1" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-05-22" firstname="Włodzimierz" gender="M" lastname="Bosowski" nation="POL" license="102611600014" athleteid="19915">
              <RESULTS>
                <RESULT eventid="1079" points="99" reactiontime="+117" swimtime="00:00:45.13" resultid="19916" heatid="24284" lane="4" entrytime="00:00:39.50" />
                <RESULT eventid="1440" status="DNS" swimtime="00:00:00.00" resultid="19917" heatid="24391" lane="0" entrytime="00:00:48.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-02-18" firstname="Genowefa" gender="F" lastname="Drużyńska" nation="POL" athleteid="19852">
              <RESULTS>
                <RESULT eventid="1187" points="78" swimtime="00:01:03.19" resultid="19853" heatid="24323" lane="5" entrytime="00:01:15.00" />
                <RESULT eventid="1222" points="81" reactiontime="+94" swimtime="00:05:21.05" resultid="19854" heatid="24338" lane="8" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.62" />
                    <SPLIT distance="100" swimtime="00:02:34.97" />
                    <SPLIT distance="150" swimtime="00:03:58.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="89" reactiontime="+93" swimtime="00:02:23.41" resultid="19855" heatid="24376" lane="6" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="97" reactiontime="+78" swimtime="00:01:03.85" resultid="19856" heatid="24455" lane="0" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-11-29" firstname="Daniel" gender="M" lastname="Fecica" nation="POL" license="102611600018" athleteid="19887">
              <RESULTS>
                <RESULT eventid="1239" points="169" reactiontime="+74" swimtime="00:03:48.88" resultid="19888" heatid="24343" lane="8" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.76" />
                    <SPLIT distance="100" swimtime="00:01:50.75" />
                    <SPLIT distance="150" swimtime="00:02:51.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="159" reactiontime="+50" swimtime="00:01:45.27" resultid="19889" heatid="24382" lane="9" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="167" reactiontime="+92" swimtime="00:00:47.10" resultid="19890" heatid="24461" lane="6" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-03-12" firstname="Krystyna" gender="F" lastname="Fecica" nation="POL" license="102611600019" athleteid="19891">
              <RESULTS>
                <RESULT eventid="1147" points="108" reactiontime="+99" swimtime="00:16:57.94" resultid="19892" heatid="24310" lane="3" entrytime="00:16:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.76" />
                    <SPLIT distance="100" swimtime="00:01:56.73" />
                    <SPLIT distance="150" swimtime="00:02:59.71" />
                    <SPLIT distance="200" swimtime="00:04:05.14" />
                    <SPLIT distance="250" swimtime="00:05:10.72" />
                    <SPLIT distance="300" swimtime="00:06:15.46" />
                    <SPLIT distance="350" swimtime="00:07:19.46" />
                    <SPLIT distance="400" swimtime="00:08:23.92" />
                    <SPLIT distance="450" swimtime="00:09:27.66" />
                    <SPLIT distance="500" swimtime="00:10:32.58" />
                    <SPLIT distance="550" swimtime="00:11:35.46" />
                    <SPLIT distance="600" swimtime="00:12:41.37" />
                    <SPLIT distance="650" swimtime="00:13:45.06" />
                    <SPLIT distance="700" swimtime="00:14:50.36" />
                    <SPLIT distance="750" swimtime="00:15:55.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="138" reactiontime="+85" swimtime="00:04:28.90" resultid="19893" heatid="24338" lane="5" entrytime="00:04:12.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:07.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="155" reactiontime="+87" swimtime="00:01:59.20" resultid="19894" heatid="24377" lane="7" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="94" reactiontime="+77" swimtime="00:00:53.57" resultid="19895" heatid="24386" lane="5" entrytime="00:00:53.00" />
                <RESULT eventid="1595" points="104" reactiontime="+105" swimtime="00:01:57.97" resultid="19896" heatid="24435" lane="7" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="163" reactiontime="+105" swimtime="00:00:53.75" resultid="19897" heatid="24455" lane="3" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-02-18" firstname="Grażyna" gender="F" lastname="Kiszczak" nation="POL" license="102611100006" athleteid="19867">
              <RESULTS>
                <RESULT eventid="1062" points="199" swimtime="00:00:40.50" resultid="19868" heatid="24277" lane="7" entrytime="00:00:39.50" />
                <RESULT eventid="1187" points="228" swimtime="00:00:44.29" resultid="19869" heatid="24325" lane="8" entrytime="00:00:47.50" />
                <RESULT eventid="1423" points="113" reactiontime="+62" swimtime="00:00:50.39" resultid="19870" heatid="24387" lane="9" entrytime="00:00:46.00" />
                <RESULT eventid="1457" points="207" reactiontime="+73" swimtime="00:01:37.92" resultid="19871" heatid="24400" lane="6" entrytime="00:01:44.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1630" points="192" reactiontime="+81" swimtime="00:03:34.90" resultid="19872" heatid="24444" lane="3" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.77" />
                    <SPLIT distance="100" swimtime="00:01:46.20" />
                    <SPLIT distance="150" swimtime="00:02:42.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-28" firstname="Wiesław" gender="M" lastname="Kornicki" nation="POL" license="102611600015" athleteid="19873">
              <RESULTS>
                <RESULT eventid="1079" points="253" reactiontime="+92" swimtime="00:00:33.02" resultid="19874" heatid="24287" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1273" points="190" reactiontime="+82" swimtime="00:01:21.46" resultid="19875" heatid="24356" lane="4" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1440" points="192" swimtime="00:00:38.56" resultid="19876" heatid="24392" lane="2" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-04-14" firstname="Gabriela" gender="F" lastname="Molenda" nation="POL" athleteid="19908">
              <RESULTS>
                <RESULT eventid="1187" points="123" swimtime="00:00:54.29" resultid="19909" heatid="24324" lane="5" entrytime="00:00:52.94" />
                <RESULT eventid="1256" points="155" reactiontime="+86" swimtime="00:01:36.14" resultid="19910" heatid="24349" lane="5" entrytime="00:01:36.57" />
                <RESULT eventid="1457" points="119" reactiontime="+89" swimtime="00:01:57.85" resultid="19911" heatid="24399" lane="5" />
                <RESULT eventid="1491" points="157" reactiontime="+77" swimtime="00:03:29.17" resultid="19912" heatid="24411" lane="7" entrytime="00:03:29.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.11" />
                    <SPLIT distance="100" swimtime="00:01:40.45" />
                    <SPLIT distance="150" swimtime="00:02:35.12" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G4 - Pływak wykonał więcej niż jedno pociągnięcie ramieniem (lub obydwoma ramionami równocześnie) w pozycji na piersiach w trakcie wykonywania nawrotu. (Time: 9:37), G-6" eventid="1630" reactiontime="+69" status="DSQ" swimtime="00:04:06.80" resultid="19913" heatid="24443" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.97" />
                    <SPLIT distance="100" swimtime="00:02:01.91" />
                    <SPLIT distance="150" swimtime="00:03:05.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1721" points="153" reactiontime="+60" swimtime="00:07:22.01" resultid="19914" heatid="24471" lane="9" entrytime="00:07:20.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.64" />
                    <SPLIT distance="100" swimtime="00:01:42.16" />
                    <SPLIT distance="150" swimtime="00:02:37.91" />
                    <SPLIT distance="200" swimtime="00:03:34.51" />
                    <SPLIT distance="250" swimtime="00:04:31.67" />
                    <SPLIT distance="300" swimtime="00:05:28.74" />
                    <SPLIT distance="350" swimtime="00:06:25.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-02-25" firstname="Bernard" gender="M" lastname="Poloczek" nation="POL" license="102611100004" athleteid="19877">
              <RESULTS>
                <RESULT eventid="1205" points="160" swimtime="00:00:44.19" resultid="19878" heatid="24331" lane="0" entrytime="00:00:44.11" />
                <RESULT eventid="1474" points="135" reactiontime="+70" swimtime="00:01:40.83" resultid="19879" heatid="24404" lane="2" entrytime="00:01:41.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="116" reactiontime="+67" swimtime="00:03:48.84" resultid="19880" heatid="24448" lane="7" entrytime="00:03:41.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.81" />
                    <SPLIT distance="100" swimtime="00:01:48.78" />
                    <SPLIT distance="150" swimtime="00:02:48.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-07-27" firstname="Danuta" gender="F" lastname="Skorupa" nation="POL" license="102611600020" athleteid="19864">
              <RESULTS>
                <RESULT eventid="1187" points="50" swimtime="00:01:12.97" resultid="19865" heatid="24324" lane="8" entrytime="00:01:02.00" />
                <RESULT eventid="1664" status="DNS" swimtime="00:00:00.00" resultid="19866" heatid="24454" lane="5" entrytime="00:01:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-03-13" firstname="Joanna" gender="F" lastname="Sulewska -Bielak" nation="POL" athleteid="19905">
              <RESULTS>
                <RESULT eventid="1062" status="DNS" swimtime="00:00:00.00" resultid="19906" heatid="24279" lane="9" entrytime="00:00:33.50" />
                <RESULT eventid="1423" status="DNS" swimtime="00:00:00.00" resultid="19907" heatid="24388" lane="9" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-11-02" firstname="Beata" gender="F" lastname="Sulewska" nation="POL" license="102611600016" athleteid="19898">
              <RESULTS>
                <RESULT eventid="1147" points="436" reactiontime="+86" swimtime="00:10:39.30" resultid="19899" heatid="24312" lane="2" entrytime="00:10:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                    <SPLIT distance="100" swimtime="00:01:15.09" />
                    <SPLIT distance="150" swimtime="00:01:54.44" />
                    <SPLIT distance="200" swimtime="00:02:34.25" />
                    <SPLIT distance="250" swimtime="00:03:14.70" />
                    <SPLIT distance="300" swimtime="00:03:54.99" />
                    <SPLIT distance="350" swimtime="00:04:35.50" />
                    <SPLIT distance="400" swimtime="00:05:16.44" />
                    <SPLIT distance="450" swimtime="00:05:57.25" />
                    <SPLIT distance="500" swimtime="00:06:37.95" />
                    <SPLIT distance="550" swimtime="00:07:18.78" />
                    <SPLIT distance="600" swimtime="00:07:59.52" />
                    <SPLIT distance="650" swimtime="00:08:39.92" />
                    <SPLIT distance="700" swimtime="00:09:20.47" />
                    <SPLIT distance="750" swimtime="00:10:00.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="410" reactiontime="+90" swimtime="00:03:07.13" resultid="19900" heatid="24340" lane="6" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.33" />
                    <SPLIT distance="100" swimtime="00:01:29.52" />
                    <SPLIT distance="150" swimtime="00:02:17.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1388" points="400" reactiontime="+57" swimtime="00:01:27.03" resultid="19901" heatid="24379" lane="8" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="435" reactiontime="+49" swimtime="00:02:29.06" resultid="19902" heatid="24414" lane="0" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.33" />
                    <SPLIT distance="100" swimtime="00:01:13.20" />
                    <SPLIT distance="150" swimtime="00:01:51.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1664" points="410" reactiontime="+46" swimtime="00:00:39.55" resultid="19903" heatid="24458" lane="0" entrytime="00:00:39.80" />
                <RESULT eventid="1721" points="424" reactiontime="+65" swimtime="00:05:14.74" resultid="19904" heatid="24473" lane="1" entrytime="00:05:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                    <SPLIT distance="100" swimtime="00:01:15.91" />
                    <SPLIT distance="150" swimtime="00:01:55.82" />
                    <SPLIT distance="200" swimtime="00:02:35.54" />
                    <SPLIT distance="250" swimtime="00:03:15.77" />
                    <SPLIT distance="300" swimtime="00:03:56.04" />
                    <SPLIT distance="350" swimtime="00:04:36.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1381" points="134" reactiontime="+67" swimtime="00:03:02.37" resultid="19923" heatid="24373" lane="6" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.81" />
                    <SPLIT distance="100" swimtime="00:01:29.40" />
                    <SPLIT distance="150" swimtime="00:02:16.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="19857" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="19887" number="2" />
                    <RELAYPOSITION athleteid="19873" number="3" reactiontime="+116" />
                    <RELAYPOSITION athleteid="19915" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="1548" points="158" reactiontime="+76" swimtime="00:02:36.86" resultid="19925" heatid="24426" lane="3" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.31" />
                    <SPLIT distance="100" swimtime="00:01:26.61" />
                    <SPLIT distance="150" swimtime="00:02:02.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="19915" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="19887" number="2" />
                    <RELAYPOSITION athleteid="19873" number="3" reactiontime="+36" />
                    <RELAYPOSITION athleteid="19857" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1358" points="154" reactiontime="+76" swimtime="00:03:18.13" resultid="19922" heatid="24372" lane="7" entrytime="00:03:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.07" />
                    <SPLIT distance="150" swimtime="00:02:38.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="19867" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="19918" number="2" />
                    <RELAYPOSITION athleteid="19891" number="3" />
                    <RELAYPOSITION athleteid="19881" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="F" number="4">
              <RESULTS>
                <RESULT eventid="1525" points="156" reactiontime="+61" swimtime="00:02:59.11" resultid="19924" heatid="24425" lane="7" entrytime="00:03:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.19" />
                    <SPLIT distance="100" swimtime="00:01:34.71" />
                    <SPLIT distance="150" swimtime="00:02:17.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="19908" number="1" reactiontime="+61" />
                    <RELAYPOSITION athleteid="19891" number="2" />
                    <RELAYPOSITION athleteid="19867" number="3" />
                    <RELAYPOSITION athleteid="19881" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1130" swimtime="00:02:44.48" resultid="19921" heatid="24308" lane="2" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.46" />
                    <SPLIT distance="100" swimtime="00:01:31.32" />
                    <SPLIT distance="150" swimtime="00:02:11.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="19867" number="1" />
                    <RELAYPOSITION athleteid="19891" number="2" />
                    <RELAYPOSITION athleteid="19887" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="19857" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="280" gender="X" number="6">
              <RESULTS>
                <RESULT eventid="1698" reactiontime="+133" swimtime="00:02:51.28" resultid="19926" heatid="24467" lane="4" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.14" />
                    <SPLIT distance="100" swimtime="00:01:32.94" />
                    <SPLIT distance="150" swimtime="00:02:11.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="19867" number="1" reactiontime="+133" />
                    <RELAYPOSITION athleteid="19887" number="2" />
                    <RELAYPOSITION athleteid="19873" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="19881" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SLAWRO" nation="POL" region="WR" clubid="20238" name="WKS Śląsk Wrocław">
          <CONTACT email="marrot68@wp.pl" name="Rother Marek" phone="785209045" />
          <ATHLETES>
            <ATHLETE birthdate="1968-03-21" firstname="Marek" gender="M" lastname="Rother" nation="POL" athleteid="20239">
              <RESULTS>
                <RESULT eventid="1205" points="439" reactiontime="+81" swimtime="00:00:31.57" resultid="20240" heatid="24335" lane="1" entrytime="00:00:30.60" />
                <RESULT eventid="1474" points="426" reactiontime="+71" swimtime="00:01:08.87" resultid="20241" heatid="24408" lane="9" entrytime="00:01:07.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1647" points="429" reactiontime="+71" swimtime="00:02:28.36" resultid="20242" heatid="24452" lane="8" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.35" />
                    <SPLIT distance="100" swimtime="00:01:12.49" />
                    <SPLIT distance="150" swimtime="00:01:51.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="LBS" clubid="20899" name="ZKS Drzonków">
          <CONTACT city="Zielona Góra" email="llfpiotr@gmail.com" fax="-" name="Barta" phone="602347348" state="LUB" street="Odrzańska" zip="66-016" />
          <ATHLETES>
            <ATHLETE birthdate="1971-03-18" firstname="Piotr" gender="M" lastname="Barta" nation="POL" license="-" athleteid="20900">
              <RESULTS>
                <RESULT eventid="1239" points="480" reactiontime="+85" swimtime="00:02:41.77" resultid="20901" heatid="24346" lane="2" entrytime="00:02:39.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.91" />
                    <SPLIT distance="100" swimtime="00:01:17.84" />
                    <SPLIT distance="150" swimtime="00:01:59.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1406" points="442" swimtime="00:01:14.91" resultid="20902" heatid="24385" lane="0" entrytime="00:01:13.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1578" points="413" reactiontime="+75" swimtime="00:05:27.36" resultid="20903" heatid="24433" lane="8" entrytime="00:05:27.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                    <SPLIT distance="100" swimtime="00:01:11.53" />
                    <SPLIT distance="150" swimtime="00:01:57.79" />
                    <SPLIT distance="200" swimtime="00:02:43.17" />
                    <SPLIT distance="250" swimtime="00:03:26.65" />
                    <SPLIT distance="300" swimtime="00:04:12.07" />
                    <SPLIT distance="350" swimtime="00:04:49.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1681" points="437" swimtime="00:00:34.19" resultid="20904" heatid="24465" lane="5" entrytime="00:00:33.50" entrycourse="LCM" />
                <RESULT eventid="1744" points="449" reactiontime="+69" swimtime="00:04:47.22" resultid="20905" heatid="24481" lane="4" entrytime="00:04:47.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.50" />
                    <SPLIT distance="100" swimtime="00:01:09.14" />
                    <SPLIT distance="150" swimtime="00:01:45.06" />
                    <SPLIT distance="200" swimtime="00:02:20.85" />
                    <SPLIT distance="250" swimtime="00:02:56.70" />
                    <SPLIT distance="300" swimtime="00:03:33.36" />
                    <SPLIT distance="350" swimtime="00:04:10.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>

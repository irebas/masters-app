<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Dolnoslaski Okregowy Zwiazek Plywacki" version="11.69132">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Wrocław" name="OTWARTE LETNIE MISTRZOSTWA DOLNEGO ŚLĄSKA – VI Memoriał im. Andrzeja Wernera" course="LCM" deadline="2019-05-20" hostclub.url="http://www.dozp.eu" organizer="Dolnośląski Okręgowy Związek Pływacki " result.url="http://ivetyming.pl" startmethod="1" timing="AUTOMATIC" nation="POL">
      <AGEDATE value="2021-01-01" type="YEAR" />
      <POOL name="im. Marka Petrusewicza" lanemax="9" />
      <FACILITY city="Wrocław" name="im. Marka Petrusewicza" nation="POL" street="Wejherowska 34" zip="50-239" />
      <POINTTABLE pointtableid="3014" name="FINA Point Scoring" version="2021" />
      <CONTACT city="Wrocław" email="nadobny@nadobny.net" />
      <QUALIFY from="2016-01-01" until="2021-05-25" conversion="ESP.CONVERSION" />
      <SESSIONS>
        <SESSION date="2021-05-28" daytime="09:00" endtime="12:17" number="1" warmupfrom="07:50" warmupuntil="08:50">
          <EVENTS>
            <EVENT eventid="44378" daytime="09:00" gender="M" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46215" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46898" />
                    <RANKING order="2" place="2" resultid="47020" />
                    <RANKING order="3" place="3" resultid="47830" />
                    <RANKING order="4" place="4" resultid="47661" />
                    <RANKING order="5" place="5" resultid="48256" />
                    <RANKING order="6" place="6" resultid="46484" />
                    <RANKING order="7" place="7" resultid="47594" />
                    <RANKING order="8" place="8" resultid="47985" />
                    <RANKING order="9" place="9" resultid="46919" />
                    <RANKING order="10" place="10" resultid="46729" />
                    <RANKING order="11" place="11" resultid="48263" />
                    <RANKING order="12" place="12" resultid="50384" />
                    <RANKING order="13" place="13" resultid="49095" />
                    <RANKING order="14" place="14" resultid="47991" />
                    <RANKING order="15" place="15" resultid="47137" />
                    <RANKING order="16" place="16" resultid="48511" />
                    <RANKING order="17" place="17" resultid="47140" />
                    <RANKING order="18" place="-1" resultid="48732" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="44379" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47163" />
                    <RANKING order="2" place="2" resultid="50314" />
                    <RANKING order="3" place="3" resultid="50363" />
                    <RANKING order="4" place="4" resultid="48727" />
                    <RANKING order="5" place="5" resultid="46912" />
                    <RANKING order="6" place="6" resultid="46646" />
                    <RANKING order="7" place="7" resultid="48056" />
                    <RANKING order="8" place="8" resultid="46477" />
                    <RANKING order="9" place="9" resultid="48742" />
                    <RANKING order="10" place="10" resultid="48502" />
                    <RANKING order="11" place="11" resultid="50321" />
                    <RANKING order="12" place="12" resultid="48631" />
                    <RANKING order="13" place="13" resultid="47959" />
                    <RANKING order="14" place="14" resultid="46905" />
                    <RANKING order="15" place="15" resultid="47034" />
                    <RANKING order="16" place="16" resultid="48491" />
                    <RANKING order="17" place="17" resultid="50370" />
                    <RANKING order="18" place="18" resultid="46626" />
                    <RANKING order="19" place="19" resultid="47972" />
                    <RANKING order="20" place="19" resultid="50377" />
                    <RANKING order="21" place="21" resultid="48235" />
                    <RANKING order="22" place="22" resultid="49074" />
                    <RANKING order="23" place="23" resultid="47924" />
                    <RANKING order="24" place="24" resultid="48240" />
                    <RANKING order="25" place="25" resultid="48413" />
                    <RANKING order="26" place="26" resultid="48250" />
                    <RANKING order="27" place="27" resultid="46717" />
                    <RANKING order="28" place="28" resultid="46857" />
                    <RANKING order="29" place="29" resultid="50336" />
                    <RANKING order="30" place="30" resultid="47603" />
                    <RANKING order="31" place="31" resultid="50330" />
                    <RANKING order="32" place="32" resultid="50390" />
                    <RANKING order="33" place="33" resultid="49088" />
                    <RANKING order="34" place="34" resultid="50326" />
                    <RANKING order="35" place="35" resultid="48737" />
                    <RANKING order="36" place="36" resultid="48062" />
                    <RANKING order="37" place="37" resultid="48245" />
                    <RANKING order="38" place="38" resultid="47100" />
                    <RANKING order="39" place="39" resultid="47112" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46318" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48682" />
                    <RANKING order="2" place="2" resultid="47654" />
                    <RANKING order="3" place="3" resultid="47886" />
                    <RANKING order="4" place="4" resultid="46530" />
                    <RANKING order="5" place="5" resultid="48693" />
                    <RANKING order="6" place="6" resultid="48387" />
                    <RANKING order="7" place="7" resultid="46867" />
                    <RANKING order="8" place="8" resultid="50343" />
                    <RANKING order="9" place="9" resultid="48227" />
                    <RANKING order="10" place="10" resultid="50350" />
                    <RANKING order="11" place="11" resultid="46808" />
                    <RANKING order="12" place="12" resultid="46519" />
                    <RANKING order="13" place="13" resultid="48162" />
                    <RANKING order="14" place="14" resultid="48701" />
                    <RANKING order="15" place="15" resultid="50357" />
                    <RANKING order="16" place="16" resultid="46879" />
                    <RANKING order="17" place="17" resultid="48074" />
                    <RANKING order="18" place="18" resultid="47598" />
                    <RANKING order="19" place="18" resultid="49081" />
                    <RANKING order="20" place="20" resultid="46723" />
                    <RANKING order="21" place="21" resultid="46636" />
                    <RANKING order="22" place="22" resultid="48218" />
                    <RANKING order="23" place="23" resultid="48636" />
                    <RANKING order="24" place="24" resultid="46524" />
                    <RANKING order="25" place="25" resultid="48211" />
                    <RANKING order="26" place="26" resultid="46864" />
                    <RANKING order="27" place="27" resultid="46606" />
                    <RANKING order="28" place="28" resultid="46596" />
                    <RANKING order="29" place="29" resultid="48205" />
                    <RANKING order="30" place="30" resultid="47151" />
                    <RANKING order="31" place="31" resultid="48068" />
                    <RANKING order="32" place="32" resultid="46616" />
                    <RANKING order="33" place="-1" resultid="47147" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46319" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47167" />
                    <RANKING order="2" place="2" resultid="46556" />
                    <RANKING order="3" place="3" resultid="48754" />
                    <RANKING order="4" place="4" resultid="46586" />
                    <RANKING order="5" place="5" resultid="48677" />
                    <RANKING order="6" place="6" resultid="47080" />
                    <RANKING order="7" place="7" resultid="48201" />
                    <RANKING order="8" place="8" resultid="49637" />
                    <RANKING order="9" place="9" resultid="47559" />
                    <RANKING order="10" place="10" resultid="48399" />
                    <RANKING order="11" place="11" resultid="49418" />
                    <RANKING order="12" place="12" resultid="46552" />
                    <RANKING order="13" place="13" resultid="48759" />
                    <RANKING order="14" place="14" resultid="50405" />
                    <RANKING order="15" place="15" resultid="47552" />
                    <RANKING order="16" place="16" resultid="47028" />
                    <RANKING order="17" place="17" resultid="47897" />
                    <RANKING order="18" place="18" resultid="47143" />
                    <RANKING order="19" place="19" resultid="48625" />
                    <RANKING order="20" place="20" resultid="48174" />
                    <RANKING order="21" place="21" resultid="49415" />
                    <RANKING order="22" place="22" resultid="50396" />
                    <RANKING order="23" place="23" resultid="47545" />
                    <RANKING order="24" place="24" resultid="47980" />
                    <RANKING order="25" place="25" resultid="49644" />
                    <RANKING order="26" place="26" resultid="46871" />
                    <RANKING order="27" place="27" resultid="48395" />
                    <RANKING order="28" place="28" resultid="48391" />
                    <RANKING order="29" place="29" resultid="48711" />
                    <RANKING order="30" place="30" resultid="48643" />
                    <RANKING order="31" place="31" resultid="48747" />
                    <RANKING order="32" place="32" resultid="50401" />
                    <RANKING order="33" place="33" resultid="47929" />
                    <RANKING order="34" place="34" resultid="46564" />
                    <RANKING order="35" place="35" resultid="46559" />
                    <RANKING order="36" place="36" resultid="47084" />
                    <RANKING order="37" place="37" resultid="49198" />
                    <RANKING order="38" place="38" resultid="48100" />
                    <RANKING order="39" place="39" resultid="46795" />
                    <RANKING order="40" place="40" resultid="48408" />
                    <RANKING order="41" place="41" resultid="48587" />
                    <RANKING order="42" place="42" resultid="48168" />
                    <RANKING order="43" place="43" resultid="48404" />
                    <RANKING order="44" place="44" resultid="47006" />
                    <RANKING order="45" place="45" resultid="46568" />
                    <RANKING order="46" place="46" resultid="47892" />
                    <RANKING order="47" place="47" resultid="47159" />
                    <RANKING order="48" place="48" resultid="47820" />
                    <RANKING order="49" place="49" resultid="47105" />
                    <RANKING order="50" place="50" resultid="47966" />
                    <RANKING order="51" place="51" resultid="47589" />
                    <RANKING order="52" place="52" resultid="49102" />
                    <RANKING order="53" place="53" resultid="48038" />
                    <RANKING order="54" place="54" resultid="47584" />
                    <RANKING order="55" place="55" resultid="46804" />
                    <RANKING order="56" place="56" resultid="46800" />
                    <RANKING order="57" place="57" resultid="46875" />
                    <RANKING order="58" place="-1" resultid="46461" />
                    <RANKING order="59" place="-1" resultid="47155" />
                    <RANKING order="60" place="-1" resultid="48723" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50663" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50664" daytime="09:03" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50665" daytime="09:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50666" daytime="09:08" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="50667" daytime="09:11" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="50668" daytime="09:13" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="50669" daytime="09:15" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="50670" daytime="09:17" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="50671" daytime="09:19" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="50672" daytime="09:22" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="50673" daytime="09:24" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="50674" daytime="09:26" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="50675" daytime="09:28" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="50676" daytime="09:30" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="50677" daytime="09:31" number="15" order="15" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="44380" daytime="09:33" gender="F" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46320" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="49140" />
                    <RANKING order="2" place="2" resultid="46491" />
                    <RANKING order="3" place="3" resultid="50460" />
                    <RANKING order="4" place="4" resultid="47997" />
                    <RANKING order="5" place="5" resultid="48321" />
                    <RANKING order="6" place="6" resultid="47047" />
                    <RANKING order="7" place="7" resultid="49133" />
                    <RANKING order="8" place="8" resultid="46706" />
                    <RANKING order="9" place="9" resultid="48328" />
                    <RANKING order="10" place="10" resultid="49161" />
                    <RANKING order="11" place="11" resultid="48002" />
                    <RANKING order="12" place="12" resultid="47170" />
                    <RANKING order="13" place="13" resultid="50442" />
                    <RANKING order="14" place="14" resultid="50448" />
                    <RANKING order="15" place="15" resultid="48192" />
                    <RANKING order="16" place="16" resultid="49105" />
                    <RANKING order="17" place="17" resultid="48518" />
                    <RANKING order="18" place="18" resultid="50454" />
                    <RANKING order="19" place="19" resultid="47876" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46321" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46956" />
                    <RANKING order="2" place="2" resultid="47839" />
                    <RANKING order="3" place="3" resultid="50435" />
                    <RANKING order="4" place="4" resultid="50479" />
                    <RANKING order="5" place="5" resultid="47933" />
                    <RANKING order="6" place="6" resultid="48079" />
                    <RANKING order="7" place="7" resultid="48269" />
                    <RANKING order="8" place="8" resultid="49126" />
                    <RANKING order="9" place="9" resultid="48418" />
                    <RANKING order="10" place="10" resultid="46891" />
                    <RANKING order="11" place="11" resultid="48650" />
                    <RANKING order="12" place="12" resultid="48432" />
                    <RANKING order="13" place="13" resultid="49147" />
                    <RANKING order="14" place="14" resultid="48617" />
                    <RANKING order="15" place="15" resultid="47052" />
                    <RANKING order="16" place="16" resultid="49652" />
                    <RANKING order="17" place="17" resultid="47848" />
                    <RANKING order="18" place="18" resultid="48315" />
                    <RANKING order="19" place="19" resultid="46947" />
                    <RANKING order="20" place="20" resultid="48105" />
                    <RANKING order="21" place="21" resultid="48185" />
                    <RANKING order="22" place="22" resultid="46885" />
                    <RANKING order="23" place="23" resultid="48288" />
                    <RANKING order="24" place="24" resultid="48275" />
                    <RANKING order="25" place="25" resultid="46686" />
                    <RANKING order="26" place="26" resultid="48299" />
                    <RANKING order="27" place="27" resultid="48110" />
                    <RANKING order="28" place="28" resultid="48293" />
                    <RANKING order="29" place="29" resultid="48310" />
                    <RANKING order="30" place="30" resultid="48305" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46322" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46961" />
                    <RANKING order="2" place="2" resultid="47043" />
                    <RANKING order="3" place="3" resultid="48427" />
                    <RANKING order="4" place="4" resultid="47677" />
                    <RANKING order="5" place="5" resultid="46739" />
                    <RANKING order="6" place="6" resultid="50424" />
                    <RANKING order="7" place="7" resultid="50410" />
                    <RANKING order="8" place="8" resultid="47039" />
                    <RANKING order="9" place="9" resultid="48592" />
                    <RANKING order="10" place="10" resultid="47180" />
                    <RANKING order="11" place="11" resultid="46933" />
                    <RANKING order="12" place="12" resultid="49119" />
                    <RANKING order="13" place="13" resultid="48280" />
                    <RANKING order="14" place="14" resultid="46696" />
                    <RANKING order="15" place="15" resultid="48529" />
                    <RANKING order="16" place="16" resultid="50417" />
                    <RANKING order="17" place="17" resultid="48284" />
                    <RANKING order="18" place="18" resultid="47184" />
                    <RANKING order="19" place="19" resultid="47613" />
                    <RANKING order="20" place="20" resultid="46676" />
                    <RANKING order="21" place="21" resultid="48536" />
                    <RANKING order="22" place="22" resultid="48657" />
                    <RANKING order="23" place="23" resultid="48180" />
                    <RANKING order="24" place="24" resultid="46656" />
                    <RANKING order="25" place="-1" resultid="49657" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46323" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47670" />
                    <RANKING order="2" place="2" resultid="50467" />
                    <RANKING order="3" place="3" resultid="50472" />
                    <RANKING order="4" place="4" resultid="50485" />
                    <RANKING order="5" place="5" resultid="46574" />
                    <RANKING order="6" place="6" resultid="46882" />
                    <RANKING order="7" place="7" resultid="50431" />
                    <RANKING order="8" place="8" resultid="47566" />
                    <RANKING order="9" place="9" resultid="49112" />
                    <RANKING order="10" place="10" resultid="47088" />
                    <RANKING order="11" place="11" resultid="46666" />
                    <RANKING order="12" place="12" resultid="46926" />
                    <RANKING order="13" place="13" resultid="46733" />
                    <RANKING order="14" place="14" resultid="46817" />
                    <RANKING order="15" place="15" resultid="47175" />
                    <RANKING order="16" place="16" resultid="47902" />
                    <RANKING order="17" place="17" resultid="48763" />
                    <RANKING order="18" place="18" resultid="47125" />
                    <RANKING order="19" place="19" resultid="48042" />
                    <RANKING order="20" place="20" resultid="46812" />
                    <RANKING order="21" place="21" resultid="46498" />
                    <RANKING order="22" place="22" resultid="47907" />
                    <RANKING order="23" place="23" resultid="47855" />
                    <RANKING order="24" place="24" resultid="47869" />
                    <RANKING order="25" place="25" resultid="47131" />
                    <RANKING order="26" place="26" resultid="47862" />
                    <RANKING order="27" place="-1" resultid="46580" />
                    <RANKING order="28" place="-1" resultid="47119" />
                    <RANKING order="29" place="-1" resultid="48423" />
                    <RANKING order="30" place="-1" resultid="49154" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50678" daytime="09:33" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50679" daytime="09:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50680" daytime="09:38" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50681" daytime="09:41" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="50682" daytime="09:43" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="50683" daytime="09:45" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="50684" daytime="09:48" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="50685" daytime="09:50" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="50686" daytime="09:52" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="50687" daytime="09:54" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="50688" daytime="09:56" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="44382" daytime="09:58" gender="M" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46324" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48796" />
                    <RANKING order="2" place="2" resultid="48776" />
                    <RANKING order="3" place="3" resultid="46542" />
                    <RANKING order="4" place="4" resultid="48347" />
                    <RANKING order="5" place="5" resultid="48771" />
                    <RANKING order="6" place="6" resultid="50385" />
                    <RANKING order="7" place="-1" resultid="48733" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46325" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48503" />
                    <RANKING order="2" place="2" resultid="46751" />
                    <RANKING order="3" place="3" resultid="47683" />
                    <RANKING order="4" place="4" resultid="47621" />
                    <RANKING order="5" place="5" resultid="47113" />
                    <RANKING order="6" place="6" resultid="49168" />
                    <RANKING order="7" place="7" resultid="50364" />
                    <RANKING order="8" place="8" resultid="48341" />
                    <RANKING order="9" place="9" resultid="48063" />
                    <RANKING order="10" place="10" resultid="50371" />
                    <RANKING order="11" place="11" resultid="50315" />
                    <RANKING order="12" place="12" resultid="46647" />
                    <RANKING order="13" place="13" resultid="47973" />
                    <RANKING order="14" place="14" resultid="46718" />
                    <RANKING order="15" place="15" resultid="48791" />
                    <RANKING order="16" place="16" resultid="48335" />
                    <RANKING order="17" place="17" resultid="48781" />
                    <RANKING order="18" place="18" resultid="47960" />
                    <RANKING order="19" place="18" resultid="48118" />
                    <RANKING order="20" place="20" resultid="46627" />
                    <RANKING order="21" place="21" resultid="48786" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46326" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46967" />
                    <RANKING order="2" place="2" resultid="46972" />
                    <RANKING order="3" place="3" resultid="46978" />
                    <RANKING order="4" place="4" resultid="50491" />
                    <RANKING order="5" place="5" resultid="48228" />
                    <RANKING order="6" place="5" resultid="48683" />
                    <RANKING order="7" place="7" resultid="46520" />
                    <RANKING order="8" place="8" resultid="48694" />
                    <RANKING order="9" place="9" resultid="47626" />
                    <RANKING order="10" place="10" resultid="48212" />
                    <RANKING order="11" place="11" resultid="46637" />
                    <RANKING order="12" place="12" resultid="48206" />
                    <RANKING order="13" place="13" resultid="46597" />
                    <RANKING order="14" place="14" resultid="46607" />
                    <RANKING order="15" place="15" resultid="46617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46327" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46827" />
                    <RANKING order="2" place="2" resultid="47059" />
                    <RANKING order="3" place="3" resultid="50498" />
                    <RANKING order="4" place="4" resultid="47560" />
                    <RANKING order="5" place="5" resultid="47055" />
                    <RANKING order="6" place="6" resultid="50503" />
                    <RANKING order="7" place="7" resultid="49421" />
                    <RANKING order="8" place="8" resultid="48047" />
                    <RANKING order="9" place="9" resultid="46823" />
                    <RANKING order="10" place="10" resultid="48626" />
                    <RANKING order="11" place="11" resultid="48175" />
                    <RANKING order="12" place="12" resultid="49175" />
                    <RANKING order="13" place="13" resultid="47092" />
                    <RANKING order="14" place="14" resultid="49645" />
                    <RANKING order="15" place="15" resultid="48644" />
                    <RANKING order="16" place="16" resultid="47013" />
                    <RANKING order="17" place="17" resultid="47967" />
                    <RANKING order="18" place="18" resultid="47665" />
                    <RANKING order="19" place="19" resultid="47106" />
                    <RANKING order="20" place="20" resultid="47188" />
                    <RANKING order="21" place="21" resultid="48010" />
                    <RANKING order="22" place="22" resultid="48114" />
                    <RANKING order="23" place="-1" resultid="46565" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50689" daytime="09:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50690" daytime="10:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50691" daytime="10:02" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50692" daytime="10:03" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="50693" daytime="10:05" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="50694" daytime="10:07" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="50695" daytime="10:09" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="44384" daytime="10:10" gender="F" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46328" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47943" />
                    <RANKING order="2" place="2" resultid="48322" />
                    <RANKING order="3" place="3" resultid="47208" />
                    <RANKING order="4" place="4" resultid="50527" />
                    <RANKING order="5" place="5" resultid="46707" />
                    <RANKING order="6" place="6" resultid="48519" />
                    <RANKING order="7" place="7" resultid="47948" />
                    <RANKING order="8" place="8" resultid="47064" />
                    <RANKING order="9" place="9" resultid="47171" />
                    <RANKING order="10" place="10" resultid="50533" />
                    <RANKING order="11" place="11" resultid="47877" />
                    <RANKING order="12" place="12" resultid="50449" />
                    <RANKING order="13" place="13" resultid="46772" />
                    <RANKING order="14" place="14" resultid="47216" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46329" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47938" />
                    <RANKING order="2" place="2" resultid="46983" />
                    <RANKING order="3" place="3" resultid="48816" />
                    <RANKING order="4" place="4" resultid="47840" />
                    <RANKING order="5" place="5" resultid="48080" />
                    <RANKING order="6" place="6" resultid="46767" />
                    <RANKING order="7" place="7" resultid="48436" />
                    <RANKING order="8" place="8" resultid="50509" />
                    <RANKING order="9" place="9" resultid="48354" />
                    <RANKING order="10" place="10" resultid="48359" />
                    <RANKING order="11" place="11" resultid="47212" />
                    <RANKING order="12" place="12" resultid="48801" />
                    <RANKING order="13" place="13" resultid="48661" />
                    <RANKING order="14" place="14" resultid="48544" />
                    <RANKING order="15" place="15" resultid="48294" />
                    <RANKING order="16" place="16" resultid="48306" />
                    <RANKING order="17" place="17" resultid="48300" />
                    <RANKING order="18" place="18" resultid="48311" />
                    <RANKING order="19" place="19" resultid="48811" />
                    <RANKING order="20" place="-1" resultid="46687" />
                    <RANKING order="21" place="-1" resultid="46892" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46330" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46503" />
                    <RANKING order="2" place="2" resultid="48122" />
                    <RANKING order="3" place="3" resultid="49182" />
                    <RANKING order="4" place="4" resultid="47913" />
                    <RANKING order="5" place="5" resultid="46761" />
                    <RANKING order="6" place="6" resultid="49120" />
                    <RANKING order="7" place="7" resultid="47204" />
                    <RANKING order="8" place="8" resultid="48665" />
                    <RANKING order="9" place="9" resultid="46697" />
                    <RANKING order="10" place="10" resultid="46677" />
                    <RANKING order="11" place="-1" resultid="46657" />
                    <RANKING order="12" place="-1" resultid="49658" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46331" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47572" />
                    <RANKING order="2" place="2" resultid="50522" />
                    <RANKING order="3" place="3" resultid="50539" />
                    <RANKING order="4" place="4" resultid="47671" />
                    <RANKING order="5" place="5" resultid="46471" />
                    <RANKING order="6" place="6" resultid="48597" />
                    <RANKING order="7" place="7" resultid="47578" />
                    <RANKING order="8" place="8" resultid="46757" />
                    <RANKING order="9" place="9" resultid="46466" />
                    <RANKING order="10" place="10" resultid="47825" />
                    <RANKING order="11" place="11" resultid="49663" />
                    <RANKING order="12" place="12" resultid="46818" />
                    <RANKING order="13" place="13" resultid="50516" />
                    <RANKING order="14" place="14" resultid="48601" />
                    <RANKING order="15" place="15" resultid="46831" />
                    <RANKING order="16" place="16" resultid="47630" />
                    <RANKING order="17" place="17" resultid="46581" />
                    <RANKING order="18" place="18" resultid="46667" />
                    <RANKING order="19" place="19" resultid="48196" />
                    <RANKING order="20" place="20" resultid="47191" />
                    <RANKING order="21" place="21" resultid="48126" />
                    <RANKING order="22" place="22" resultid="47195" />
                    <RANKING order="23" place="23" resultid="47199" />
                    <RANKING order="24" place="24" resultid="47863" />
                    <RANKING order="25" place="-1" resultid="47120" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50696" daytime="10:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50697" daytime="10:12" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50698" daytime="10:14" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50699" daytime="10:16" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="50700" daytime="10:18" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="50701" daytime="10:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="50702" daytime="10:21" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="50703" daytime="10:23" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="44386" daytime="10:24" gender="M" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46332" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47831" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46333" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46776" />
                    <RANKING order="2" place="2" resultid="48085" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46334" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50351" />
                    <RANKING order="2" place="2" resultid="46525" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46335" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48824" />
                    <RANKING order="2" place="2" resultid="48821" />
                    <RANKING order="3" place="3" resultid="46587" />
                    <RANKING order="4" place="4" resultid="48442" />
                    <RANKING order="5" place="5" resultid="50541" />
                    <RANKING order="6" place="6" resultid="48130" />
                    <RANKING order="7" place="7" resultid="50886" />
                    <RANKING order="8" place="-1" resultid="46560" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50704" daytime="10:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50705" daytime="10:28" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="44388" daytime="10:32" gender="F" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46336" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50546" />
                    <RANKING order="2" place="2" resultid="48329" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46337" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48446" />
                    <RANKING order="2" place="2" resultid="48828" />
                    <RANKING order="3" place="3" resultid="46782" />
                    <RANKING order="4" place="4" resultid="47849" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46338" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50411" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46339" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50549" />
                    <RANKING order="2" place="2" resultid="47856" />
                    <RANKING order="3" place="3" resultid="48134" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50706" daytime="10:32" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="44390" daytime="10:36" gender="M" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46340" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48797" />
                    <RANKING order="2" place="2" resultid="47832" />
                    <RANKING order="3" place="3" resultid="48264" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46341" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46478" />
                    <RANKING order="2" place="2" resultid="46648" />
                    <RANKING order="3" place="3" resultid="48492" />
                    <RANKING order="4" place="4" resultid="46628" />
                    <RANKING order="5" place="5" resultid="50337" />
                    <RANKING order="6" place="6" resultid="48792" />
                    <RANKING order="7" place="7" resultid="49169" />
                    <RANKING order="8" place="8" resultid="48336" />
                    <RANKING order="9" place="9" resultid="48787" />
                    <RANKING order="10" place="-1" resultid="48504" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46342" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46973" />
                    <RANKING order="2" place="2" resultid="48450" />
                    <RANKING order="3" place="3" resultid="48684" />
                    <RANKING order="4" place="4" resultid="46979" />
                    <RANKING order="5" place="5" resultid="46531" />
                    <RANKING order="6" place="6" resultid="48075" />
                    <RANKING order="7" place="7" resultid="46638" />
                    <RANKING order="8" place="8" resultid="48229" />
                    <RANKING order="9" place="9" resultid="48219" />
                    <RANKING order="10" place="10" resultid="46608" />
                    <RANKING order="11" place="11" resultid="46598" />
                    <RANKING order="12" place="12" resultid="48069" />
                    <RANKING order="13" place="13" resultid="46618" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46343" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48822" />
                    <RANKING order="2" place="2" resultid="48669" />
                    <RANKING order="3" place="3" resultid="50567" />
                    <RANKING order="4" place="4" resultid="49638" />
                    <RANKING order="5" place="5" resultid="46872" />
                    <RANKING order="6" place="6" resultid="50561" />
                    <RANKING order="7" place="7" resultid="48454" />
                    <RANKING order="8" place="8" resultid="46836" />
                    <RANKING order="9" place="9" resultid="49199" />
                    <RANKING order="10" place="10" resultid="50555" />
                    <RANKING order="11" place="11" resultid="49646" />
                    <RANKING order="12" place="12" resultid="48138" />
                    <RANKING order="13" place="13" resultid="49176" />
                    <RANKING order="14" place="14" resultid="47007" />
                    <RANKING order="15" place="15" resultid="46805" />
                    <RANKING order="16" place="16" resultid="46569" />
                    <RANKING order="17" place="17" resultid="47107" />
                    <RANKING order="18" place="-1" resultid="48748" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50707" daytime="10:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50708" daytime="10:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50709" daytime="10:44" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50710" daytime="10:48" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="50711" daytime="10:51" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="44392" daytime="10:55" gender="F" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46344" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="49141" />
                    <RANKING order="2" place="2" resultid="48833" />
                    <RANKING order="3" place="3" resultid="46708" />
                    <RANKING order="4" place="4" resultid="50528" />
                    <RANKING order="5" place="5" resultid="48365" />
                    <RANKING order="6" place="6" resultid="48520" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46345" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47841" />
                    <RANKING order="2" place="2" resultid="46984" />
                    <RANKING order="3" place="3" resultid="47939" />
                    <RANKING order="4" place="4" resultid="50480" />
                    <RANKING order="5" place="5" resultid="48270" />
                    <RANKING order="6" place="6" resultid="48437" />
                    <RANKING order="7" place="7" resultid="50510" />
                    <RANKING order="8" place="8" resultid="46768" />
                    <RANKING order="9" place="9" resultid="48618" />
                    <RANKING order="10" place="10" resultid="48817" />
                    <RANKING order="11" place="11" resultid="46688" />
                    <RANKING order="12" place="12" resultid="48186" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46346" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48458" />
                    <RANKING order="2" place="2" resultid="50572" />
                    <RANKING order="3" place="3" resultid="49183" />
                    <RANKING order="4" place="4" resultid="50425" />
                    <RANKING order="5" place="5" resultid="50418" />
                    <RANKING order="6" place="6" resultid="47914" />
                    <RANKING order="7" place="7" resultid="46698" />
                    <RANKING order="8" place="8" resultid="48530" />
                    <RANKING order="9" place="9" resultid="46678" />
                    <RANKING order="10" place="10" resultid="46658" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46347" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50589" />
                    <RANKING order="2" place="2" resultid="46472" />
                    <RANKING order="3" place="3" resultid="50486" />
                    <RANKING order="4" place="4" resultid="50473" />
                    <RANKING order="5" place="5" resultid="50579" />
                    <RANKING order="6" place="6" resultid="46467" />
                    <RANKING order="7" place="7" resultid="46575" />
                    <RANKING order="8" place="8" resultid="47918" />
                    <RANKING order="9" place="9" resultid="50584" />
                    <RANKING order="10" place="10" resultid="46668" />
                    <RANKING order="11" place="11" resultid="47126" />
                    <RANKING order="12" place="12" resultid="46841" />
                    <RANKING order="13" place="13" resultid="47132" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50712" daytime="10:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50713" daytime="10:59" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50714" daytime="11:03" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50715" daytime="11:07" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="50716" daytime="11:11" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="44394" daytime="11:14" gender="M" number="9" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46348" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47021" />
                    <RANKING order="2" place="2" resultid="46899" />
                    <RANKING order="3" place="3" resultid="48257" />
                    <RANKING order="4" place="4" resultid="47986" />
                    <RANKING order="5" place="5" resultid="46513" />
                    <RANKING order="6" place="6" resultid="47219" />
                    <RANKING order="7" place="7" resultid="46485" />
                    <RANKING order="8" place="7" resultid="47595" />
                    <RANKING order="9" place="9" resultid="46920" />
                    <RANKING order="10" place="10" resultid="48348" />
                    <RANKING order="11" place="11" resultid="49096" />
                    <RANKING order="12" place="12" resultid="48512" />
                    <RANKING order="13" place="13" resultid="47992" />
                    <RANKING order="14" place="-1" resultid="48146" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46349" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48091" />
                    <RANKING order="2" place="2" resultid="47688" />
                    <RANKING order="3" place="3" resultid="46906" />
                    <RANKING order="4" place="4" resultid="48142" />
                    <RANKING order="5" place="5" resultid="48463" />
                    <RANKING order="6" place="6" resultid="48838" />
                    <RANKING order="7" place="7" resultid="46913" />
                    <RANKING order="8" place="8" resultid="46988" />
                    <RANKING order="9" place="9" resultid="48086" />
                    <RANKING order="10" place="10" resultid="48371" />
                    <RANKING order="11" place="11" resultid="48493" />
                    <RANKING order="12" place="12" resultid="50378" />
                    <RANKING order="13" place="13" resultid="47925" />
                    <RANKING order="14" place="14" resultid="49089" />
                    <RANKING order="15" place="15" resultid="49075" />
                    <RANKING order="16" place="16" resultid="46858" />
                    <RANKING order="17" place="17" resultid="48738" />
                    <RANKING order="18" place="18" resultid="48342" />
                    <RANKING order="19" place="19" resultid="48241" />
                    <RANKING order="20" place="20" resultid="50391" />
                    <RANKING order="21" place="21" resultid="47223" />
                    <RANKING order="22" place="-1" resultid="48843" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46350" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50344" />
                    <RANKING order="2" place="2" resultid="48163" />
                    <RANKING order="3" place="3" resultid="48220" />
                    <RANKING order="4" place="4" resultid="48702" />
                    <RANKING order="5" place="5" resultid="49082" />
                    <RANKING order="6" place="6" resultid="46992" />
                    <RANKING order="7" place="7" resultid="48637" />
                    <RANKING order="8" place="8" resultid="50492" />
                    <RANKING order="9" place="9" resultid="47638" />
                    <RANKING order="10" place="9" resultid="50358" />
                    <RANKING order="11" place="11" resultid="46508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46351" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47095" />
                    <RANKING order="2" place="2" resultid="48467" />
                    <RANKING order="3" place="3" resultid="47553" />
                    <RANKING order="4" place="4" resultid="46845" />
                    <RANKING order="5" place="5" resultid="48470" />
                    <RANKING order="6" place="6" resultid="48712" />
                    <RANKING order="7" place="7" resultid="47546" />
                    <RANKING order="8" place="8" resultid="47069" />
                    <RANKING order="9" place="9" resultid="47634" />
                    <RANKING order="10" place="10" resultid="47930" />
                    <RANKING order="11" place="11" resultid="48169" />
                    <RANKING order="12" place="12" resultid="48039" />
                    <RANKING order="13" place="13" resultid="47968" />
                    <RANKING order="14" place="14" resultid="46876" />
                    <RANKING order="15" place="15" resultid="50885" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50717" daytime="11:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50718" daytime="11:17" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50719" daytime="11:19" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50720" daytime="11:22" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="50721" daytime="11:24" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="50722" daytime="11:26" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="50723" daytime="11:29" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="44396" daytime="11:31" gender="F" number="10" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46352" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50461" />
                    <RANKING order="2" place="2" resultid="50443" />
                    <RANKING order="3" place="3" resultid="49162" />
                    <RANKING order="4" place="4" resultid="48003" />
                    <RANKING order="5" place="5" resultid="49134" />
                    <RANKING order="6" place="6" resultid="47949" />
                    <RANKING order="7" place="7" resultid="47209" />
                    <RANKING order="8" place="8" resultid="49106" />
                    <RANKING order="9" place="9" resultid="47065" />
                    <RANKING order="10" place="10" resultid="50455" />
                    <RANKING order="11" place="11" resultid="50534" />
                    <RANKING order="12" place="12" resultid="48521" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46353" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50436" />
                    <RANKING order="2" place="2" resultid="49127" />
                    <RANKING order="3" place="3" resultid="47953" />
                    <RANKING order="4" place="4" resultid="48848" />
                    <RANKING order="5" place="5" resultid="46789" />
                    <RANKING order="6" place="6" resultid="48651" />
                    <RANKING order="7" place="7" resultid="48483" />
                    <RANKING order="8" place="8" resultid="46948" />
                    <RANKING order="9" place="9" resultid="48316" />
                    <RANKING order="10" place="10" resultid="48376" />
                    <RANKING order="11" place="11" resultid="48802" />
                    <RANKING order="12" place="12" resultid="48276" />
                    <RANKING order="13" place="13" resultid="48027" />
                    <RANKING order="14" place="14" resultid="48812" />
                    <RANKING order="15" place="15" resultid="48187" />
                    <RANKING order="16" place="16" resultid="46886" />
                    <RANKING order="17" place="17" resultid="48360" />
                    <RANKING order="18" place="-1" resultid="49148" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46354" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50573" />
                    <RANKING order="2" place="2" resultid="46934" />
                    <RANKING order="3" place="3" resultid="48537" />
                    <RANKING order="4" place="4" resultid="48475" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46355" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="49676" />
                    <RANKING order="2" place="2" resultid="48478" />
                    <RANKING order="3" place="3" resultid="49669" />
                    <RANKING order="4" place="4" resultid="50468" />
                    <RANKING order="5" place="5" resultid="50517" />
                    <RANKING order="6" place="6" resultid="49113" />
                    <RANKING order="7" place="7" resultid="48150" />
                    <RANKING order="8" place="8" resultid="48032" />
                    <RANKING order="9" place="9" resultid="46927" />
                    <RANKING order="10" place="10" resultid="48019" />
                    <RANKING order="11" place="11" resultid="48043" />
                    <RANKING order="12" place="12" resultid="48605" />
                    <RANKING order="13" place="13" resultid="47908" />
                    <RANKING order="14" place="14" resultid="47227" />
                    <RANKING order="15" place="15" resultid="48155" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50724" daytime="11:31" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50725" daytime="11:33" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50726" daytime="11:36" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50727" daytime="11:38" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="50728" daytime="11:41" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="44399" daytime="11:43" gender="M" number="11" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46230" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="46231" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48096" />
                    <RANKING order="2" place="2" resultid="46951" />
                    <RANKING order="3" place="3" resultid="48852" />
                    <RANKING order="4" place="4" resultid="48380" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46436" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47000" />
                    <RANKING order="2" place="2" resultid="50598" />
                    <RANKING order="3" place="3" resultid="48379" />
                    <RANKING order="4" place="-1" resultid="47642" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46437" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46849" />
                    <RANKING order="2" place="2" resultid="47530" />
                    <RANKING order="3" place="3" resultid="47076" />
                    <RANKING order="4" place="4" resultid="48674" />
                    <RANKING order="5" place="5" resultid="46850" />
                    <RANKING order="6" place="6" resultid="49188" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50729" daytime="11:43" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50730" daytime="11:49" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="44401" daytime="11:55" gender="F" number="12" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46438" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="49190" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46439" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48853" />
                    <RANKING order="2" place="2" resultid="48381" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46440" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50601" />
                    <RANKING order="2" place="-1" resultid="47001" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46441" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50600" />
                    <RANKING order="2" place="2" resultid="50599" />
                    <RANKING order="3" place="3" resultid="49189" />
                    <RANKING order="4" place="4" resultid="50888" />
                    <RANKING order="5" place="5" resultid="46851" />
                    <RANKING order="6" place="6" resultid="47881" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50731" daytime="11:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50887" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2021-05-28" daytime="13:15" endtime="17:37" number="2" warmupfrom="12:15">
          <EVENTS>
            <EVENT eventid="44403" daytime="13:15" gender="M" number="13" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46356" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46900" />
                    <RANKING order="2" place="2" resultid="47833" />
                    <RANKING order="3" place="3" resultid="47022" />
                    <RANKING order="4" place="4" resultid="47662" />
                    <RANKING order="5" place="5" resultid="48258" />
                    <RANKING order="6" place="6" resultid="46486" />
                    <RANKING order="7" place="7" resultid="46730" />
                    <RANKING order="8" place="8" resultid="46921" />
                    <RANKING order="9" place="9" resultid="49097" />
                    <RANKING order="10" place="-1" resultid="48734" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46357" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48092" />
                    <RANKING order="2" place="2" resultid="46479" />
                    <RANKING order="3" place="3" resultid="48057" />
                    <RANKING order="4" place="4" resultid="46649" />
                    <RANKING order="5" place="5" resultid="50316" />
                    <RANKING order="6" place="6" resultid="46914" />
                    <RANKING order="7" place="7" resultid="46907" />
                    <RANKING order="8" place="8" resultid="46629" />
                    <RANKING order="9" place="9" resultid="47961" />
                    <RANKING order="10" place="10" resultid="50322" />
                    <RANKING order="11" place="11" resultid="47974" />
                    <RANKING order="12" place="12" resultid="46719" />
                    <RANKING order="13" place="13" resultid="49076" />
                    <RANKING order="14" place="14" resultid="50338" />
                    <RANKING order="15" place="15" resultid="50331" />
                    <RANKING order="16" place="16" resultid="48236" />
                    <RANKING order="17" place="17" resultid="46859" />
                    <RANKING order="18" place="18" resultid="50392" />
                    <RANKING order="19" place="19" resultid="48251" />
                    <RANKING order="20" place="20" resultid="49090" />
                    <RANKING order="21" place="21" resultid="47604" />
                    <RANKING order="22" place="22" resultid="47101" />
                    <RANKING order="23" place="-1" resultid="48494" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46358" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47655" />
                    <RANKING order="2" place="2" resultid="48685" />
                    <RANKING order="3" place="3" resultid="48451" />
                    <RANKING order="4" place="4" resultid="46532" />
                    <RANKING order="5" place="5" resultid="46809" />
                    <RANKING order="6" place="6" resultid="48703" />
                    <RANKING order="7" place="7" resultid="50359" />
                    <RANKING order="8" place="8" resultid="48695" />
                    <RANKING order="9" place="9" resultid="46639" />
                    <RANKING order="10" place="10" resultid="50352" />
                    <RANKING order="11" place="11" resultid="46724" />
                    <RANKING order="12" place="12" resultid="46609" />
                    <RANKING order="13" place="13" resultid="46599" />
                    <RANKING order="14" place="14" resultid="46619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46359" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46588" />
                    <RANKING order="2" place="2" resultid="48755" />
                    <RANKING order="3" place="3" resultid="48678" />
                    <RANKING order="4" place="4" resultid="48443" />
                    <RANKING order="5" place="5" resultid="50406" />
                    <RANKING order="6" place="6" resultid="47029" />
                    <RANKING order="7" place="7" resultid="49639" />
                    <RANKING order="8" place="8" resultid="50562" />
                    <RANKING order="9" place="9" resultid="50397" />
                    <RANKING order="10" place="10" resultid="48400" />
                    <RANKING order="11" place="11" resultid="48670" />
                    <RANKING order="12" place="12" resultid="47554" />
                    <RANKING order="13" place="13" resultid="47981" />
                    <RANKING order="14" place="14" resultid="48396" />
                    <RANKING order="15" place="15" resultid="49419" />
                    <RANKING order="16" place="16" resultid="47547" />
                    <RANKING order="17" place="17" resultid="50556" />
                    <RANKING order="18" place="18" resultid="48392" />
                    <RANKING order="19" place="19" resultid="47821" />
                    <RANKING order="20" place="20" resultid="48405" />
                    <RANKING order="21" place="21" resultid="47666" />
                    <RANKING order="22" place="22" resultid="47590" />
                    <RANKING order="23" place="23" resultid="48749" />
                    <RANKING order="24" place="24" resultid="47008" />
                    <RANKING order="25" place="25" resultid="46801" />
                    <RANKING order="26" place="26" resultid="46570" />
                    <RANKING order="27" place="27" resultid="49895" />
                    <RANKING order="28" place="28" resultid="48040" />
                    <RANKING order="29" place="29" resultid="47585" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50732" daytime="13:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50733" daytime="13:19" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50734" daytime="13:23" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50735" daytime="13:26" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="50736" daytime="13:30" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="50737" daytime="13:33" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="50738" daytime="13:36" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="50739" daytime="13:39" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="44405" daytime="13:42" gender="F" number="14" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46360" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="49142" />
                    <RANKING order="2" place="2" resultid="46492" />
                    <RANKING order="3" place="3" resultid="48330" />
                    <RANKING order="4" place="4" resultid="49163" />
                    <RANKING order="5" place="5" resultid="47998" />
                    <RANKING order="6" place="6" resultid="48323" />
                    <RANKING order="7" place="7" resultid="47048" />
                    <RANKING order="8" place="8" resultid="46709" />
                    <RANKING order="9" place="9" resultid="49135" />
                    <RANKING order="10" place="10" resultid="49107" />
                    <RANKING order="11" place="-1" resultid="50879" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46361" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47842" />
                    <RANKING order="2" place="2" resultid="50437" />
                    <RANKING order="3" place="3" resultid="48829" />
                    <RANKING order="4" place="4" resultid="50481" />
                    <RANKING order="5" place="5" resultid="46957" />
                    <RANKING order="6" place="6" resultid="48419" />
                    <RANKING order="7" place="7" resultid="49128" />
                    <RANKING order="8" place="8" resultid="48619" />
                    <RANKING order="9" place="9" resultid="46949" />
                    <RANKING order="10" place="10" resultid="46689" />
                    <RANKING order="11" place="11" resultid="48289" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46362" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48459" />
                    <RANKING order="2" place="2" resultid="48428" />
                    <RANKING order="3" place="3" resultid="46962" />
                    <RANKING order="4" place="4" resultid="46740" />
                    <RANKING order="5" place="5" resultid="47040" />
                    <RANKING order="6" place="6" resultid="48281" />
                    <RANKING order="7" place="7" resultid="46699" />
                    <RANKING order="8" place="8" resultid="50426" />
                    <RANKING order="9" place="9" resultid="50412" />
                    <RANKING order="10" place="10" resultid="50419" />
                    <RANKING order="11" place="11" resultid="46935" />
                    <RANKING order="12" place="12" resultid="46679" />
                    <RANKING order="13" place="13" resultid="46659" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46363" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50590" />
                    <RANKING order="2" place="2" resultid="47672" />
                    <RANKING order="3" place="3" resultid="47567" />
                    <RANKING order="4" place="4" resultid="50487" />
                    <RANKING order="5" place="5" resultid="50432" />
                    <RANKING order="6" place="6" resultid="50474" />
                    <RANKING order="7" place="7" resultid="50550" />
                    <RANKING order="8" place="8" resultid="46669" />
                    <RANKING order="9" place="9" resultid="46734" />
                    <RANKING order="10" place="10" resultid="49156" />
                    <RANKING order="11" place="11" resultid="46819" />
                    <RANKING order="12" place="12" resultid="46928" />
                    <RANKING order="13" place="13" resultid="47870" />
                    <RANKING order="14" place="14" resultid="47133" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50740" daytime="13:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50741" daytime="13:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50742" daytime="13:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50743" daytime="13:54" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="50744" daytime="13:57" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="44407" daytime="14:00" gender="M" number="15" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46364" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48798" />
                    <RANKING order="2" place="2" resultid="48777" />
                    <RANKING order="3" place="3" resultid="46543" />
                    <RANKING order="4" place="4" resultid="47987" />
                    <RANKING order="5" place="5" resultid="48349" />
                    <RANKING order="6" place="6" resultid="50386" />
                    <RANKING order="7" place="7" resultid="49098" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46365" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48505" />
                    <RANKING order="2" place="2" resultid="46752" />
                    <RANKING order="3" place="3" resultid="47684" />
                    <RANKING order="4" place="4" resultid="47114" />
                    <RANKING order="5" place="5" resultid="47622" />
                    <RANKING order="6" place="6" resultid="50372" />
                    <RANKING order="7" place="7" resultid="48343" />
                    <RANKING order="8" place="8" resultid="50365" />
                    <RANKING order="9" place="9" resultid="49170" />
                    <RANKING order="10" place="10" resultid="48064" />
                    <RANKING order="11" place="11" resultid="50327" />
                    <RANKING order="12" place="12" resultid="48793" />
                    <RANKING order="13" place="13" resultid="47975" />
                    <RANKING order="14" place="14" resultid="48337" />
                    <RANKING order="15" place="15" resultid="48739" />
                    <RANKING order="16" place="16" resultid="48788" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46366" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46980" />
                    <RANKING order="2" place="2" resultid="50493" />
                    <RANKING order="3" place="3" resultid="46974" />
                    <RANKING order="4" place="4" resultid="48230" />
                    <RANKING order="5" place="5" resultid="48686" />
                    <RANKING order="6" place="6" resultid="47627" />
                    <RANKING order="7" place="7" resultid="48213" />
                    <RANKING order="8" place="8" resultid="48070" />
                    <RANKING order="9" place="9" resultid="48207" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46367" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50568" />
                    <RANKING order="2" place="2" resultid="47561" />
                    <RANKING order="3" place="3" resultid="47056" />
                    <RANKING order="4" place="4" resultid="50504" />
                    <RANKING order="5" place="5" resultid="50499" />
                    <RANKING order="6" place="6" resultid="46824" />
                    <RANKING order="7" place="7" resultid="49177" />
                    <RANKING order="8" place="8" resultid="47093" />
                    <RANKING order="9" place="9" resultid="48455" />
                    <RANKING order="10" place="10" resultid="49197" />
                    <RANKING order="11" place="11" resultid="49647" />
                    <RANKING order="12" place="12" resultid="49422" />
                    <RANKING order="13" place="13" resultid="50402" />
                    <RANKING order="14" place="14" resultid="49896" />
                    <RANKING order="15" place="15" resultid="48645" />
                    <RANKING order="16" place="16" resultid="48139" />
                    <RANKING order="17" place="17" resultid="47969" />
                    <RANKING order="18" place="18" resultid="47108" />
                    <RANKING order="19" place="19" resultid="47014" />
                    <RANKING order="20" place="20" resultid="48011" />
                    <RANKING order="21" place="21" resultid="50889" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50745" daytime="14:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50746" daytime="14:03" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50747" daytime="14:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50748" daytime="14:08" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="50749" daytime="14:11" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="50750" daytime="14:13" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="44409" daytime="14:15" gender="F" number="16" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46368" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48324" />
                    <RANKING order="2" place="2" resultid="47944" />
                    <RANKING order="3" place="3" resultid="50529" />
                    <RANKING order="4" place="4" resultid="48366" />
                    <RANKING order="5" place="5" resultid="47950" />
                    <RANKING order="6" place="6" resultid="47878" />
                    <RANKING order="7" place="7" resultid="48522" />
                    <RANKING order="8" place="8" resultid="50450" />
                    <RANKING order="9" place="9" resultid="50535" />
                    <RANKING order="10" place="10" resultid="46773" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46369" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48447" />
                    <RANKING order="2" place="2" resultid="47940" />
                    <RANKING order="3" place="3" resultid="46985" />
                    <RANKING order="4" place="4" resultid="48818" />
                    <RANKING order="5" place="5" resultid="46769" />
                    <RANKING order="6" place="6" resultid="48081" />
                    <RANKING order="7" place="7" resultid="48438" />
                    <RANKING order="8" place="8" resultid="50511" />
                    <RANKING order="9" place="9" resultid="48355" />
                    <RANKING order="10" place="10" resultid="48361" />
                    <RANKING order="11" place="11" resultid="48662" />
                    <RANKING order="12" place="12" resultid="48803" />
                    <RANKING order="13" place="13" resultid="48295" />
                    <RANKING order="14" place="14" resultid="48545" />
                    <RANKING order="15" place="15" resultid="48307" />
                    <RANKING order="16" place="16" resultid="48312" />
                    <RANKING order="17" place="17" resultid="48813" />
                    <RANKING order="18" place="-1" resultid="47843" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46370" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="49184" />
                    <RANKING order="2" place="2" resultid="47915" />
                    <RANKING order="3" place="3" resultid="46504" />
                    <RANKING order="4" place="4" resultid="48123" />
                    <RANKING order="5" place="5" resultid="46762" />
                    <RANKING order="6" place="6" resultid="47205" />
                    <RANKING order="7" place="7" resultid="48666" />
                    <RANKING order="8" place="-1" resultid="49659" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46371" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47573" />
                    <RANKING order="2" place="2" resultid="50523" />
                    <RANKING order="3" place="3" resultid="46473" />
                    <RANKING order="4" place="4" resultid="46758" />
                    <RANKING order="5" place="5" resultid="47579" />
                    <RANKING order="6" place="6" resultid="49664" />
                    <RANKING order="7" place="7" resultid="48598" />
                    <RANKING order="8" place="8" resultid="46468" />
                    <RANKING order="9" place="9" resultid="48602" />
                    <RANKING order="10" place="10" resultid="47826" />
                    <RANKING order="11" place="11" resultid="47919" />
                    <RANKING order="12" place="12" resultid="46832" />
                    <RANKING order="13" place="13" resultid="47631" />
                    <RANKING order="14" place="14" resultid="47864" />
                    <RANKING order="15" place="-1" resultid="47121" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50751" daytime="14:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50752" daytime="14:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50753" daytime="14:21" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50754" daytime="14:24" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="50755" daytime="14:26" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="50756" daytime="14:29" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="44411" daytime="14:31" gender="M" number="17" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46372" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46901" />
                    <RANKING order="2" place="2" resultid="47023" />
                    <RANKING order="3" place="3" resultid="47834" />
                    <RANKING order="4" place="4" resultid="48772" />
                    <RANKING order="5" place="5" resultid="48778" />
                    <RANKING order="6" place="6" resultid="46544" />
                    <RANKING order="7" place="7" resultid="47220" />
                    <RANKING order="8" place="8" resultid="48259" />
                    <RANKING order="9" place="9" resultid="48265" />
                    <RANKING order="10" place="10" resultid="50873" />
                    <RANKING order="11" place="11" resultid="46922" />
                    <RANKING order="12" place="12" resultid="47993" />
                    <RANKING order="13" place="13" resultid="50387" />
                    <RANKING order="14" place="14" resultid="48513" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46373" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47689" />
                    <RANKING order="2" place="2" resultid="48743" />
                    <RANKING order="3" place="3" resultid="46753" />
                    <RANKING order="4" place="4" resultid="47164" />
                    <RANKING order="5" place="5" resultid="50317" />
                    <RANKING order="6" place="6" resultid="48728" />
                    <RANKING order="7" place="7" resultid="46908" />
                    <RANKING order="8" place="8" resultid="48087" />
                    <RANKING order="9" place="9" resultid="46915" />
                    <RANKING order="10" place="10" resultid="46989" />
                    <RANKING order="11" place="11" resultid="46650" />
                    <RANKING order="12" place="12" resultid="50366" />
                    <RANKING order="13" place="13" resultid="48495" />
                    <RANKING order="14" place="13" resultid="50323" />
                    <RANKING order="15" place="15" resultid="47976" />
                    <RANKING order="16" place="16" resultid="48414" />
                    <RANKING order="17" place="17" resultid="48632" />
                    <RANKING order="18" place="18" resultid="48506" />
                    <RANKING order="19" place="19" resultid="46630" />
                    <RANKING order="20" place="20" resultid="48058" />
                    <RANKING order="21" place="21" resultid="49077" />
                    <RANKING order="22" place="22" resultid="46860" />
                    <RANKING order="23" place="23" resultid="47962" />
                    <RANKING order="24" place="24" resultid="47035" />
                    <RANKING order="25" place="25" resultid="50328" />
                    <RANKING order="26" place="26" resultid="49171" />
                    <RANKING order="27" place="27" resultid="48119" />
                    <RANKING order="28" place="28" resultid="50379" />
                    <RANKING order="29" place="29" resultid="50339" />
                    <RANKING order="30" place="30" resultid="48338" />
                    <RANKING order="31" place="31" resultid="47224" />
                    <RANKING order="32" place="32" resultid="48782" />
                    <RANKING order="33" place="-1" resultid="47926" />
                    <RANKING order="34" place="-1" resultid="48237" />
                    <RANKING order="35" place="-1" resultid="48844" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46374" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46968" />
                    <RANKING order="2" place="2" resultid="50353" />
                    <RANKING order="3" place="3" resultid="47656" />
                    <RANKING order="4" place="4" resultid="47887" />
                    <RANKING order="5" place="5" resultid="48388" />
                    <RANKING order="6" place="6" resultid="48696" />
                    <RANKING order="7" place="7" resultid="47599" />
                    <RANKING order="8" place="8" resultid="46533" />
                    <RANKING order="9" place="9" resultid="46868" />
                    <RANKING order="10" place="10" resultid="46521" />
                    <RANKING order="11" place="10" resultid="48704" />
                    <RANKING order="12" place="12" resultid="48687" />
                    <RANKING order="13" place="13" resultid="46993" />
                    <RANKING order="14" place="14" resultid="49083" />
                    <RANKING order="15" place="15" resultid="46526" />
                    <RANKING order="16" place="16" resultid="46880" />
                    <RANKING order="17" place="17" resultid="50345" />
                    <RANKING order="18" place="18" resultid="48638" />
                    <RANKING order="19" place="19" resultid="46610" />
                    <RANKING order="20" place="20" resultid="46640" />
                    <RANKING order="21" place="21" resultid="46865" />
                    <RANKING order="22" place="22" resultid="47152" />
                    <RANKING order="23" place="23" resultid="46725" />
                    <RANKING order="24" place="24" resultid="46600" />
                    <RANKING order="25" place="25" resultid="46620" />
                    <RANKING order="26" place="26" resultid="48071" />
                    <RANKING order="27" place="27" resultid="50494" />
                    <RANKING order="28" place="-1" resultid="47148" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46375" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46462" />
                    <RANKING order="2" place="2" resultid="47081" />
                    <RANKING order="3" place="3" resultid="49640" />
                    <RANKING order="4" place="4" resultid="48679" />
                    <RANKING order="5" place="5" resultid="47074" />
                    <RANKING order="6" place="6" resultid="48756" />
                    <RANKING order="7" place="7" resultid="48176" />
                    <RANKING order="8" place="8" resultid="50594" />
                    <RANKING order="9" place="9" resultid="50569" />
                    <RANKING order="10" place="10" resultid="47562" />
                    <RANKING order="11" place="11" resultid="48627" />
                    <RANKING order="12" place="12" resultid="48750" />
                    <RANKING order="13" place="13" resultid="46589" />
                    <RANKING order="14" place="14" resultid="47030" />
                    <RANKING order="15" place="15" resultid="48760" />
                    <RANKING order="16" place="16" resultid="49416" />
                    <RANKING order="17" place="17" resultid="46553" />
                    <RANKING order="18" place="17" resultid="47144" />
                    <RANKING order="19" place="19" resultid="48401" />
                    <RANKING order="20" place="20" resultid="49648" />
                    <RANKING order="21" place="21" resultid="47070" />
                    <RANKING order="22" place="22" resultid="47060" />
                    <RANKING order="23" place="23" resultid="50557" />
                    <RANKING order="24" place="24" resultid="48101" />
                    <RANKING order="25" place="25" resultid="48671" />
                    <RANKING order="26" place="26" resultid="48409" />
                    <RANKING order="27" place="27" resultid="48170" />
                    <RANKING order="28" place="28" resultid="47898" />
                    <RANKING order="29" place="29" resultid="47548" />
                    <RANKING order="30" place="30" resultid="50563" />
                    <RANKING order="31" place="31" resultid="46873" />
                    <RANKING order="32" place="32" resultid="50542" />
                    <RANKING order="33" place="33" resultid="48048" />
                    <RANKING order="34" place="34" resultid="50505" />
                    <RANKING order="35" place="35" resultid="46837" />
                    <RANKING order="36" place="36" resultid="47009" />
                    <RANKING order="37" place="36" resultid="48588" />
                    <RANKING order="38" place="38" resultid="48646" />
                    <RANKING order="39" place="39" resultid="49178" />
                    <RANKING order="40" place="40" resultid="47160" />
                    <RANKING order="41" place="41" resultid="48131" />
                    <RANKING order="42" place="42" resultid="47591" />
                    <RANKING order="43" place="43" resultid="47015" />
                    <RANKING order="44" place="44" resultid="47586" />
                    <RANKING order="45" place="45" resultid="47232" />
                    <RANKING order="46" place="-1" resultid="47156" />
                    <RANKING order="47" place="-1" resultid="47893" />
                    <RANKING order="48" place="-1" resultid="48051" />
                    <RANKING order="49" place="-1" resultid="48724" />
                    <RANKING order="50" place="-1" resultid="50893" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50757" daytime="14:31" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50758" daytime="14:33" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50759" daytime="14:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50760" daytime="14:37" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="50761" daytime="14:38" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="50762" daytime="14:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="50763" daytime="14:42" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="50764" daytime="14:44" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="50765" daytime="14:45" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="50766" daytime="14:47" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="50767" daytime="14:48" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="50768" daytime="14:50" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="50769" daytime="14:51" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="50894" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="44413" daytime="14:53" gender="F" number="18" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46376" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50462" />
                    <RANKING order="2" place="2" resultid="48004" />
                    <RANKING order="3" place="3" resultid="47945" />
                    <RANKING order="4" place="4" resultid="46710" />
                    <RANKING order="5" place="5" resultid="48331" />
                    <RANKING order="6" place="6" resultid="49108" />
                    <RANKING order="7" place="7" resultid="48193" />
                    <RANKING order="8" place="8" resultid="49136" />
                    <RANKING order="9" place="9" resultid="49164" />
                    <RANKING order="10" place="10" resultid="48367" />
                    <RANKING order="11" place="11" resultid="48523" />
                    <RANKING order="12" place="12" resultid="47049" />
                    <RANKING order="13" place="13" resultid="47172" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46377" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46997" />
                    <RANKING order="2" place="2" resultid="46958" />
                    <RANKING order="3" place="3" resultid="47934" />
                    <RANKING order="4" place="4" resultid="48652" />
                    <RANKING order="5" place="5" resultid="50482" />
                    <RANKING order="6" place="6" resultid="47844" />
                    <RANKING order="7" place="7" resultid="48830" />
                    <RANKING order="8" place="8" resultid="48271" />
                    <RANKING order="9" place="9" resultid="48849" />
                    <RANKING order="10" place="10" resultid="48082" />
                    <RANKING order="11" place="11" resultid="48106" />
                    <RANKING order="12" place="12" resultid="48486" />
                    <RANKING order="13" place="13" resultid="50512" />
                    <RANKING order="14" place="14" resultid="49149" />
                    <RANKING order="15" place="15" resultid="49653" />
                    <RANKING order="16" place="16" resultid="46950" />
                    <RANKING order="17" place="17" resultid="46893" />
                    <RANKING order="18" place="18" resultid="48439" />
                    <RANKING order="19" place="19" resultid="47213" />
                    <RANKING order="20" place="20" resultid="47850" />
                    <RANKING order="21" place="21" resultid="48620" />
                    <RANKING order="22" place="22" resultid="48317" />
                    <RANKING order="23" place="23" resultid="48301" />
                    <RANKING order="24" place="24" resultid="48188" />
                    <RANKING order="25" place="25" resultid="48277" />
                    <RANKING order="26" place="26" resultid="46887" />
                    <RANKING order="27" place="27" resultid="48028" />
                    <RANKING order="28" place="28" resultid="48111" />
                    <RANKING order="29" place="29" resultid="48356" />
                    <RANKING order="30" place="30" resultid="46690" />
                    <RANKING order="31" place="31" resultid="48546" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46378" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46963" />
                    <RANKING order="2" place="2" resultid="50427" />
                    <RANKING order="3" place="3" resultid="46537" />
                    <RANKING order="4" place="4" resultid="50413" />
                    <RANKING order="5" place="5" resultid="47181" />
                    <RANKING order="6" place="6" resultid="47678" />
                    <RANKING order="7" place="7" resultid="49185" />
                    <RANKING order="8" place="8" resultid="46763" />
                    <RANKING order="9" place="9" resultid="48531" />
                    <RANKING order="10" place="10" resultid="46936" />
                    <RANKING order="11" place="11" resultid="48593" />
                    <RANKING order="12" place="12" resultid="48181" />
                    <RANKING order="13" place="13" resultid="48285" />
                    <RANKING order="14" place="14" resultid="48658" />
                    <RANKING order="15" place="15" resultid="47185" />
                    <RANKING order="16" place="16" resultid="46700" />
                    <RANKING order="17" place="17" resultid="46505" />
                    <RANKING order="18" place="18" resultid="47614" />
                    <RANKING order="19" place="19" resultid="46680" />
                    <RANKING order="20" place="20" resultid="46660" />
                    <RANKING order="21" place="-1" resultid="48538" />
                    <RANKING order="22" place="-1" resultid="49121" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46379" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="49670" />
                    <RANKING order="2" place="2" resultid="48479" />
                    <RANKING order="3" place="3" resultid="46576" />
                    <RANKING order="4" place="4" resultid="47235" />
                    <RANKING order="5" place="5" resultid="50475" />
                    <RANKING order="6" place="6" resultid="47673" />
                    <RANKING order="7" place="7" resultid="50524" />
                    <RANKING order="8" place="8" resultid="50591" />
                    <RANKING order="9" place="9" resultid="49665" />
                    <RANKING order="10" place="10" resultid="47574" />
                    <RANKING order="11" place="11" resultid="49114" />
                    <RANKING order="12" place="12" resultid="47903" />
                    <RANKING order="13" place="13" resultid="46820" />
                    <RANKING order="14" place="14" resultid="47176" />
                    <RANKING order="15" place="15" resultid="48764" />
                    <RANKING order="16" place="16" resultid="46670" />
                    <RANKING order="17" place="17" resultid="48020" />
                    <RANKING order="18" place="18" resultid="47127" />
                    <RANKING order="19" place="19" resultid="46929" />
                    <RANKING order="20" place="20" resultid="47920" />
                    <RANKING order="21" place="21" resultid="48135" />
                    <RANKING order="22" place="22" resultid="47857" />
                    <RANKING order="23" place="23" resultid="46833" />
                    <RANKING order="24" place="24" resultid="48156" />
                    <RANKING order="25" place="25" resultid="46813" />
                    <RANKING order="26" place="26" resultid="46842" />
                    <RANKING order="27" place="27" resultid="47909" />
                    <RANKING order="28" place="28" resultid="47196" />
                    <RANKING order="29" place="29" resultid="47865" />
                    <RANKING order="30" place="30" resultid="47871" />
                    <RANKING order="31" place="31" resultid="47200" />
                    <RANKING order="32" place="-1" resultid="48424" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50770" daytime="14:53" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50771" daytime="14:54" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50772" daytime="14:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50773" daytime="14:58" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="50774" daytime="15:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="50775" daytime="15:02" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="50776" daytime="15:03" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="50777" daytime="15:05" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="50778" daytime="15:07" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="50779" daytime="15:08" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="44415" daytime="15:10" gender="M" number="19" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46380" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47024" />
                    <RANKING order="2" place="2" resultid="46514" />
                    <RANKING order="3" place="3" resultid="48350" />
                    <RANKING order="4" place="-1" resultid="48147" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46381" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47690" />
                    <RANKING order="2" place="2" resultid="48093" />
                    <RANKING order="3" place="3" resultid="48464" />
                    <RANKING order="4" place="4" resultid="50373" />
                    <RANKING order="5" place="5" resultid="48839" />
                    <RANKING order="6" place="6" resultid="48143" />
                    <RANKING order="7" place="7" resultid="50380" />
                    <RANKING order="8" place="8" resultid="48496" />
                    <RANKING order="9" place="9" resultid="49091" />
                    <RANKING order="10" place="10" resultid="48372" />
                    <RANKING order="11" place="11" resultid="46631" />
                    <RANKING order="12" place="12" resultid="46651" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46382" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48705" />
                    <RANKING order="2" place="2" resultid="48221" />
                    <RANKING order="3" place="3" resultid="48164" />
                    <RANKING order="4" place="4" resultid="50346" />
                    <RANKING order="5" place="5" resultid="48639" />
                    <RANKING order="6" place="6" resultid="49084" />
                    <RANKING order="7" place="7" resultid="46509" />
                    <RANKING order="8" place="8" resultid="46641" />
                    <RANKING order="9" place="9" resultid="47639" />
                    <RANKING order="10" place="10" resultid="46611" />
                    <RANKING order="11" place="11" resultid="46601" />
                    <RANKING order="12" place="12" resultid="46621" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46383" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48826" />
                    <RANKING order="2" place="2" resultid="47096" />
                    <RANKING order="3" place="3" resultid="47555" />
                    <RANKING order="4" place="4" resultid="48471" />
                    <RANKING order="5" place="5" resultid="46846" />
                    <RANKING order="6" place="6" resultid="50543" />
                    <RANKING order="7" place="7" resultid="48713" />
                    <RANKING order="8" place="8" resultid="49071" />
                    <RANKING order="9" place="9" resultid="47635" />
                    <RANKING order="10" place="10" resultid="47931" />
                    <RANKING order="11" place="11" resultid="46796" />
                    <RANKING order="12" place="12" resultid="46877" />
                    <RANKING order="13" place="13" resultid="48115" />
                    <RANKING order="14" place="14" resultid="50890" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50780" daytime="15:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50781" daytime="15:13" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50782" daytime="15:17" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50783" daytime="15:21" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="50784" daytime="15:25" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="44417" daytime="15:28" gender="F" number="20" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46384" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="49143" />
                    <RANKING order="2" place="2" resultid="48834" />
                    <RANKING order="3" place="3" resultid="50463" />
                    <RANKING order="4" place="4" resultid="46711" />
                    <RANKING order="5" place="5" resultid="50444" />
                    <RANKING order="6" place="6" resultid="48005" />
                    <RANKING order="7" place="7" resultid="50456" />
                    <RANKING order="8" place="-1" resultid="48524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46385" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="49129" />
                    <RANKING order="2" place="2" resultid="50438" />
                    <RANKING order="3" place="3" resultid="47954" />
                    <RANKING order="4" place="4" resultid="46790" />
                    <RANKING order="5" place="5" resultid="48850" />
                    <RANKING order="6" place="6" resultid="49150" />
                    <RANKING order="7" place="7" resultid="48377" />
                    <RANKING order="8" place="8" resultid="46691" />
                    <RANKING order="9" place="9" resultid="48107" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46386" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50574" />
                    <RANKING order="2" place="2" resultid="46701" />
                    <RANKING order="3" place="3" resultid="48539" />
                    <RANKING order="4" place="4" resultid="46681" />
                    <RANKING order="5" place="5" resultid="46661" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46387" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="49677" />
                    <RANKING order="2" place="2" resultid="49671" />
                    <RANKING order="3" place="3" resultid="50580" />
                    <RANKING order="4" place="4" resultid="50518" />
                    <RANKING order="5" place="5" resultid="50585" />
                    <RANKING order="6" place="6" resultid="49115" />
                    <RANKING order="7" place="7" resultid="48151" />
                    <RANKING order="8" place="8" resultid="48033" />
                    <RANKING order="9" place="9" resultid="46671" />
                    <RANKING order="10" place="10" resultid="48021" />
                    <RANKING order="11" place="11" resultid="48606" />
                    <RANKING order="12" place="12" resultid="46499" />
                    <RANKING order="13" place="13" resultid="47228" />
                    <RANKING order="14" place="14" resultid="48157" />
                    <RANKING order="15" place="15" resultid="48127" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50785" daytime="15:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50786" daytime="15:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50787" daytime="15:37" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50788" daytime="15:41" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="46285" daytime="15:45" gender="M" number="21" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46388" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="46389" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46480" />
                    <RANKING order="2" place="2" resultid="46778" />
                    <RANKING order="3" place="3" resultid="50332" />
                    <RANKING order="4" place="4" resultid="48252" />
                    <RANKING order="5" place="5" resultid="48246" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46390" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48076" />
                    <RANKING order="2" place="2" resultid="48222" />
                    <RANKING order="3" place="3" resultid="48214" />
                    <RANKING order="4" place="4" resultid="48208" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46391" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46590" />
                    <RANKING order="2" place="2" resultid="47085" />
                    <RANKING order="3" place="3" resultid="50398" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50789" daytime="15:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50790" daytime="16:04" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="46287" daytime="16:24" gender="F" number="22" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46392" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46493" />
                    <RANKING order="2" place="2" resultid="46547" />
                    <RANKING order="3" place="3" resultid="48325" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46393" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46785" />
                    <RANKING order="2" place="2" resultid="48433" />
                    <RANKING order="3" place="3" resultid="48487" />
                    <RANKING order="4" place="4" resultid="48420" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46394" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48460" />
                    <RANKING order="2" place="2" resultid="50575" />
                    <RANKING order="3" place="3" resultid="50420" />
                    <RANKING order="4" place="-1" resultid="46741" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46395" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47089" />
                    <RANKING order="2" place="2" resultid="47568" />
                    <RANKING order="3" place="3" resultid="46735" />
                    <RANKING order="4" place="4" resultid="50551" />
                    <RANKING order="5" place="5" resultid="47872" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50791" daytime="16:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50792" daytime="16:38" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="46289" daytime="16:51" gender="M" number="23" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46442" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="46443" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48097" />
                    <RANKING order="2" place="2" resultid="48854" />
                    <RANKING order="3" place="3" resultid="46952" />
                    <RANKING order="4" place="4" resultid="48383" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46444" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47002" />
                    <RANKING order="2" place="2" resultid="50662" />
                    <RANKING order="3" place="3" resultid="48382" />
                    <RANKING order="4" place="-1" resultid="47643" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46445" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46583" />
                    <RANKING order="2" place="2" resultid="50603" />
                    <RANKING order="3" place="3" resultid="47077" />
                    <RANKING order="4" place="4" resultid="46852" />
                    <RANKING order="5" place="5" resultid="50604" />
                    <RANKING order="6" place="6" resultid="46853" />
                    <RANKING order="7" place="7" resultid="49191" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50793" daytime="16:51" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50794" daytime="16:57" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="46291" daytime="17:02" gender="F" number="24" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46446" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="49193" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46447" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48855" />
                    <RANKING order="2" place="2" resultid="48384" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46448" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47003" />
                    <RANKING order="2" place="2" resultid="50607" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46449" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50606" />
                    <RANKING order="2" place="2" resultid="50605" />
                    <RANKING order="3" place="3" resultid="49192" />
                    <RANKING order="4" place="4" resultid="46854" />
                    <RANKING order="5" place="5" resultid="47882" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50795" daytime="17:02" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2021-05-29" daytime="09:00" endtime="12:37" number="3" warmupfrom="07:50" warmupuntil="08:50">
          <EVENTS>
            <EVENT eventid="46294" daytime="09:00" gender="M" number="25" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46396" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47835" />
                    <RANKING order="2" place="2" resultid="46487" />
                    <RANKING order="3" place="3" resultid="50874" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46397" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48094" />
                    <RANKING order="2" place="2" resultid="46481" />
                    <RANKING order="3" place="3" resultid="46652" />
                    <RANKING order="4" place="4" resultid="46779" />
                    <RANKING order="5" place="5" resultid="48059" />
                    <RANKING order="6" place="6" resultid="47623" />
                    <RANKING order="7" place="7" resultid="48840" />
                    <RANKING order="8" place="8" resultid="46632" />
                    <RANKING order="9" place="9" resultid="50340" />
                    <RANKING order="10" place="10" resultid="48497" />
                    <RANKING order="11" place="11" resultid="50333" />
                    <RANKING order="12" place="12" resultid="48253" />
                    <RANKING order="13" place="13" resultid="47102" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46398" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47657" />
                    <RANKING order="2" place="2" resultid="48688" />
                    <RANKING order="3" place="3" resultid="48697" />
                    <RANKING order="4" place="4" resultid="50354" />
                    <RANKING order="5" place="5" resultid="46642" />
                    <RANKING order="6" place="6" resultid="50360" />
                    <RANKING order="7" place="7" resultid="48706" />
                    <RANKING order="8" place="8" resultid="46726" />
                    <RANKING order="9" place="9" resultid="48077" />
                    <RANKING order="10" place="10" resultid="48223" />
                    <RANKING order="11" place="11" resultid="48231" />
                    <RANKING order="12" place="12" resultid="46612" />
                    <RANKING order="13" place="13" resultid="46602" />
                    <RANKING order="14" place="14" resultid="46622" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46399" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46591" />
                    <RANKING order="2" place="2" resultid="48444" />
                    <RANKING order="3" place="3" resultid="50407" />
                    <RANKING order="4" place="4" resultid="47086" />
                    <RANKING order="5" place="5" resultid="47556" />
                    <RANKING order="6" place="6" resultid="50399" />
                    <RANKING order="7" place="7" resultid="47822" />
                    <RANKING order="8" place="8" resultid="47549" />
                    <RANKING order="9" place="9" resultid="48406" />
                    <RANKING order="10" place="10" resultid="49200" />
                    <RANKING order="11" place="11" resultid="49179" />
                    <RANKING order="12" place="12" resultid="47667" />
                    <RANKING order="13" place="13" resultid="46802" />
                    <RANKING order="14" place="14" resultid="48132" />
                    <RANKING order="15" place="-1" resultid="50891" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50796" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50797" daytime="09:07" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50798" daytime="09:13" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50799" daytime="09:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="50800" daytime="09:26" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="46296" daytime="09:31" gender="F" number="26" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46400" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="49144" />
                    <RANKING order="2" place="2" resultid="48332" />
                    <RANKING order="3" place="3" resultid="48835" />
                    <RANKING order="4" place="4" resultid="49165" />
                    <RANKING order="5" place="5" resultid="50530" />
                    <RANKING order="6" place="6" resultid="46712" />
                    <RANKING order="7" place="7" resultid="46548" />
                    <RANKING order="8" place="8" resultid="49137" />
                    <RANKING order="9" place="9" resultid="49109" />
                    <RANKING order="10" place="-1" resultid="46494" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46401" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47845" />
                    <RANKING order="2" place="2" resultid="50439" />
                    <RANKING order="3" place="3" resultid="46786" />
                    <RANKING order="4" place="4" resultid="48434" />
                    <RANKING order="5" place="5" resultid="49130" />
                    <RANKING order="6" place="6" resultid="47955" />
                    <RANKING order="7" place="7" resultid="46692" />
                    <RANKING order="8" place="8" resultid="48290" />
                    <RANKING order="9" place="-1" resultid="49151" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46402" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48461" />
                    <RANKING order="2" place="2" resultid="50576" />
                    <RANKING order="3" place="3" resultid="48429" />
                    <RANKING order="4" place="4" resultid="47679" />
                    <RANKING order="5" place="5" resultid="46742" />
                    <RANKING order="6" place="6" resultid="46702" />
                    <RANKING order="7" place="7" resultid="48282" />
                    <RANKING order="8" place="8" resultid="50421" />
                    <RANKING order="9" place="9" resultid="46682" />
                    <RANKING order="10" place="10" resultid="46662" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46403" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47090" />
                    <RANKING order="2" place="2" resultid="50488" />
                    <RANKING order="3" place="3" resultid="47569" />
                    <RANKING order="4" place="4" resultid="47674" />
                    <RANKING order="5" place="5" resultid="50581" />
                    <RANKING order="6" place="6" resultid="50552" />
                    <RANKING order="7" place="7" resultid="46736" />
                    <RANKING order="8" place="8" resultid="46672" />
                    <RANKING order="9" place="9" resultid="46843" />
                    <RANKING order="10" place="10" resultid="46814" />
                    <RANKING order="11" place="11" resultid="47873" />
                    <RANKING order="12" place="12" resultid="48158" />
                    <RANKING order="13" place="-1" resultid="49158" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50801" daytime="09:31" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50802" daytime="09:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50803" daytime="09:44" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50804" daytime="09:51" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="50805" daytime="09:58" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="46298" daytime="10:04" gender="M" number="27" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46404" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46902" />
                    <RANKING order="2" place="2" resultid="47025" />
                    <RANKING order="3" place="3" resultid="47663" />
                    <RANKING order="4" place="4" resultid="48260" />
                    <RANKING order="5" place="5" resultid="47836" />
                    <RANKING order="6" place="6" resultid="46488" />
                    <RANKING order="7" place="7" resultid="47596" />
                    <RANKING order="8" place="8" resultid="50875" />
                    <RANKING order="9" place="9" resultid="48773" />
                    <RANKING order="10" place="10" resultid="47221" />
                    <RANKING order="11" place="11" resultid="47988" />
                    <RANKING order="12" place="12" resultid="46731" />
                    <RANKING order="13" place="13" resultid="47138" />
                    <RANKING order="14" place="14" resultid="48266" />
                    <RANKING order="15" place="15" resultid="46923" />
                    <RANKING order="16" place="16" resultid="46515" />
                    <RANKING order="17" place="17" resultid="49099" />
                    <RANKING order="18" place="18" resultid="47994" />
                    <RANKING order="19" place="19" resultid="50388" />
                    <RANKING order="20" place="20" resultid="48514" />
                    <RANKING order="21" place="21" resultid="47141" />
                    <RANKING order="22" place="-1" resultid="48735" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46405" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47691" />
                    <RANKING order="2" place="2" resultid="47165" />
                    <RANKING order="3" place="3" resultid="50318" />
                    <RANKING order="4" place="4" resultid="48744" />
                    <RANKING order="5" place="5" resultid="46754" />
                    <RANKING order="6" place="6" resultid="47685" />
                    <RANKING order="7" place="7" resultid="48729" />
                    <RANKING order="8" place="8" resultid="50367" />
                    <RANKING order="9" place="9" resultid="46653" />
                    <RANKING order="10" place="10" resultid="48507" />
                    <RANKING order="11" place="11" resultid="46916" />
                    <RANKING order="12" place="12" resultid="50324" />
                    <RANKING order="13" place="13" resultid="47927" />
                    <RANKING order="14" place="14" resultid="47647" />
                    <RANKING order="15" place="15" resultid="47963" />
                    <RANKING order="16" place="16" resultid="47036" />
                    <RANKING order="17" place="17" resultid="46909" />
                    <RANKING order="18" place="18" resultid="48415" />
                    <RANKING order="19" place="19" resultid="46633" />
                    <RANKING order="20" place="19" resultid="48238" />
                    <RANKING order="21" place="21" resultid="47977" />
                    <RANKING order="22" place="22" resultid="48498" />
                    <RANKING order="23" place="23" resultid="48242" />
                    <RANKING order="24" place="24" resultid="49078" />
                    <RANKING order="25" place="25" resultid="50374" />
                    <RANKING order="26" place="26" resultid="46990" />
                    <RANKING order="27" place="27" resultid="50381" />
                    <RANKING order="28" place="28" resultid="48254" />
                    <RANKING order="29" place="29" resultid="46861" />
                    <RANKING order="30" place="30" resultid="47605" />
                    <RANKING order="31" place="31" resultid="46720" />
                    <RANKING order="32" place="32" resultid="49172" />
                    <RANKING order="33" place="33" resultid="50393" />
                    <RANKING order="34" place="34" resultid="48373" />
                    <RANKING order="35" place="35" resultid="49092" />
                    <RANKING order="36" place="36" resultid="47225" />
                    <RANKING order="37" place="37" resultid="48120" />
                    <RANKING order="38" place="38" resultid="48247" />
                    <RANKING order="39" place="39" resultid="48783" />
                    <RANKING order="40" place="40" resultid="48065" />
                    <RANKING order="41" place="41" resultid="47115" />
                    <RANKING order="42" place="-1" resultid="47103" />
                    <RANKING order="43" place="-1" resultid="48633" />
                    <RANKING order="44" place="-1" resultid="48845" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46406" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46969" />
                    <RANKING order="2" place="2" resultid="47888" />
                    <RANKING order="3" place="3" resultid="47658" />
                    <RANKING order="4" place="4" resultid="48452" />
                    <RANKING order="5" place="5" resultid="46975" />
                    <RANKING order="6" place="6" resultid="48698" />
                    <RANKING order="7" place="7" resultid="46534" />
                    <RANKING order="8" place="8" resultid="48232" />
                    <RANKING order="9" place="9" resultid="48165" />
                    <RANKING order="10" place="10" resultid="50347" />
                    <RANKING order="11" place="11" resultid="48689" />
                    <RANKING order="12" place="12" resultid="46522" />
                    <RANKING order="13" place="13" resultid="46810" />
                    <RANKING order="14" place="14" resultid="49085" />
                    <RANKING order="15" place="15" resultid="48707" />
                    <RANKING order="16" place="15" resultid="50361" />
                    <RANKING order="17" place="17" resultid="46527" />
                    <RANKING order="18" place="18" resultid="47600" />
                    <RANKING order="19" place="19" resultid="47640" />
                    <RANKING order="20" place="20" resultid="46994" />
                    <RANKING order="21" place="21" resultid="48640" />
                    <RANKING order="22" place="22" resultid="46643" />
                    <RANKING order="23" place="23" resultid="46603" />
                    <RANKING order="24" place="24" resultid="46727" />
                    <RANKING order="25" place="25" resultid="48215" />
                    <RANKING order="26" place="26" resultid="46613" />
                    <RANKING order="27" place="27" resultid="46510" />
                    <RANKING order="28" place="28" resultid="48209" />
                    <RANKING order="29" place="29" resultid="48072" />
                    <RANKING order="30" place="30" resultid="46623" />
                    <RANKING order="31" place="-1" resultid="46869" />
                    <RANKING order="32" place="-1" resultid="47153" />
                    <RANKING order="33" place="-1" resultid="47149" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46407" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47168" />
                    <RANKING order="2" place="2" resultid="46557" />
                    <RANKING order="3" place="3" resultid="48680" />
                    <RANKING order="4" place="4" resultid="46463" />
                    <RANKING order="5" place="5" resultid="48757" />
                    <RANKING order="6" place="6" resultid="49641" />
                    <RANKING order="7" place="7" resultid="47563" />
                    <RANKING order="8" place="8" resultid="47082" />
                    <RANKING order="9" place="9" resultid="46592" />
                    <RANKING order="10" place="10" resultid="46554" />
                    <RANKING order="11" place="11" resultid="48177" />
                    <RANKING order="12" place="12" resultid="47075" />
                    <RANKING order="13" place="13" resultid="48402" />
                    <RANKING order="14" place="14" resultid="47031" />
                    <RANKING order="15" place="15" resultid="47071" />
                    <RANKING order="16" place="16" resultid="47550" />
                    <RANKING order="17" place="16" resultid="48202" />
                    <RANKING order="18" place="18" resultid="48628" />
                    <RANKING order="19" place="19" resultid="50595" />
                    <RANKING order="20" place="20" resultid="49649" />
                    <RANKING order="21" place="21" resultid="48140" />
                    <RANKING order="22" place="21" resultid="48751" />
                    <RANKING order="23" place="23" resultid="47145" />
                    <RANKING order="24" place="24" resultid="47061" />
                    <RANKING order="25" place="25" resultid="46561" />
                    <RANKING order="26" place="26" resultid="46566" />
                    <RANKING order="27" place="27" resultid="48472" />
                    <RANKING order="28" place="28" resultid="50558" />
                    <RANKING order="29" place="29" resultid="47899" />
                    <RANKING order="30" place="30" resultid="48102" />
                    <RANKING order="31" place="31" resultid="48761" />
                    <RANKING order="32" place="32" resultid="48714" />
                    <RANKING order="33" place="33" resultid="46838" />
                    <RANKING order="34" place="34" resultid="49897" />
                    <RANKING order="35" place="35" resultid="48647" />
                    <RANKING order="36" place="36" resultid="48410" />
                    <RANKING order="37" place="36" resultid="50564" />
                    <RANKING order="38" place="38" resultid="50500" />
                    <RANKING order="39" place="39" resultid="49103" />
                    <RANKING order="40" place="40" resultid="50506" />
                    <RANKING order="41" place="41" resultid="48393" />
                    <RANKING order="42" place="42" resultid="48397" />
                    <RANKING order="43" place="43" resultid="46797" />
                    <RANKING order="44" place="44" resultid="47161" />
                    <RANKING order="45" place="45" resultid="47982" />
                    <RANKING order="46" place="46" resultid="48049" />
                    <RANKING order="47" place="47" resultid="48171" />
                    <RANKING order="48" place="48" resultid="47010" />
                    <RANKING order="49" place="49" resultid="47650" />
                    <RANKING order="50" place="50" resultid="48052" />
                    <RANKING order="51" place="51" resultid="48589" />
                    <RANKING order="52" place="52" resultid="47894" />
                    <RANKING order="53" place="53" resultid="46571" />
                    <RANKING order="54" place="54" resultid="47189" />
                    <RANKING order="55" place="55" resultid="47970" />
                    <RANKING order="56" place="56" resultid="47016" />
                    <RANKING order="57" place="57" resultid="47109" />
                    <RANKING order="58" place="58" resultid="48012" />
                    <RANKING order="59" place="59" resultid="49072" />
                    <RANKING order="60" place="60" resultid="47587" />
                    <RANKING order="61" place="61" resultid="47233" />
                    <RANKING order="62" place="62" resultid="48116" />
                    <RANKING order="63" place="63" resultid="50910" />
                    <RANKING order="64" place="-1" resultid="47157" />
                    <RANKING order="65" place="-1" resultid="47239" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50806" daytime="10:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50807" daytime="10:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50808" daytime="10:07" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50809" daytime="10:09" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="50810" daytime="10:11" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="50811" daytime="10:13" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="50812" daytime="10:14" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="50813" daytime="10:16" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="50814" daytime="10:18" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="50815" daytime="10:19" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="50816" daytime="10:21" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="50817" daytime="10:22" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="50818" daytime="10:24" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="50819" daytime="10:25" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="50820" daytime="10:27" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="50821" daytime="10:28" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="50822" daytime="10:29" number="17" order="17" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="46300" daytime="10:31" gender="F" number="28" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46408" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="49145" />
                    <RANKING order="2" place="2" resultid="50464" />
                    <RANKING order="3" place="3" resultid="46495" />
                    <RANKING order="4" place="4" resultid="46713" />
                    <RANKING order="5" place="5" resultid="47999" />
                    <RANKING order="6" place="6" resultid="47050" />
                    <RANKING order="7" place="7" resultid="48006" />
                    <RANKING order="8" place="8" resultid="47210" />
                    <RANKING order="9" place="9" resultid="50445" />
                    <RANKING order="10" place="10" resultid="47173" />
                    <RANKING order="11" place="11" resultid="48194" />
                    <RANKING order="12" place="12" resultid="50531" />
                    <RANKING order="13" place="13" resultid="50451" />
                    <RANKING order="14" place="14" resultid="50536" />
                    <RANKING order="15" place="15" resultid="47066" />
                    <RANKING order="16" place="16" resultid="48525" />
                    <RANKING order="17" place="17" resultid="47879" />
                    <RANKING order="18" place="18" resultid="50457" />
                    <RANKING order="19" place="19" resultid="50878" />
                    <RANKING order="20" place="20" resultid="46774" />
                    <RANKING order="21" place="21" resultid="47217" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46409" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46998" />
                    <RANKING order="2" place="2" resultid="50440" />
                    <RANKING order="3" place="3" resultid="47846" />
                    <RANKING order="4" place="4" resultid="48272" />
                    <RANKING order="5" place="5" resultid="50483" />
                    <RANKING order="6" place="6" resultid="48421" />
                    <RANKING order="7" place="7" resultid="47851" />
                    <RANKING order="8" place="8" resultid="48083" />
                    <RANKING order="9" place="9" resultid="49654" />
                    <RANKING order="10" place="10" resultid="48653" />
                    <RANKING order="11" place="11" resultid="48621" />
                    <RANKING order="12" place="12" resultid="47053" />
                    <RANKING order="13" place="13" resultid="48318" />
                    <RANKING order="14" place="14" resultid="48029" />
                    <RANKING order="15" place="15" resultid="48189" />
                    <RANKING order="16" place="16" resultid="46888" />
                    <RANKING order="17" place="17" resultid="47214" />
                    <RANKING order="18" place="18" resultid="48663" />
                    <RANKING order="19" place="19" resultid="46693" />
                    <RANKING order="20" place="19" resultid="48112" />
                    <RANKING order="21" place="21" resultid="48291" />
                    <RANKING order="22" place="22" resultid="48302" />
                    <RANKING order="23" place="23" resultid="48547" />
                    <RANKING order="24" place="24" resultid="48296" />
                    <RANKING order="25" place="25" resultid="48313" />
                    <RANKING order="26" place="26" resultid="48308" />
                    <RANKING order="27" place="-1" resultid="46894" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46410" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46964" />
                    <RANKING order="2" place="2" resultid="47044" />
                    <RANKING order="3" place="3" resultid="48430" />
                    <RANKING order="4" place="4" resultid="46538" />
                    <RANKING order="5" place="4" resultid="50428" />
                    <RANKING order="6" place="6" resultid="47680" />
                    <RANKING order="7" place="7" resultid="50414" />
                    <RANKING order="8" place="8" resultid="48532" />
                    <RANKING order="9" place="9" resultid="46743" />
                    <RANKING order="10" place="10" resultid="47182" />
                    <RANKING order="11" place="11" resultid="46937" />
                    <RANKING order="12" place="12" resultid="48594" />
                    <RANKING order="13" place="13" resultid="48286" />
                    <RANKING order="14" place="14" resultid="46764" />
                    <RANKING order="15" place="15" resultid="47186" />
                    <RANKING order="16" place="16" resultid="46703" />
                    <RANKING order="17" place="17" resultid="47206" />
                    <RANKING order="18" place="18" resultid="48182" />
                    <RANKING order="19" place="19" resultid="47615" />
                    <RANKING order="20" place="20" resultid="48540" />
                    <RANKING order="21" place="21" resultid="48659" />
                    <RANKING order="22" place="22" resultid="46683" />
                    <RANKING order="23" place="23" resultid="46663" />
                    <RANKING order="24" place="-1" resultid="49122" />
                    <RANKING order="25" place="-1" resultid="49660" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46411" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50592" />
                    <RANKING order="2" place="2" resultid="47675" />
                    <RANKING order="3" place="3" resultid="50469" />
                    <RANKING order="4" place="4" resultid="50525" />
                    <RANKING order="5" place="5" resultid="50476" />
                    <RANKING order="6" place="6" resultid="48480" />
                    <RANKING order="7" place="7" resultid="47236" />
                    <RANKING order="8" place="8" resultid="49672" />
                    <RANKING order="9" place="9" resultid="46577" />
                    <RANKING order="10" place="10" resultid="50519" />
                    <RANKING order="11" place="11" resultid="50586" />
                    <RANKING order="12" place="12" resultid="50489" />
                    <RANKING order="13" place="13" resultid="50433" />
                    <RANKING order="14" place="14" resultid="46883" />
                    <RANKING order="15" place="15" resultid="49116" />
                    <RANKING order="16" place="16" resultid="46930" />
                    <RANKING order="17" place="17" resultid="46469" />
                    <RANKING order="18" place="18" resultid="46821" />
                    <RANKING order="19" place="19" resultid="46673" />
                    <RANKING order="20" place="20" resultid="49666" />
                    <RANKING order="21" place="21" resultid="47575" />
                    <RANKING order="22" place="22" resultid="47580" />
                    <RANKING order="23" place="23" resultid="48765" />
                    <RANKING order="24" place="24" resultid="48152" />
                    <RANKING order="25" place="25" resultid="48034" />
                    <RANKING order="26" place="26" resultid="47904" />
                    <RANKING order="27" place="27" resultid="47177" />
                    <RANKING order="28" place="28" resultid="49159" />
                    <RANKING order="29" place="29" resultid="46737" />
                    <RANKING order="30" place="30" resultid="48044" />
                    <RANKING order="31" place="31" resultid="47128" />
                    <RANKING order="32" place="32" resultid="47910" />
                    <RANKING order="33" place="33" resultid="46834" />
                    <RANKING order="34" place="34" resultid="48023" />
                    <RANKING order="35" place="35" resultid="48136" />
                    <RANKING order="36" place="36" resultid="46500" />
                    <RANKING order="37" place="37" resultid="46815" />
                    <RANKING order="38" place="38" resultid="48197" />
                    <RANKING order="39" place="39" resultid="47858" />
                    <RANKING order="40" place="40" resultid="47134" />
                    <RANKING order="41" place="41" resultid="47229" />
                    <RANKING order="42" place="42" resultid="46582" />
                    <RANKING order="43" place="43" resultid="47874" />
                    <RANKING order="44" place="44" resultid="47241" />
                    <RANKING order="45" place="45" resultid="47197" />
                    <RANKING order="46" place="46" resultid="47866" />
                    <RANKING order="47" place="47" resultid="47201" />
                    <RANKING order="48" place="-1" resultid="47122" />
                    <RANKING order="49" place="-1" resultid="47192" />
                    <RANKING order="50" place="-1" resultid="48425" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50823" daytime="10:31" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50824" daytime="10:33" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50825" daytime="10:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50826" daytime="10:36" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="50827" daytime="10:37" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="50828" daytime="10:39" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="50829" daytime="10:41" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="50830" daytime="10:42" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="50831" daytime="10:44" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="50832" daytime="10:45" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="50833" daytime="10:47" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="50834" daytime="10:48" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="50835" daytime="10:50" number="13" order="13" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="46302" daytime="10:51" gender="M" number="29" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46412" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48799" />
                    <RANKING order="2" place="2" resultid="46545" />
                    <RANKING order="3" place="3" resultid="48351" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46413" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47686" />
                    <RANKING order="2" place="2" resultid="48508" />
                    <RANKING order="3" place="3" resultid="46755" />
                    <RANKING order="4" place="4" resultid="47624" />
                    <RANKING order="5" place="5" resultid="50368" />
                    <RANKING order="6" place="6" resultid="47116" />
                    <RANKING order="7" place="7" resultid="48066" />
                    <RANKING order="8" place="8" resultid="46482" />
                    <RANKING order="9" place="9" resultid="48344" />
                    <RANKING order="10" place="10" resultid="48794" />
                    <RANKING order="11" place="11" resultid="49173" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46414" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50495" />
                    <RANKING order="2" place="2" resultid="48690" />
                    <RANKING order="3" place="3" resultid="48233" />
                    <RANKING order="4" place="4" resultid="48216" />
                    <RANKING order="5" place="-1" resultid="47628" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46415" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="49892" />
                    <RANKING order="2" place="2" resultid="46828" />
                    <RANKING order="3" place="3" resultid="50570" />
                    <RANKING order="4" place="4" resultid="50507" />
                    <RANKING order="5" place="5" resultid="48456" />
                    <RANKING order="6" place="6" resultid="46825" />
                    <RANKING order="7" place="7" resultid="47057" />
                    <RANKING order="8" place="8" resultid="50501" />
                    <RANKING order="9" place="9" resultid="49650" />
                    <RANKING order="10" place="10" resultid="49180" />
                    <RANKING order="11" place="11" resultid="50403" />
                    <RANKING order="12" place="12" resultid="49898" />
                    <RANKING order="13" place="13" resultid="47110" />
                    <RANKING order="14" place="-1" resultid="47017" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50836" daytime="10:51" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50837" daytime="10:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50838" daytime="11:01" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50839" daytime="11:06" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="46304" daytime="11:10" gender="F" number="30" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46416" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48326" />
                    <RANKING order="2" place="2" resultid="47946" />
                    <RANKING order="3" place="3" resultid="47951" />
                    <RANKING order="4" place="4" resultid="48368" />
                    <RANKING order="5" place="5" resultid="47880" />
                    <RANKING order="6" place="6" resultid="50452" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46417" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48448" />
                    <RANKING order="2" place="2" resultid="47941" />
                    <RANKING order="3" place="3" resultid="46986" />
                    <RANKING order="4" place="4" resultid="50513" />
                    <RANKING order="5" place="5" resultid="46770" />
                    <RANKING order="6" place="6" resultid="48440" />
                    <RANKING order="7" place="7" resultid="48362" />
                    <RANKING order="8" place="8" resultid="48357" />
                    <RANKING order="9" place="9" resultid="48819" />
                    <RANKING order="10" place="10" resultid="48297" />
                    <RANKING order="11" place="11" resultid="48548" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46418" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47916" />
                    <RANKING order="2" place="2" resultid="48124" />
                    <RANKING order="3" place="3" resultid="46765" />
                    <RANKING order="4" place="4" resultid="46506" />
                    <RANKING order="5" place="5" resultid="49123" />
                    <RANKING order="6" place="-1" resultid="49661" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46419" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47576" />
                    <RANKING order="2" place="2" resultid="46474" />
                    <RANKING order="3" place="3" resultid="46759" />
                    <RANKING order="4" place="4" resultid="47581" />
                    <RANKING order="5" place="5" resultid="48603" />
                    <RANKING order="6" place="6" resultid="47827" />
                    <RANKING order="7" place="7" resultid="48599" />
                    <RANKING order="8" place="8" resultid="47632" />
                    <RANKING order="9" place="-1" resultid="47123" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50840" daytime="11:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50841" daytime="11:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50842" daytime="11:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50843" daytime="11:24" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="46306" daytime="11:28" gender="M" number="31" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46420" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46903" />
                    <RANKING order="2" place="2" resultid="47837" />
                    <RANKING order="3" place="3" resultid="48779" />
                    <RANKING order="4" place="4" resultid="48267" />
                    <RANKING order="5" place="-1" resultid="48515" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46421" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48745" />
                    <RANKING order="2" place="2" resultid="50896" />
                    <RANKING order="3" place="3" resultid="48088" />
                    <RANKING order="4" place="4" resultid="46917" />
                    <RANKING order="5" place="5" resultid="46654" />
                    <RANKING order="6" place="6" resultid="50382" />
                    <RANKING order="7" place="7" resultid="50341" />
                    <RANKING order="8" place="8" resultid="48499" />
                    <RANKING order="9" place="9" resultid="46634" />
                    <RANKING order="10" place="10" resultid="48060" />
                    <RANKING order="11" place="11" resultid="46721" />
                    <RANKING order="12" place="12" resultid="47964" />
                    <RANKING order="13" place="13" resultid="48339" />
                    <RANKING order="14" place="14" resultid="48789" />
                    <RANKING order="15" place="15" resultid="47978" />
                    <RANKING order="16" place="16" resultid="47648" />
                    <RANKING order="17" place="17" resultid="50334" />
                    <RANKING order="18" place="-1" resultid="48634" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46422" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50355" />
                    <RANKING order="2" place="2" resultid="48389" />
                    <RANKING order="3" place="3" resultid="46535" />
                    <RANKING order="4" place="4" resultid="48699" />
                    <RANKING order="5" place="5" resultid="46981" />
                    <RANKING order="6" place="6" resultid="48708" />
                    <RANKING order="7" place="7" resultid="48691" />
                    <RANKING order="8" place="8" resultid="47889" />
                    <RANKING order="9" place="9" resultid="47601" />
                    <RANKING order="10" place="10" resultid="46644" />
                    <RANKING order="11" place="11" resultid="46528" />
                    <RANKING order="12" place="12" resultid="48224" />
                    <RANKING order="13" place="13" resultid="46604" />
                    <RANKING order="14" place="14" resultid="46624" />
                    <RANKING order="15" place="15" resultid="46614" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46423" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48672" />
                    <RANKING order="2" place="2" resultid="49642" />
                    <RANKING order="3" place="3" resultid="46593" />
                    <RANKING order="4" place="4" resultid="50596" />
                    <RANKING order="5" place="5" resultid="47032" />
                    <RANKING order="6" place="6" resultid="46847" />
                    <RANKING order="7" place="7" resultid="50408" />
                    <RANKING order="8" place="8" resultid="47564" />
                    <RANKING order="9" place="9" resultid="50559" />
                    <RANKING order="10" place="10" resultid="48752" />
                    <RANKING order="11" place="11" resultid="50544" />
                    <RANKING order="12" place="12" resultid="48629" />
                    <RANKING order="13" place="13" resultid="46562" />
                    <RANKING order="14" place="14" resultid="47651" />
                    <RANKING order="15" place="15" resultid="47900" />
                    <RANKING order="16" place="16" resultid="48590" />
                    <RANKING order="17" place="17" resultid="48172" />
                    <RANKING order="18" place="18" resultid="47011" />
                    <RANKING order="19" place="19" resultid="47592" />
                    <RANKING order="20" place="20" resultid="50892" />
                    <RANKING order="21" place="-1" resultid="47983" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50844" daytime="11:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50845" daytime="11:31" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50846" daytime="11:33" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50847" daytime="11:36" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="50848" daytime="11:38" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="50849" daytime="11:40" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="46308" daytime="11:42" gender="F" number="32" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46424" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50547" />
                    <RANKING order="2" place="2" resultid="48007" />
                    <RANKING order="3" place="3" resultid="48333" />
                    <RANKING order="4" place="4" resultid="49166" />
                    <RANKING order="5" place="5" resultid="48369" />
                    <RANKING order="6" place="6" resultid="46549" />
                    <RANKING order="7" place="7" resultid="46714" />
                    <RANKING order="8" place="8" resultid="48000" />
                    <RANKING order="9" place="9" resultid="48526" />
                    <RANKING order="10" place="-1" resultid="49138" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46425" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46959" />
                    <RANKING order="2" place="2" resultid="48831" />
                    <RANKING order="3" place="3" resultid="47935" />
                    <RANKING order="4" place="4" resultid="46787" />
                    <RANKING order="5" place="5" resultid="48273" />
                    <RANKING order="6" place="6" resultid="48654" />
                    <RANKING order="7" place="7" resultid="48108" />
                    <RANKING order="8" place="8" resultid="48851" />
                    <RANKING order="9" place="9" resultid="50514" />
                    <RANKING order="10" place="10" resultid="48488" />
                    <RANKING order="11" place="11" resultid="46791" />
                    <RANKING order="12" place="12" resultid="47852" />
                    <RANKING order="13" place="13" resultid="48303" />
                    <RANKING order="14" place="14" resultid="46694" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46426" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46965" />
                    <RANKING order="2" place="2" resultid="50577" />
                    <RANKING order="3" place="3" resultid="50415" />
                    <RANKING order="4" place="4" resultid="48595" />
                    <RANKING order="5" place="5" resultid="48541" />
                    <RANKING order="6" place="6" resultid="50422" />
                    <RANKING order="7" place="7" resultid="48533" />
                    <RANKING order="8" place="8" resultid="48183" />
                    <RANKING order="9" place="9" resultid="46704" />
                    <RANKING order="10" place="10" resultid="46684" />
                    <RANKING order="11" place="11" resultid="46664" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46427" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50882" />
                    <RANKING order="2" place="2" resultid="49673" />
                    <RANKING order="3" place="3" resultid="46578" />
                    <RANKING order="4" place="4" resultid="49667" />
                    <RANKING order="5" place="5" resultid="47905" />
                    <RANKING order="6" place="6" resultid="50553" />
                    <RANKING order="7" place="7" resultid="50477" />
                    <RANKING order="8" place="8" resultid="47570" />
                    <RANKING order="9" place="9" resultid="47921" />
                    <RANKING order="10" place="10" resultid="46674" />
                    <RANKING order="11" place="11" resultid="47129" />
                    <RANKING order="12" place="12" resultid="47859" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50897" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50898" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50899" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50900" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="50901" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="46310" daytime="11:55" gender="M" number="33" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46428" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47026" />
                    <RANKING order="2" place="2" resultid="48261" />
                    <RANKING order="3" place="3" resultid="50876" />
                    <RANKING order="4" place="4" resultid="46924" />
                    <RANKING order="5" place="5" resultid="47989" />
                    <RANKING order="6" place="6" resultid="46516" />
                    <RANKING order="7" place="7" resultid="46489" />
                    <RANKING order="8" place="8" resultid="48352" />
                    <RANKING order="9" place="9" resultid="48774" />
                    <RANKING order="10" place="10" resultid="49100" />
                    <RANKING order="11" place="11" resultid="48516" />
                    <RANKING order="12" place="12" resultid="47995" />
                    <RANKING order="13" place="-1" resultid="48148" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46429" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47692" />
                    <RANKING order="2" place="2" resultid="48095" />
                    <RANKING order="3" place="3" resultid="46910" />
                    <RANKING order="4" place="4" resultid="48730" />
                    <RANKING order="5" place="5" resultid="48144" />
                    <RANKING order="6" place="6" resultid="50319" />
                    <RANKING order="7" place="7" resultid="48465" />
                    <RANKING order="8" place="8" resultid="48374" />
                    <RANKING order="9" place="9" resultid="48841" />
                    <RANKING order="10" place="10" resultid="50375" />
                    <RANKING order="11" place="11" resultid="48089" />
                    <RANKING order="12" place="12" resultid="48500" />
                    <RANKING order="13" place="13" resultid="46862" />
                    <RANKING order="14" place="14" resultid="48740" />
                    <RANKING order="15" place="15" resultid="49093" />
                    <RANKING order="16" place="16" resultid="48345" />
                    <RANKING order="17" place="17" resultid="48509" />
                    <RANKING order="18" place="18" resultid="48416" />
                    <RANKING order="19" place="19" resultid="49079" />
                    <RANKING order="20" place="20" resultid="48243" />
                    <RANKING order="21" place="21" resultid="50394" />
                    <RANKING order="22" place="22" resultid="47037" />
                    <RANKING order="23" place="23" resultid="48248" />
                    <RANKING order="24" place="24" resultid="48784" />
                    <RANKING order="25" place="25" resultid="47117" />
                    <RANKING order="26" place="-1" resultid="48846" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46430" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46970" />
                    <RANKING order="2" place="2" resultid="46976" />
                    <RANKING order="3" place="3" resultid="50348" />
                    <RANKING order="4" place="4" resultid="47890" />
                    <RANKING order="5" place="5" resultid="48166" />
                    <RANKING order="6" place="6" resultid="48709" />
                    <RANKING order="7" place="7" resultid="48641" />
                    <RANKING order="8" place="8" resultid="48225" />
                    <RANKING order="9" place="9" resultid="49086" />
                    <RANKING order="10" place="10" resultid="46995" />
                    <RANKING order="11" place="11" resultid="47641" />
                    <RANKING order="12" place="12" resultid="50496" />
                    <RANKING order="13" place="13" resultid="46511" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46431" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48468" />
                    <RANKING order="2" place="2" resultid="47097" />
                    <RANKING order="3" place="3" resultid="47557" />
                    <RANKING order="4" place="4" resultid="48673" />
                    <RANKING order="5" place="5" resultid="46848" />
                    <RANKING order="6" place="6" resultid="48715" />
                    <RANKING order="7" place="7" resultid="46839" />
                    <RANKING order="8" place="8" resultid="48473" />
                    <RANKING order="9" place="9" resultid="48178" />
                    <RANKING order="10" place="10" resultid="47072" />
                    <RANKING order="11" place="11" resultid="47636" />
                    <RANKING order="12" place="12" resultid="50565" />
                    <RANKING order="13" place="13" resultid="46798" />
                    <RANKING order="14" place="14" resultid="48411" />
                    <RANKING order="15" place="15" resultid="47062" />
                    <RANKING order="16" place="16" resultid="48053" />
                    <RANKING order="17" place="17" resultid="47895" />
                    <RANKING order="18" place="18" resultid="48648" />
                    <RANKING order="19" place="19" resultid="46572" />
                    <RANKING order="20" place="-1" resultid="48725" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50855" daytime="11:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50856" daytime="11:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50857" daytime="11:58" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50858" daytime="12:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="50859" daytime="12:02" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="50860" daytime="12:04" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="50861" daytime="12:05" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="50862" daytime="12:07" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="46312" daytime="12:08" gender="F" number="34" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46432" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50465" />
                    <RANKING order="2" place="2" resultid="46496" />
                    <RANKING order="3" place="3" resultid="48836" />
                    <RANKING order="4" place="4" resultid="50446" />
                    <RANKING order="5" place="5" resultid="48008" />
                    <RANKING order="6" place="6" resultid="47067" />
                    <RANKING order="7" place="7" resultid="50458" />
                    <RANKING order="8" place="8" resultid="48527" />
                    <RANKING order="9" place="9" resultid="50537" />
                    <RANKING order="10" place="10" resultid="49110" />
                    <RANKING order="11" place="11" resultid="50880" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46433" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46999" />
                    <RANKING order="2" place="2" resultid="49131" />
                    <RANKING order="3" place="3" resultid="47936" />
                    <RANKING order="4" place="4" resultid="48655" />
                    <RANKING order="5" place="5" resultid="46792" />
                    <RANKING order="6" place="6" resultid="47956" />
                    <RANKING order="7" place="7" resultid="49655" />
                    <RANKING order="8" place="8" resultid="48622" />
                    <RANKING order="9" place="9" resultid="48484" />
                    <RANKING order="10" place="10" resultid="47853" />
                    <RANKING order="11" place="11" resultid="48319" />
                    <RANKING order="12" place="12" resultid="48378" />
                    <RANKING order="13" place="13" resultid="48278" />
                    <RANKING order="14" place="14" resultid="48030" />
                    <RANKING order="15" place="15" resultid="48814" />
                    <RANKING order="16" place="16" resultid="48190" />
                    <RANKING order="17" place="17" resultid="46889" />
                    <RANKING order="18" place="18" resultid="48363" />
                    <RANKING order="19" place="-1" resultid="46895" />
                    <RANKING order="20" place="-1" resultid="48549" />
                    <RANKING order="21" place="-1" resultid="48804" />
                    <RANKING order="22" place="-1" resultid="49152" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46434" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="47045" />
                    <RANKING order="2" place="2" resultid="46539" />
                    <RANKING order="3" place="3" resultid="47681" />
                    <RANKING order="4" place="4" resultid="50429" />
                    <RANKING order="5" place="5" resultid="48476" />
                    <RANKING order="6" place="6" resultid="46938" />
                    <RANKING order="7" place="7" resultid="48542" />
                    <RANKING order="8" place="8" resultid="48667" />
                    <RANKING order="9" place="9" resultid="49124" />
                    <RANKING order="10" place="-1" resultid="48534" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46435" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50883" />
                    <RANKING order="2" place="2" resultid="49678" />
                    <RANKING order="3" place="3" resultid="48481" />
                    <RANKING order="4" place="4" resultid="50470" />
                    <RANKING order="5" place="5" resultid="49674" />
                    <RANKING order="6" place="6" resultid="50520" />
                    <RANKING order="7" place="7" resultid="50582" />
                    <RANKING order="8" place="8" resultid="50587" />
                    <RANKING order="9" place="9" resultid="49117" />
                    <RANKING order="10" place="10" resultid="46931" />
                    <RANKING order="11" place="11" resultid="47237" />
                    <RANKING order="12" place="12" resultid="48153" />
                    <RANKING order="13" place="13" resultid="47178" />
                    <RANKING order="14" place="14" resultid="48035" />
                    <RANKING order="15" place="15" resultid="48045" />
                    <RANKING order="16" place="16" resultid="48607" />
                    <RANKING order="17" place="17" resultid="47911" />
                    <RANKING order="18" place="18" resultid="48025" />
                    <RANKING order="19" place="19" resultid="48159" />
                    <RANKING order="20" place="20" resultid="46501" />
                    <RANKING order="21" place="21" resultid="48198" />
                    <RANKING order="22" place="22" resultid="47230" />
                    <RANKING order="23" place="23" resultid="47860" />
                    <RANKING order="24" place="24" resultid="47867" />
                    <RANKING order="25" place="25" resultid="47242" />
                    <RANKING order="26" place="26" resultid="47202" />
                    <RANKING order="27" place="-1" resultid="47193" />
                    <RANKING order="28" place="-1" resultid="48128" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50902" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="50903" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="50904" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="50905" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="50906" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="50907" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="50908" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="50909" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="46314" daytime="12:20" gender="M" number="35" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46450" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="46451" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="46953" />
                    <RANKING order="2" place="2" resultid="48856" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46452" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="46453" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50608" />
                    <RANKING order="2" place="2" resultid="47644" />
                    <RANKING order="3" place="3" resultid="49194" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50870" daytime="12:20" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="46316" daytime="12:31" gender="F" number="36" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="46454" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="49196" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46455" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="48857" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="46456" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="46457" agemax="95" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="50609" />
                    <RANKING order="2" place="2" resultid="49195" />
                    <RANKING order="3" place="3" resultid="47883" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="50871" daytime="12:31" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="00701" nation="POL" region="01" clubid="47135" name="MKS Dziewiątka Dzierżoniów">
          <ATHLETES>
            <ATHLETE firstname="Mateusz" lastname="Kut" birthdate="2004-10-03" gender="M" nation="POL" license="100701700088" swrid="5287590" athleteid="47154">
              <RESULTS>
                <RESULT eventid="44378" status="DNS" swimtime="00:00:00.00" resultid="47155" heatid="50664" lane="0" />
                <RESULT eventid="44411" status="DNS" swimtime="00:00:00.00" resultid="47156" heatid="50762" lane="2" entrytime="00:00:38.48" entrycourse="LCM" />
                <RESULT eventid="46298" status="DNS" swimtime="00:00:00.00" resultid="47157" heatid="50814" lane="9" entrytime="00:00:32.86" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominik" lastname="Pietrewicz" birthdate="2003-10-13" gender="M" nation="POL" license="100701700071" swrid="4012815" athleteid="47187">
              <RESULTS>
                <RESULT eventid="44382" points="314" reactiontime="+67" swimtime="00:00:38.14" resultid="47188" heatid="50693" lane="6" entrytime="00:00:38.50" entrycourse="LCM" />
                <RESULT eventid="46298" points="422" reactiontime="+64" swimtime="00:00:27.87" resultid="47189" heatid="50817" lane="2" entrytime="00:00:28.16" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lateef" lastname="Hanus" birthdate="2005-06-29" gender="M" nation="POL" license="100701700087" swrid="5143702" athleteid="47231">
              <RESULTS>
                <RESULT eventid="44411" points="277" reactiontime="+71" swimtime="00:00:34.14" resultid="47232" heatid="50758" lane="7" />
                <RESULT eventid="46298" points="366" reactiontime="+75" swimtime="00:00:29.22" resultid="47233" heatid="50813" lane="8" entrytime="00:00:33.58" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Gutkowska" birthdate="2007-06-12" gender="F" nation="POL" license="100701600132" swrid="5094202" athleteid="47211">
              <RESULTS>
                <RESULT eventid="44384" points="313" reactiontime="+71" swimtime="00:00:43.26" resultid="47212" heatid="50698" lane="3" />
                <RESULT eventid="44413" points="330" swimtime="00:00:35.32" resultid="47213" heatid="50771" lane="4" />
                <RESULT eventid="46300" points="362" reactiontime="+64" swimtime="00:00:33.20" resultid="47214" heatid="50827" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Magdalena" lastname="Ramilowska" birthdate="2006-04-19" gender="F" nation="POL" license="100701600078" swrid="4995335" athleteid="47183">
              <RESULTS>
                <RESULT eventid="44380" points="397" reactiontime="+68" swimtime="00:01:10.30" resultid="47184" heatid="50679" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="342" reactiontime="+49" swimtime="00:00:34.90" resultid="47185" heatid="50774" lane="4" entrytime="00:00:37.98" entrycourse="LCM" />
                <RESULT eventid="46300" points="427" reactiontime="+69" swimtime="00:00:31.42" resultid="47186" heatid="50826" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Raszewska" birthdate="2008-03-01" gender="F" nation="POL" license="100701600127" swrid="5165952" athleteid="47169">
              <RESULTS>
                <RESULT eventid="44380" points="393" reactiontime="+70" swimtime="00:01:10.59" resultid="47170" heatid="50678" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44384" points="322" reactiontime="+53" swimtime="00:00:42.89" resultid="47171" heatid="50698" lane="4" />
                <RESULT eventid="44413" points="280" reactiontime="+75" swimtime="00:00:37.31" resultid="47172" heatid="50772" lane="8" />
                <RESULT eventid="46300" points="395" reactiontime="+72" swimtime="00:00:32.24" resultid="47173" heatid="50824" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hanna" lastname="Nawrot" birthdate="2006-05-23" gender="F" nation="POL" license="100701600080" swrid="4995338" athleteid="47179">
              <RESULTS>
                <RESULT eventid="44380" points="465" reactiontime="+68" swimtime="00:01:06.73" resultid="47180" heatid="50679" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="424" reactiontime="+69" swimtime="00:00:32.50" resultid="47181" heatid="50775" lane="1" entrytime="00:00:37.48" entrycourse="LCM" />
                <RESULT eventid="46300" points="502" reactiontime="+64" swimtime="00:00:29.78" resultid="47182" heatid="50830" lane="0" entrytime="00:00:32.46" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Grondkowska" birthdate="2006-01-05" gender="F" nation="POL" license="100701600126" swrid="5112206" athleteid="47203">
              <RESULTS>
                <RESULT eventid="44384" points="408" reactiontime="+94" swimtime="00:00:39.62" resultid="47204" heatid="50699" lane="9" />
                <RESULT eventid="44409" points="355" swimtime="00:01:30.55" resultid="47205" heatid="50751" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="420" reactiontime="+71" swimtime="00:00:31.59" resultid="47206" heatid="50824" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hubert" lastname="Falkowski" birthdate="2008-06-23" gender="M" nation="POL" license="100701700104" swrid="5009407" athleteid="47139">
              <RESULTS>
                <RESULT eventid="44378" points="160" reactiontime="+86" swimtime="00:01:26.39" resultid="47140" heatid="50663" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="194" reactiontime="+79" swimtime="00:00:36.11" resultid="47141" heatid="50808" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Pietrewicz" birthdate="2008-06-22" gender="M" nation="POL" license="100701700096" swrid="5441183" athleteid="47218">
              <RESULTS>
                <RESULT eventid="44394" points="272" reactiontime="+66" swimtime="00:01:19.99" resultid="47219" heatid="50718" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="267" reactiontime="+79" swimtime="00:00:34.57" resultid="47220" heatid="50757" lane="2" />
                <RESULT eventid="46298" points="290" reactiontime="+82" swimtime="00:00:31.56" resultid="47221" heatid="50812" lane="3" entrytime="00:00:35.81" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miłosz" lastname="Sztachelek" birthdate="2005-02-27" gender="M" nation="POL" license="100701700077" swrid="5186702" athleteid="47158">
              <RESULTS>
                <RESULT eventid="44378" points="448" reactiontime="+78" swimtime="00:01:01.29" resultid="47159" heatid="50664" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="399" reactiontime="+66" swimtime="00:00:30.25" resultid="47160" heatid="50764" lane="9" entrytime="00:00:32.87" entrycourse="LCM" />
                <RESULT eventid="46298" points="474" reactiontime="+65" swimtime="00:00:26.81" resultid="47161" heatid="50815" lane="3" entrytime="00:00:29.90" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gaja" lastname="Kopera" birthdate="2008-12-16" gender="F" nation="POL" license="100701600129" swrid="5157137" athleteid="47207">
              <RESULTS>
                <RESULT eventid="44384" points="430" reactiontime="+67" swimtime="00:00:38.95" resultid="47208" heatid="50697" lane="2" />
                <RESULT eventid="44396" points="292" reactiontime="+67" swimtime="00:01:26.76" resultid="47209" heatid="50724" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="402" reactiontime="+79" swimtime="00:00:32.05" resultid="47210" heatid="50826" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Kędzierski" birthdate="2006-06-16" gender="M" nation="POL" license="100701700086" swrid="5395492" athleteid="47150">
              <RESULTS>
                <RESULT eventid="44378" points="328" reactiontime="+54" swimtime="00:01:07.99" resultid="47151" heatid="50663" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="302" reactiontime="+57" swimtime="00:00:33.16" resultid="47152" heatid="50762" lane="7" entrytime="00:00:39.59" entrycourse="LCM" />
                <RESULT comment="O-1" eventid="46298" reactiontime="+49" status="DSQ" swimtime="00:00:00.00" resultid="47153" heatid="50814" lane="2" entrytime="00:00:32.01" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Juraszek" birthdate="1994-10-08" gender="M" nation="POL" license="100701700068" swrid="4114468" athleteid="47166">
              <RESULTS>
                <RESULT eventid="44378" points="825" reactiontime="+63" swimtime="00:00:50.01" resultid="47167" heatid="50677" lane="4" entrytime="00:00:49.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="851" reactiontime="+68" swimtime="00:00:22.06" resultid="47168" heatid="50822" lane="4" entrytime="00:00:21.45" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Tatarzyn" birthdate="2007-06-20" gender="M" nation="POL" license="100701700100" swrid="5088583" athleteid="47222">
              <RESULTS>
                <RESULT eventid="44394" points="224" reactiontime="+52" swimtime="00:01:25.36" resultid="47223" heatid="50719" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="222" reactiontime="+66" swimtime="00:00:36.77" resultid="47224" heatid="50761" lane="4" />
                <RESULT eventid="46298" points="296" reactiontime="+73" swimtime="00:00:31.35" resultid="47225" heatid="50809" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krystian" lastname="Bełtowski" birthdate="2001-02-06" gender="M" nation="POL" license="100701700057" swrid="4711914" athleteid="47142">
              <RESULTS>
                <RESULT eventid="44378" points="584" reactiontime="+67" swimtime="00:00:56.10" resultid="47143" heatid="50675" lane="7" entrytime="00:00:57.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="547" reactiontime="+65" swimtime="00:00:27.22" resultid="47144" heatid="50766" lane="7" entrytime="00:00:29.61" entrycourse="LCM" />
                <RESULT eventid="46298" points="540" reactiontime="+63" swimtime="00:00:25.67" resultid="47145" heatid="50821" lane="8" entrytime="00:00:25.75" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edyta" lastname="Bejster" birthdate="1981-05-21" gender="F" nation="POL" license="100701600124" athleteid="47198">
              <RESULTS>
                <RESULT eventid="44384" points="226" reactiontime="+83" swimtime="00:00:48.23" resultid="47199" heatid="50698" lane="0" />
                <RESULT eventid="44413" points="153" reactiontime="+79" swimtime="00:00:45.64" resultid="47200" heatid="50772" lane="9" />
                <RESULT eventid="46300" points="230" reactiontime="+75" swimtime="00:00:38.59" resultid="47201" heatid="50825" lane="0" />
                <RESULT eventid="46312" points="146" reactiontime="+65" swimtime="00:00:51.21" resultid="47202" heatid="50905" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Wierzbicki" birthdate="2007-01-03" gender="M" nation="POL" license="100701700085" swrid="4995342" athleteid="47162">
              <RESULTS>
                <RESULT eventid="44378" points="498" reactiontime="+79" swimtime="00:00:59.15" resultid="47163" heatid="50664" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="433" reactiontime="+76" swimtime="00:00:29.42" resultid="47164" heatid="50764" lane="2" entrytime="00:00:32.41" entrycourse="LCM" />
                <RESULT eventid="46298" points="496" reactiontime="+75" swimtime="00:00:26.41" resultid="47165" heatid="50818" lane="9" entrytime="00:00:27.66" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Bejster" birthdate="2005-02-28" gender="F" nation="POL" license="100701600082" swrid="5088555" athleteid="47190">
              <RESULTS>
                <RESULT eventid="44384" points="307" reactiontime="+65" swimtime="00:00:43.54" resultid="47191" heatid="50696" lane="3" />
                <RESULT eventid="46300" status="DNS" swimtime="00:00:00.00" resultid="47192" heatid="50832" lane="1" entrytime="00:00:29.94" entrycourse="LCM" />
                <RESULT eventid="46312" status="DNS" swimtime="00:00:00.00" resultid="47193" heatid="50908" lane="8" entrytime="00:00:35.20" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Kwaśny" birthdate="1984-04-02" gender="M" nation="POL" license="100701700117" athleteid="47238">
              <RESULTS>
                <RESULT eventid="46298" status="DNS" swimtime="00:00:00.00" resultid="47239" heatid="50807" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alicja" lastname="Kaucka" birthdate="1988-09-22" gender="F" nation="POL" license="100701600118" athleteid="47240">
              <RESULTS>
                <RESULT eventid="46300" points="322" reactiontime="+79" swimtime="00:00:34.53" resultid="47241" heatid="50827" lane="3" />
                <RESULT eventid="46312" points="224" reactiontime="+75" swimtime="00:00:44.36" resultid="47242" heatid="50903" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patryk" lastname="Falkowski" birthdate="2008-06-23" gender="M" nation="POL" license="100701700105" swrid="5049932" athleteid="47136">
              <RESULTS>
                <RESULT eventid="44378" points="233" reactiontime="+88" swimtime="00:01:16.21" resultid="47137" heatid="50664" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="281" reactiontime="+83" swimtime="00:00:31.90" resultid="47138" heatid="50807" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulina" lastname="Porębska" birthdate="2003-05-09" gender="F" nation="POL" license="100701600075" swrid="4012816" athleteid="47174">
              <RESULTS>
                <RESULT eventid="44380" points="535" reactiontime="+66" swimtime="00:01:03.67" resultid="47175" heatid="50685" lane="4" entrytime="00:01:04.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="479" reactiontime="+76" swimtime="00:00:31.21" resultid="47176" heatid="50778" lane="0" entrytime="00:00:32.10" entrycourse="LCM" />
                <RESULT eventid="46300" points="522" reactiontime="+70" swimtime="00:00:29.39" resultid="47177" heatid="50832" lane="9" entrytime="00:00:30.03" entrycourse="LCM" />
                <RESULT eventid="46312" points="523" reactiontime="+67" swimtime="00:00:33.48" resultid="47178" heatid="50902" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Kwiatkowska" birthdate="2008-10-09" gender="F" nation="POL" license="100701600133" athleteid="47215">
              <RESULTS>
                <RESULT eventid="44384" points="171" reactiontime="+69" swimtime="00:00:52.89" resultid="47216" heatid="50698" lane="6" />
                <RESULT eventid="46300" points="223" reactiontime="+62" swimtime="00:00:39.01" resultid="47217" heatid="50826" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Pisarska" birthdate="1981-11-06" gender="F" nation="POL" license="100701600113" athleteid="47234">
              <RESULTS>
                <RESULT eventid="44413" points="562" reactiontime="+64" swimtime="00:00:29.60" resultid="47235" heatid="50772" lane="1" />
                <RESULT eventid="46300" points="609" reactiontime="+63" swimtime="00:00:27.92" resultid="47236" heatid="50826" lane="8" />
                <RESULT eventid="46312" points="563" reactiontime="+60" swimtime="00:00:32.67" resultid="47237" heatid="50904" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Kwinta" birthdate="2006-11-07" gender="M" nation="POL" license="100701700102" swrid="4995339" athleteid="47146">
              <RESULTS>
                <RESULT eventid="44378" status="DNS" swimtime="00:00:00.00" resultid="47147" heatid="50664" lane="8" />
                <RESULT eventid="44411" status="DNS" swimtime="00:00:00.00" resultid="47148" heatid="50759" lane="0" />
                <RESULT eventid="46298" status="DNS" swimtime="00:00:00.00" resultid="47149" heatid="50811" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Babicka" birthdate="1986-11-23" gender="F" nation="POL" license="100701600122" athleteid="47194">
              <RESULTS>
                <RESULT eventid="44384" points="247" reactiontime="+62" swimtime="00:00:46.83" resultid="47195" heatid="50696" lane="5" />
                <RESULT eventid="44413" points="221" reactiontime="+73" swimtime="00:00:40.36" resultid="47196" heatid="50770" lane="7" />
                <RESULT eventid="46300" points="320" reactiontime="+66" swimtime="00:00:34.59" resultid="47197" heatid="50826" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Wojnowska" birthdate="2005-05-21" gender="F" nation="POL" license="100701600083" swrid="5088568" athleteid="47226">
              <RESULTS>
                <RESULT eventid="44396" points="359" reactiontime="+61" swimtime="00:01:20.95" resultid="47227" heatid="50725" lane="7" entrytime="00:01:25.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44417" points="336" reactiontime="+62" swimtime="00:02:57.30" resultid="47228" heatid="50787" lane="5" entrytime="00:03:14.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.51" />
                    <SPLIT distance="100" swimtime="00:01:26.28" />
                    <SPLIT distance="150" swimtime="00:02:12.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="358" reactiontime="+59" swimtime="00:00:33.32" resultid="47229" heatid="50828" lane="4" entrytime="00:00:35.12" entrycourse="LCM" />
                <RESULT eventid="46312" points="353" reactiontime="+64" swimtime="00:00:38.14" resultid="47230" heatid="50906" lane="7" entrytime="00:00:40.07" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="05801" nation="POL" region="01" clubid="47828" name="UKS &quot;Krośnicka Przystań&quot;">
          <ATHLETES>
            <ATHLETE firstname="Kinga" lastname="Filipiak" birthdate="2005-12-07" gender="F" nation="POL" license="105801600017" swrid="5249608" athleteid="47861">
              <RESULTS>
                <RESULT eventid="44380" points="277" reactiontime="+70" swimtime="00:01:19.29" resultid="47862" heatid="50681" lane="9" entrytime="00:01:17.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44384" points="220" reactiontime="+76" swimtime="00:00:48.66" resultid="47863" heatid="50700" lane="9" entrytime="00:00:46.28" entrycourse="LCM" />
                <RESULT eventid="44409" points="218" reactiontime="+73" swimtime="00:01:46.44" resultid="47864" heatid="50753" lane="0" entrytime="00:01:41.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="219" reactiontime="+88" swimtime="00:00:40.50" resultid="47865" heatid="50774" lane="1" entrytime="00:00:39.90" entrycourse="LCM" />
                <RESULT eventid="46300" points="295" reactiontime="+74" swimtime="00:00:35.52" resultid="47866" heatid="50828" lane="6" entrytime="00:00:35.94" entrycourse="LCM" />
                <RESULT eventid="46312" points="286" reactiontime="+63" swimtime="00:00:40.91" resultid="47867" heatid="50905" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Kułakowska" birthdate="2008-12-19" gender="F" nation="POL" license="105801600030" swrid="5398288" athleteid="47875">
              <RESULTS>
                <RESULT eventid="44380" points="271" reactiontime="+57" swimtime="00:01:19.87" resultid="47876" heatid="50680" lane="1" entrytime="00:01:21.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44384" points="273" reactiontime="+62" swimtime="00:00:45.32" resultid="47877" heatid="50699" lane="5" entrytime="00:00:49.76" entrycourse="LCM" />
                <RESULT eventid="44409" points="282" swimtime="00:01:37.77" resultid="47878" heatid="50752" lane="4" entrytime="00:01:45.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="295" reactiontime="+70" swimtime="00:00:35.53" resultid="47879" heatid="50828" lane="3" entrytime="00:00:35.21" entrycourse="LCM" />
                <RESULT eventid="46304" points="299" reactiontime="+58" swimtime="00:03:27.98" resultid="47880" heatid="50842" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.95" />
                    <SPLIT distance="100" swimtime="00:01:40.54" />
                    <SPLIT distance="150" swimtime="00:02:34.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Bocheńska" birthdate="2005-03-27" gender="F" nation="POL" license="105801600018" swrid="5249552" athleteid="47868">
              <RESULTS>
                <RESULT eventid="44380" points="343" reactiontime="+76" swimtime="00:01:13.82" resultid="47869" heatid="50681" lane="8" entrytime="00:01:16.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="333" reactiontime="+76" swimtime="00:02:42.92" resultid="47870" heatid="50740" lane="3" entrytime="00:02:40.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                    <SPLIT distance="100" swimtime="00:01:19.20" />
                    <SPLIT distance="150" swimtime="00:02:03.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="217" reactiontime="+73" swimtime="00:00:40.65" resultid="47871" heatid="50773" lane="5" entrytime="00:00:44.13" entrycourse="LCM" />
                <RESULT eventid="46287" points="314" reactiontime="+78" swimtime="00:11:53.01" resultid="47872" heatid="50791" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                    <SPLIT distance="100" swimtime="00:01:19.12" />
                    <SPLIT distance="150" swimtime="00:02:04.74" />
                    <SPLIT distance="200" swimtime="00:02:50.09" />
                    <SPLIT distance="250" swimtime="00:03:35.60" />
                    <SPLIT distance="300" swimtime="00:04:21.09" />
                    <SPLIT distance="350" swimtime="00:05:07.13" />
                    <SPLIT distance="400" swimtime="00:05:52.20" />
                    <SPLIT distance="450" swimtime="00:06:38.03" />
                    <SPLIT distance="500" swimtime="00:07:24.32" />
                    <SPLIT distance="550" swimtime="00:08:10.22" />
                    <SPLIT distance="600" swimtime="00:08:55.90" />
                    <SPLIT distance="650" swimtime="00:09:41.12" />
                    <SPLIT distance="700" swimtime="00:10:26.81" />
                    <SPLIT distance="750" swimtime="00:11:11.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="319" reactiontime="+80" swimtime="00:05:45.99" resultid="47873" heatid="50804" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.78" />
                    <SPLIT distance="100" swimtime="00:01:18.29" />
                    <SPLIT distance="150" swimtime="00:02:02.90" />
                    <SPLIT distance="200" swimtime="00:02:47.40" />
                    <SPLIT distance="250" swimtime="00:03:32.73" />
                    <SPLIT distance="300" swimtime="00:04:18.87" />
                    <SPLIT distance="350" swimtime="00:05:04.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="332" reactiontime="+77" swimtime="00:00:34.18" resultid="47874" heatid="50828" lane="2" entrytime="00:00:37.36" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patrycja" lastname="Giewiada" birthdate="2007-06-20" gender="F" nation="POL" license="105801600014" swrid="5214751" athleteid="47838">
              <RESULTS>
                <RESULT eventid="44380" points="583" reactiontime="+75" swimtime="00:01:01.88" resultid="47839" heatid="50688" lane="8" entrytime="00:01:01.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44384" points="531" reactiontime="+78" swimtime="00:00:36.30" resultid="47840" heatid="50701" lane="1" entrytime="00:00:42.29" entrycourse="LCM" />
                <RESULT eventid="44392" points="548" reactiontime="+75" swimtime="00:02:34.05" resultid="47841" heatid="50716" lane="8" entrytime="00:02:33.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                    <SPLIT distance="100" swimtime="00:01:15.26" />
                    <SPLIT distance="150" swimtime="00:01:59.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="581" reactiontime="+69" swimtime="00:02:15.36" resultid="47842" heatid="50744" lane="0" entrytime="00:02:15.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.31" />
                    <SPLIT distance="100" swimtime="00:01:05.60" />
                    <SPLIT distance="150" swimtime="00:01:40.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44409" status="DNS" swimtime="00:00:00.00" resultid="47843" heatid="50755" lane="3" entrytime="00:01:19.06" entrycourse="LCM" />
                <RESULT eventid="44413" points="435" reactiontime="+75" swimtime="00:00:32.22" resultid="47844" heatid="50777" lane="3" entrytime="00:00:32.75" entrycourse="LCM" />
                <RESULT eventid="46296" points="545" reactiontime="+73" swimtime="00:04:49.47" resultid="47845" heatid="50804" lane="7" entrytime="00:05:26.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                    <SPLIT distance="100" swimtime="00:01:08.31" />
                    <SPLIT distance="150" swimtime="00:01:46.33" />
                    <SPLIT distance="200" swimtime="00:02:24.37" />
                    <SPLIT distance="250" swimtime="00:03:01.85" />
                    <SPLIT distance="300" swimtime="00:03:39.11" />
                    <SPLIT distance="350" swimtime="00:04:15.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="548" reactiontime="+72" swimtime="00:00:28.91" resultid="47846" heatid="50834" lane="1" entrytime="00:00:28.59" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Twaróg" birthdate="2008-04-30" gender="M" nation="POL" license="105801700012" swrid="5249551" athleteid="47829">
              <RESULTS>
                <RESULT eventid="44378" points="409" reactiontime="+85" swimtime="00:01:03.18" resultid="47830" heatid="50672" lane="0" entrytime="00:01:02.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44386" points="357" reactiontime="+71" swimtime="00:02:35.99" resultid="47831" heatid="50704" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                    <SPLIT distance="100" swimtime="00:01:11.00" />
                    <SPLIT distance="150" swimtime="00:01:53.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44390" points="358" reactiontime="+77" swimtime="00:02:40.45" resultid="47832" heatid="50710" lane="9" entrytime="00:02:42.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                    <SPLIT distance="100" swimtime="00:01:17.08" />
                    <SPLIT distance="150" swimtime="00:02:07.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="422" reactiontime="+79" swimtime="00:02:15.90" resultid="47833" heatid="50736" lane="6" entrytime="00:02:16.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.03" />
                    <SPLIT distance="100" swimtime="00:01:05.25" />
                    <SPLIT distance="150" swimtime="00:01:41.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="351" swimtime="00:00:31.57" resultid="47834" heatid="50764" lane="4" entrytime="00:00:31.79" entrycourse="LCM" />
                <RESULT eventid="46294" points="431" reactiontime="+74" swimtime="00:04:51.27" resultid="47835" heatid="50798" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                    <SPLIT distance="100" swimtime="00:01:07.40" />
                    <SPLIT distance="150" swimtime="00:01:46.82" />
                    <SPLIT distance="200" swimtime="00:02:24.41" />
                    <SPLIT distance="250" swimtime="00:03:02.29" />
                    <SPLIT distance="300" swimtime="00:03:39.09" />
                    <SPLIT distance="350" swimtime="00:04:16.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="357" reactiontime="+73" swimtime="00:00:29.45" resultid="47836" heatid="50815" lane="9" entrytime="00:00:30.90" entrycourse="LCM" />
                <RESULT eventid="46306" points="381" reactiontime="+72" swimtime="00:01:08.27" resultid="47837" heatid="50847" lane="5" entrytime="00:01:09.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Zakrzewska" birthdate="2007-07-28" gender="F" nation="POL" license="105801600013" swrid="5214645" athleteid="47847">
              <RESULTS>
                <RESULT eventid="44380" points="399" swimtime="00:01:10.22" resultid="47848" heatid="50683" lane="0" entrytime="00:01:09.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44388" points="265" reactiontime="+64" swimtime="00:03:09.54" resultid="47849" heatid="50706" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                    <SPLIT distance="100" swimtime="00:01:26.29" />
                    <SPLIT distance="150" swimtime="00:02:18.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="323" reactiontime="+72" swimtime="00:00:35.59" resultid="47850" heatid="50775" lane="3" entrytime="00:00:35.35" entrycourse="LCM" />
                <RESULT eventid="46300" points="484" reactiontime="+68" swimtime="00:00:30.13" resultid="47851" heatid="50831" lane="7" entrytime="00:00:30.69" entrycourse="LCM" />
                <RESULT eventid="46308" points="292" reactiontime="+71" swimtime="00:01:23.57" resultid="47852" heatid="50899" lane="8" entrytime="00:01:21.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="354" reactiontime="+68" swimtime="00:00:38.11" resultid="47853" heatid="50903" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Barbara" lastname="Zakrzewska" birthdate="2005-11-26" gender="F" nation="POL" license="105801600016" swrid="5249588" athleteid="47854">
              <RESULTS>
                <RESULT eventid="44380" points="387" reactiontime="+75" swimtime="00:01:10.90" resultid="47855" heatid="50683" lane="8" entrytime="00:01:09.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44388" points="296" reactiontime="+76" swimtime="00:03:02.66" resultid="47856" heatid="50706" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                    <SPLIT distance="100" swimtime="00:01:26.34" />
                    <SPLIT distance="150" swimtime="00:02:15.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="364" reactiontime="+73" swimtime="00:00:34.20" resultid="47857" heatid="50775" lane="0" entrytime="00:00:37.76" entrycourse="LCM" />
                <RESULT eventid="46300" points="428" reactiontime="+73" swimtime="00:00:31.39" resultid="47858" heatid="50829" lane="7" entrytime="00:00:33.52" entrycourse="LCM" />
                <RESULT eventid="46308" points="302" reactiontime="+74" swimtime="00:01:22.69" resultid="47859" heatid="50897" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="331" reactiontime="+58" swimtime="00:00:38.99" resultid="47860" heatid="50906" lane="6" entrytime="00:00:39.70" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="95" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="44401" points="364" reactiontime="+64" swimtime="00:05:22.42" resultid="47881" heatid="50731" lane="7" entrytime="00:05:19.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                    <SPLIT distance="100" swimtime="00:01:23.36" />
                    <SPLIT distance="150" swimtime="00:02:00.30" />
                    <SPLIT distance="200" swimtime="00:02:44.90" />
                    <SPLIT distance="250" swimtime="00:03:22.42" />
                    <SPLIT distance="300" swimtime="00:04:10.75" />
                    <SPLIT distance="350" swimtime="00:04:44.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="47854" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="47838" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="47847" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="47868" number="4" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46291" points="448" reactiontime="+71" swimtime="00:04:34.44" resultid="47882" heatid="50795" lane="8" entrytime="00:04:35.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                    <SPLIT distance="100" swimtime="00:01:09.63" />
                    <SPLIT distance="150" swimtime="00:01:44.83" />
                    <SPLIT distance="200" swimtime="00:02:23.36" />
                    <SPLIT distance="250" swimtime="00:02:55.93" />
                    <SPLIT distance="300" swimtime="00:03:31.99" />
                    <SPLIT distance="350" swimtime="00:04:00.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="47847" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="47868" number="2" reactiontime="+22" />
                    <RELAYPOSITION athleteid="47854" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="47838" number="4" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46316" points="446" reactiontime="+74" swimtime="00:10:03.96" resultid="47883" heatid="50871" lane="3" entrytime="00:09:59.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.26" />
                    <SPLIT distance="100" swimtime="00:01:04.61" />
                    <SPLIT distance="150" swimtime="00:01:40.66" />
                    <SPLIT distance="200" swimtime="00:02:16.10" />
                    <SPLIT distance="250" swimtime="00:02:51.44" />
                    <SPLIT distance="300" swimtime="00:03:32.35" />
                    <SPLIT distance="350" swimtime="00:04:15.20" />
                    <SPLIT distance="400" swimtime="00:04:54.41" />
                    <SPLIT distance="450" swimtime="00:05:28.00" />
                    <SPLIT distance="500" swimtime="00:06:07.40" />
                    <SPLIT distance="550" swimtime="00:06:49.06" />
                    <SPLIT distance="600" swimtime="00:07:28.16" />
                    <SPLIT distance="650" swimtime="00:08:01.14" />
                    <SPLIT distance="700" swimtime="00:08:40.84" />
                    <SPLIT distance="750" swimtime="00:09:23.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="47838" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="47868" number="2" reactiontime="+29" />
                    <RELAYPOSITION athleteid="47854" number="3" reactiontime="+67" />
                    <RELAYPOSITION athleteid="47847" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="05601" nation="POL" region="01" clubid="46475" name="Gminny Klub Pływacki 7 Zdrój Trzebnica">
          <ATHLETES>
            <ATHLETE firstname="Monika" lastname="Michalczuk" birthdate="2008-07-30" gender="F" nation="POL" license="105601600012" swrid="5287611" athleteid="46490">
              <RESULTS>
                <RESULT eventid="44380" points="498" reactiontime="+70" swimtime="00:01:05.21" resultid="46491" heatid="50686" lane="8" entrytime="00:01:04.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="466" reactiontime="+73" swimtime="00:02:25.68" resultid="46492" heatid="50742" lane="6" entrytime="00:02:24.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                    <SPLIT distance="100" swimtime="00:01:10.91" />
                    <SPLIT distance="150" swimtime="00:01:49.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46287" points="459" reactiontime="+61" swimtime="00:10:28.46" resultid="46493" heatid="50791" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                    <SPLIT distance="100" swimtime="00:01:12.25" />
                    <SPLIT distance="150" swimtime="00:01:51.06" />
                    <SPLIT distance="200" swimtime="00:02:30.44" />
                    <SPLIT distance="250" swimtime="00:03:10.14" />
                    <SPLIT distance="300" swimtime="00:03:50.19" />
                    <SPLIT distance="350" swimtime="00:04:30.23" />
                    <SPLIT distance="400" swimtime="00:05:10.11" />
                    <SPLIT distance="450" swimtime="00:05:50.18" />
                    <SPLIT distance="500" swimtime="00:06:29.93" />
                    <SPLIT distance="550" swimtime="00:07:10.45" />
                    <SPLIT distance="600" swimtime="00:07:50.82" />
                    <SPLIT distance="650" swimtime="00:08:31.17" />
                    <SPLIT distance="700" swimtime="00:09:11.07" />
                    <SPLIT distance="750" swimtime="00:09:50.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" status="DNS" swimtime="00:00:00.00" resultid="46494" heatid="50802" lane="0" />
                <RESULT eventid="46300" points="484" reactiontime="+69" swimtime="00:00:30.14" resultid="46495" heatid="50832" lane="7" entrytime="00:00:29.93" entrycourse="LCM" />
                <RESULT eventid="46312" points="420" reactiontime="+77" swimtime="00:00:36.02" resultid="46496" heatid="50907" lane="3" entrytime="00:00:35.80" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Okoń" birthdate="2007-02-22" gender="M" nation="POL" license="105601700009" swrid="5165911" athleteid="46476">
              <RESULTS>
                <RESULT eventid="44378" points="435" reactiontime="+64" swimtime="00:01:01.91" resultid="46477" heatid="50672" lane="5" entrytime="00:01:01.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44390" points="397" reactiontime="+64" swimtime="00:02:35.09" resultid="46478" heatid="50710" lane="8" entrytime="00:02:36.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.06" />
                    <SPLIT distance="100" swimtime="00:01:14.35" />
                    <SPLIT distance="150" swimtime="00:02:00.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="459" reactiontime="+48" swimtime="00:02:12.15" resultid="46479" heatid="50736" lane="4" entrytime="00:02:15.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.57" />
                    <SPLIT distance="100" swimtime="00:01:03.36" />
                    <SPLIT distance="150" swimtime="00:01:38.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46285" points="477" reactiontime="+63" swimtime="00:18:34.67" resultid="46480" heatid="50790" lane="3" entrytime="00:18:44.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.69" />
                    <SPLIT distance="100" swimtime="00:01:05.13" />
                    <SPLIT distance="150" swimtime="00:01:41.06" />
                    <SPLIT distance="200" swimtime="00:02:18.04" />
                    <SPLIT distance="250" swimtime="00:02:55.10" />
                    <SPLIT distance="300" swimtime="00:03:31.94" />
                    <SPLIT distance="350" swimtime="00:04:09.24" />
                    <SPLIT distance="400" swimtime="00:04:46.53" />
                    <SPLIT distance="450" swimtime="00:05:23.96" />
                    <SPLIT distance="500" swimtime="00:06:01.70" />
                    <SPLIT distance="550" swimtime="00:06:39.20" />
                    <SPLIT distance="600" swimtime="00:07:16.83" />
                    <SPLIT distance="650" swimtime="00:07:55.24" />
                    <SPLIT distance="700" swimtime="00:08:32.77" />
                    <SPLIT distance="750" swimtime="00:09:10.17" />
                    <SPLIT distance="800" swimtime="00:09:47.45" />
                    <SPLIT distance="850" swimtime="00:10:25.20" />
                    <SPLIT distance="900" swimtime="00:11:02.46" />
                    <SPLIT distance="950" swimtime="00:11:40.35" />
                    <SPLIT distance="1000" swimtime="00:12:18.24" />
                    <SPLIT distance="1050" swimtime="00:12:56.23" />
                    <SPLIT distance="1100" swimtime="00:13:34.37" />
                    <SPLIT distance="1150" swimtime="00:14:12.37" />
                    <SPLIT distance="1200" swimtime="00:14:50.27" />
                    <SPLIT distance="1250" swimtime="00:15:28.43" />
                    <SPLIT distance="1300" swimtime="00:16:06.46" />
                    <SPLIT distance="1350" swimtime="00:16:43.57" />
                    <SPLIT distance="1400" swimtime="00:17:21.57" />
                    <SPLIT distance="1450" swimtime="00:17:58.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="483" reactiontime="+63" swimtime="00:04:40.42" resultid="46481" heatid="50799" lane="6" entrytime="00:04:48.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.79" />
                    <SPLIT distance="100" swimtime="00:01:04.25" />
                    <SPLIT distance="150" swimtime="00:01:39.95" />
                    <SPLIT distance="200" swimtime="00:02:15.97" />
                    <SPLIT distance="250" swimtime="00:02:52.50" />
                    <SPLIT distance="300" swimtime="00:03:29.15" />
                    <SPLIT distance="350" swimtime="00:04:05.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46302" points="320" reactiontime="+66" swimtime="00:03:04.23" resultid="46482" heatid="50838" lane="7" entrytime="00:04:00.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.52" />
                    <SPLIT distance="100" swimtime="00:01:28.59" />
                    <SPLIT distance="150" swimtime="00:02:16.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Angelika" lastname="Zys" birthdate="2004-03-27" gender="F" nation="POL" license="105601600052" swrid="5088656" athleteid="46497">
              <RESULTS>
                <RESULT eventid="44380" points="431" reactiontime="+88" swimtime="00:01:08.43" resultid="46498" heatid="50679" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44417" points="340" swimtime="00:02:56.61" resultid="46499" heatid="50787" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.51" />
                    <SPLIT distance="100" swimtime="00:01:28.69" />
                    <SPLIT distance="150" swimtime="00:02:14.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="451" reactiontime="+84" swimtime="00:00:30.85" resultid="46500" heatid="50825" lane="9" />
                <RESULT eventid="46312" points="386" reactiontime="+88" swimtime="00:00:37.04" resultid="46501" heatid="50904" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Kunicki" birthdate="2008-01-01" gender="M" nation="POL" athleteid="50872">
              <RESULTS>
                <RESULT eventid="44411" points="243" reactiontime="+76" swimtime="00:00:35.68" resultid="50873" heatid="50757" lane="7" late="yes" />
                <RESULT eventid="46294" points="277" reactiontime="+71" swimtime="00:05:37.34" resultid="50874" heatid="50796" lane="6" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                    <SPLIT distance="100" swimtime="00:01:14.24" />
                    <SPLIT distance="150" swimtime="00:01:57.65" />
                    <SPLIT distance="200" swimtime="00:02:41.79" />
                    <SPLIT distance="250" swimtime="00:03:26.96" />
                    <SPLIT distance="300" swimtime="00:04:11.54" />
                    <SPLIT distance="350" swimtime="00:04:56.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="305" reactiontime="+68" swimtime="00:00:31.06" resultid="50875" heatid="50806" lane="6" late="yes" />
                <RESULT eventid="46310" points="281" reactiontime="+57" swimtime="00:00:36.64" resultid="50876" heatid="50855" lane="6" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antoni" lastname="Tomalik" birthdate="2008-05-12" gender="M" nation="POL" license="105601700014" swrid="5244071" athleteid="46512">
              <RESULTS>
                <RESULT eventid="44394" points="272" reactiontime="+59" swimtime="00:01:19.94" resultid="46513" heatid="50720" lane="1" entrytime="00:01:20.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="270" reactiontime="+64" swimtime="00:02:53.06" resultid="46514" heatid="50782" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.83" />
                    <SPLIT distance="100" swimtime="00:01:24.79" />
                    <SPLIT distance="150" swimtime="00:02:09.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="264" reactiontime="+65" swimtime="00:00:32.59" resultid="46515" heatid="50814" lane="8" entrytime="00:00:32.68" entrycourse="LCM" />
                <RESULT eventid="46310" points="263" reactiontime="+64" swimtime="00:00:37.45" resultid="46516" heatid="50859" lane="7" entrytime="00:00:41.37" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Michalczuk" birthdate="2008-07-30" gender="M" nation="POL" license="105601700011" swrid="5287614" athleteid="46483">
              <RESULTS>
                <RESULT eventid="44378" points="340" reactiontime="+63" swimtime="00:01:07.20" resultid="46484" heatid="50668" lane="2" entrytime="00:01:06.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="262" reactiontime="+79" swimtime="00:01:21.03" resultid="46485" heatid="50719" lane="4" entrytime="00:01:21.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="317" reactiontime="+70" swimtime="00:02:29.54" resultid="46486" heatid="50735" lane="8" entrytime="00:02:27.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                    <SPLIT distance="100" swimtime="00:01:14.05" />
                    <SPLIT distance="150" swimtime="00:01:54.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="323" swimtime="00:05:20.52" resultid="46487" heatid="50796" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                    <SPLIT distance="100" swimtime="00:01:14.00" />
                    <SPLIT distance="150" swimtime="00:01:55.40" />
                    <SPLIT distance="200" swimtime="00:02:37.38" />
                    <SPLIT distance="250" swimtime="00:03:19.60" />
                    <SPLIT distance="300" swimtime="00:04:02.10" />
                    <SPLIT distance="350" swimtime="00:04:43.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="327" reactiontime="+67" swimtime="00:00:30.35" resultid="46488" heatid="50815" lane="7" entrytime="00:00:30.27" entrycourse="LCM" />
                <RESULT eventid="46310" points="256" reactiontime="+73" swimtime="00:00:37.75" resultid="46489" heatid="50859" lane="4" entrytime="00:00:38.07" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Majchrzak" birthdate="2006-10-09" gender="F" nation="POL" license="105601600004" swrid="5281330" athleteid="46502">
              <RESULTS>
                <RESULT eventid="44384" points="545" reactiontime="+75" swimtime="00:00:35.99" resultid="46503" heatid="50701" lane="3" entrytime="00:00:38.78" entrycourse="LCM" />
                <RESULT eventid="44409" points="480" reactiontime="+66" swimtime="00:01:21.89" resultid="46504" heatid="50755" lane="8" entrytime="00:01:22.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="304" reactiontime="+72" swimtime="00:00:36.31" resultid="46505" heatid="50774" lane="5" entrytime="00:00:38.17" entrycourse="LCM" />
                <RESULT eventid="46304" points="395" reactiontime="+75" swimtime="00:03:09.52" resultid="46506" heatid="50840" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.91" />
                    <SPLIT distance="100" swimtime="00:01:29.94" />
                    <SPLIT distance="150" swimtime="00:02:20.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zofia" lastname="Kunicka" birthdate="2008-01-01" gender="F" nation="POL" athleteid="50877">
              <RESULTS>
                <RESULT eventid="46300" points="283" reactiontime="+90" swimtime="00:00:36.05" resultid="50878" heatid="50823" lane="6" late="yes" />
                <RESULT eventid="44405" reactiontime="+89" status="DNF" swimtime="00:00:00.00" resultid="50879" heatid="50740" lane="0" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                    <SPLIT distance="100" swimtime="00:01:26.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="266" reactiontime="+71" swimtime="00:00:41.93" resultid="50880" heatid="50903" lane="2" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksander" lastname="Tomalik" birthdate="2006-04-05" gender="M" nation="POL" license="105601700015" swrid="5212908" athleteid="46507">
              <RESULTS>
                <RESULT eventid="44394" points="330" reactiontime="+71" swimtime="00:01:14.97" resultid="46508" heatid="50721" lane="7" entrytime="00:01:15.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="330" reactiontime="+71" swimtime="00:02:41.93" resultid="46509" heatid="50783" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.48" />
                    <SPLIT distance="100" swimtime="00:01:19.86" />
                    <SPLIT distance="150" swimtime="00:02:01.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="326" reactiontime="+79" swimtime="00:00:30.36" resultid="46510" heatid="50813" lane="9" entrytime="00:00:34.95" entrycourse="LCM" />
                <RESULT eventid="46310" points="315" reactiontime="+70" swimtime="00:00:35.27" resultid="46511" heatid="50859" lane="5" entrytime="00:00:39.29" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01507" nation="POL" region="07" clubid="48385" name="UKS MOS w Opolu">
          <ATHLETES>
            <ATHLETE firstname="Oliwier" lastname="Sosnowski" birthdate="2005-07-07" gender="M" nation="POL" license="101507700068" swrid="5168603" athleteid="48390">
              <RESULTS>
                <RESULT eventid="44378" points="542" reactiontime="+68" swimtime="00:00:57.53" resultid="48391" heatid="50674" lane="3" entrytime="00:00:58.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="491" reactiontime="+66" swimtime="00:02:09.27" resultid="48392" heatid="50738" lane="0" entrytime="00:02:10.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.48" />
                    <SPLIT distance="100" swimtime="00:01:02.43" />
                    <SPLIT distance="150" swimtime="00:01:36.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="484" reactiontime="+68" swimtime="00:00:26.63" resultid="48393" heatid="50818" lane="5" entrytime="00:00:26.75" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Rakowska" birthdate="2006-02-07" gender="F" nation="POL" license="101507600070" swrid="4973679" athleteid="48457">
              <RESULTS>
                <RESULT eventid="44392" points="627" reactiontime="+66" swimtime="00:02:27.30" resultid="48458" heatid="50716" lane="5" entrytime="00:02:27.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                    <SPLIT distance="100" swimtime="00:01:11.47" />
                    <SPLIT distance="150" swimtime="00:01:54.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="636" reactiontime="+73" swimtime="00:02:11.32" resultid="48459" heatid="50744" lane="3" entrytime="00:02:10.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                    <SPLIT distance="100" swimtime="00:01:05.00" />
                    <SPLIT distance="150" swimtime="00:01:39.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46287" points="574" reactiontime="+70" swimtime="00:09:43.18" resultid="48460" heatid="50791" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.97" />
                    <SPLIT distance="100" swimtime="00:01:09.27" />
                    <SPLIT distance="150" swimtime="00:01:46.16" />
                    <SPLIT distance="200" swimtime="00:02:23.87" />
                    <SPLIT distance="250" swimtime="00:03:00.77" />
                    <SPLIT distance="300" swimtime="00:03:38.13" />
                    <SPLIT distance="350" swimtime="00:04:15.08" />
                    <SPLIT distance="400" swimtime="00:04:52.18" />
                    <SPLIT distance="450" swimtime="00:05:29.00" />
                    <SPLIT distance="500" swimtime="00:06:06.22" />
                    <SPLIT distance="550" swimtime="00:06:43.13" />
                    <SPLIT distance="600" swimtime="00:07:20.52" />
                    <SPLIT distance="650" swimtime="00:07:57.27" />
                    <SPLIT distance="700" swimtime="00:08:34.91" />
                    <SPLIT distance="750" swimtime="00:09:10.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="594" reactiontime="+72" swimtime="00:04:41.29" resultid="48461" heatid="50805" lane="6" entrytime="00:04:43.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                    <SPLIT distance="100" swimtime="00:01:07.88" />
                    <SPLIT distance="150" swimtime="00:01:44.26" />
                    <SPLIT distance="200" swimtime="00:02:20.71" />
                    <SPLIT distance="250" swimtime="00:02:56.81" />
                    <SPLIT distance="300" swimtime="00:03:32.82" />
                    <SPLIT distance="350" swimtime="00:04:08.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cezary" lastname="Górowski" birthdate="2004-08-28" gender="M" nation="POL" license="101507700038" swrid="5117194" athleteid="48403">
              <RESULTS>
                <RESULT eventid="44378" points="483" reactiontime="+74" swimtime="00:00:59.78" resultid="48404" heatid="50673" lane="0" entrytime="00:01:00.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="486" reactiontime="+73" swimtime="00:02:09.71" resultid="48405" heatid="50737" lane="5" entrytime="00:02:11.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.84" />
                    <SPLIT distance="100" swimtime="00:01:02.84" />
                    <SPLIT distance="150" swimtime="00:01:36.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="477" reactiontime="+65" swimtime="00:04:41.53" resultid="48406" heatid="50799" lane="4" entrytime="00:04:38.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.86" />
                    <SPLIT distance="100" swimtime="00:01:04.85" />
                    <SPLIT distance="150" swimtime="00:01:40.18" />
                    <SPLIT distance="200" swimtime="00:02:16.31" />
                    <SPLIT distance="250" swimtime="00:02:52.82" />
                    <SPLIT distance="300" swimtime="00:03:30.56" />
                    <SPLIT distance="350" swimtime="00:04:06.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marco" lastname="Czaja" birthdate="2003-12-09" gender="M" nation="POL" license="101507700002" swrid="4926616" athleteid="48466">
              <RESULTS>
                <RESULT eventid="44394" points="633" reactiontime="+65" swimtime="00:01:00.36" resultid="48467" heatid="50723" lane="3" entrytime="00:01:01.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46310" points="670" reactiontime="+61" swimtime="00:00:27.42" resultid="48468" heatid="50862" lane="6" entrytime="00:00:28.06" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Pasternak" birthdate="2005-05-19" gender="M" nation="POL" license="101507700057" swrid="5112218" athleteid="48407">
              <RESULTS>
                <RESULT eventid="44378" points="492" reactiontime="+66" swimtime="00:00:59.39" resultid="48408" heatid="50663" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="517" reactiontime="+60" swimtime="00:00:27.74" resultid="48409" heatid="50762" lane="9" entrytime="00:00:48.33" entrycourse="LCM" />
                <RESULT eventid="46298" points="501" reactiontime="+64" swimtime="00:00:26.32" resultid="48410" heatid="50812" lane="0" entrytime="00:00:37.90" entrycourse="LCM" />
                <RESULT eventid="46310" points="471" reactiontime="+63" swimtime="00:00:30.84" resultid="48411" heatid="50859" lane="8" entrytime="00:00:43.47" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulina" lastname="Jaśniecka" birthdate="2007-05-31" gender="F" nation="POL" license="101507600067" swrid="5269049" athleteid="48431">
              <RESULTS>
                <RESULT eventid="44380" points="443" reactiontime="+76" swimtime="00:01:07.80" resultid="48432" heatid="50684" lane="1" entrytime="00:01:07.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46287" points="463" reactiontime="+76" swimtime="00:10:26.41" resultid="48433" heatid="50791" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                    <SPLIT distance="100" swimtime="00:01:12.51" />
                    <SPLIT distance="150" swimtime="00:01:51.82" />
                    <SPLIT distance="200" swimtime="00:02:31.21" />
                    <SPLIT distance="250" swimtime="00:03:10.93" />
                    <SPLIT distance="300" swimtime="00:03:50.28" />
                    <SPLIT distance="350" swimtime="00:04:29.90" />
                    <SPLIT distance="400" swimtime="00:05:09.60" />
                    <SPLIT distance="450" swimtime="00:05:49.14" />
                    <SPLIT distance="500" swimtime="00:06:28.53" />
                    <SPLIT distance="550" swimtime="00:07:09.02" />
                    <SPLIT distance="600" swimtime="00:07:49.57" />
                    <SPLIT distance="650" swimtime="00:08:29.59" />
                    <SPLIT distance="700" swimtime="00:09:09.87" />
                    <SPLIT distance="750" swimtime="00:09:48.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="460" reactiontime="+77" swimtime="00:05:06.31" resultid="48434" heatid="50804" lane="6" entrytime="00:05:03.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                    <SPLIT distance="100" swimtime="00:01:11.82" />
                    <SPLIT distance="150" swimtime="00:01:51.16" />
                    <SPLIT distance="200" swimtime="00:02:30.36" />
                    <SPLIT distance="250" swimtime="00:03:09.77" />
                    <SPLIT distance="300" swimtime="00:03:49.16" />
                    <SPLIT distance="350" swimtime="00:04:28.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maksymilian" lastname="Topolnicki" birthdate="2006-04-08" gender="M" nation="POL" license="101507700094" swrid="4918010" athleteid="48449">
              <RESULTS>
                <RESULT eventid="44390" points="516" reactiontime="+56" swimtime="00:02:22.11" resultid="48450" heatid="50710" lane="4" entrytime="00:02:28.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.29" />
                    <SPLIT distance="100" swimtime="00:01:09.13" />
                    <SPLIT distance="150" swimtime="00:01:50.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="497" reactiontime="+70" swimtime="00:02:08.75" resultid="48451" heatid="50732" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                    <SPLIT distance="100" swimtime="00:01:02.55" />
                    <SPLIT distance="150" swimtime="00:01:36.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="527" reactiontime="+62" swimtime="00:00:25.88" resultid="48452" heatid="50810" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Żaba" birthdate="2005-09-19" gender="M" nation="POL" license="101507700013" swrid="5085199" athleteid="48453">
              <RESULTS>
                <RESULT eventid="44390" points="519" reactiontime="+76" swimtime="00:02:21.79" resultid="48454" heatid="50710" lane="3" entrytime="00:02:28.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.09" />
                    <SPLIT distance="100" swimtime="00:01:09.77" />
                    <SPLIT distance="150" swimtime="00:01:50.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="482" reactiontime="+77" swimtime="00:01:12.52" resultid="48455" heatid="50749" lane="7" entrytime="00:01:18.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46302" points="507" reactiontime="+78" swimtime="00:02:38.15" resultid="48456" heatid="50839" lane="9" entrytime="00:02:41.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.21" />
                    <SPLIT distance="100" swimtime="00:01:16.31" />
                    <SPLIT distance="150" swimtime="00:01:57.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alicja" lastname="Czuryło" birthdate="2007-10-12" gender="F" nation="POL" license="101507600060" swrid="5269054" athleteid="48482">
              <RESULTS>
                <RESULT eventid="44396" points="362" reactiontime="+86" swimtime="00:01:20.71" resultid="48483" heatid="50724" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="364" reactiontime="+80" swimtime="00:00:37.78" resultid="48484" heatid="50904" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Szymczykowski" birthdate="2003-05-12" gender="M" nation="POL" license="101507700005" swrid="5097700" athleteid="48441">
              <RESULTS>
                <RESULT eventid="44386" points="609" reactiontime="+77" swimtime="00:02:10.62" resultid="48442" heatid="50705" lane="3" entrytime="00:02:11.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.91" />
                    <SPLIT distance="100" swimtime="00:01:01.81" />
                    <SPLIT distance="150" swimtime="00:01:36.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="632" reactiontime="+70" swimtime="00:01:58.82" resultid="48443" heatid="50739" lane="2" entrytime="00:01:59.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.71" />
                    <SPLIT distance="100" swimtime="00:00:58.11" />
                    <SPLIT distance="150" swimtime="00:01:28.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="628" reactiontime="+71" swimtime="00:04:16.91" resultid="48444" heatid="50800" lane="6" entrytime="00:04:18.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.42" />
                    <SPLIT distance="100" swimtime="00:01:01.81" />
                    <SPLIT distance="150" swimtime="00:01:34.70" />
                    <SPLIT distance="200" swimtime="00:02:07.91" />
                    <SPLIT distance="250" swimtime="00:02:41.23" />
                    <SPLIT distance="300" swimtime="00:03:14.55" />
                    <SPLIT distance="350" swimtime="00:03:46.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Trentkiewicz" birthdate="2004-03-07" gender="F" nation="POL" license="101507600009" swrid="5013985" athleteid="48477">
              <RESULTS>
                <RESULT eventid="44396" points="721" reactiontime="+53" swimtime="00:01:04.18" resultid="48478" heatid="50728" lane="5" entrytime="00:01:03.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="615" reactiontime="+65" swimtime="00:00:28.72" resultid="48479" heatid="50779" lane="5" entrytime="00:00:29.00" entrycourse="LCM" />
                <RESULT eventid="46300" points="615" reactiontime="+64" swimtime="00:00:27.82" resultid="48480" heatid="50834" lane="9" entrytime="00:00:28.73" entrycourse="LCM" />
                <RESULT eventid="46312" points="725" reactiontime="+56" swimtime="00:00:30.03" resultid="48481" heatid="50909" lane="3" entrytime="00:00:29.95" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mikołaj" lastname="Adamek" birthdate="2004-05-01" gender="M" nation="POL" license="101507700054" swrid="5082344" athleteid="48394">
              <RESULTS>
                <RESULT eventid="44378" points="545" reactiontime="+71" swimtime="00:00:57.41" resultid="48395" heatid="50674" lane="1" entrytime="00:00:58.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="512" reactiontime="+71" swimtime="00:02:07.45" resultid="48396" heatid="50737" lane="4" entrytime="00:02:10.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.29" />
                    <SPLIT distance="100" swimtime="00:01:01.18" />
                    <SPLIT distance="150" swimtime="00:01:34.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="480" reactiontime="+72" swimtime="00:00:26.69" resultid="48397" heatid="50819" lane="0" entrytime="00:00:26.62" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Gilowska" birthdate="2006-05-13" gender="F" nation="POL" license="101507600059" swrid="5250810" athleteid="48474">
              <RESULTS>
                <RESULT eventid="44396" points="387" reactiontime="+82" swimtime="00:01:18.96" resultid="48475" heatid="50727" lane="7" entrytime="00:01:15.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="443" reactiontime="+73" swimtime="00:00:35.38" resultid="48476" heatid="50908" lane="1" entrytime="00:00:34.68" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Szczygieł" birthdate="2007-06-19" gender="M" nation="POL" license="101507700058" swrid="5120220" athleteid="48462">
              <RESULTS>
                <RESULT eventid="44394" points="372" reactiontime="+75" swimtime="00:01:12.04" resultid="48463" heatid="50721" lane="4" entrytime="00:01:12.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="374" reactiontime="+75" swimtime="00:02:35.33" resultid="48464" heatid="50783" lane="3" entrytime="00:02:37.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.88" />
                    <SPLIT distance="100" swimtime="00:01:17.18" />
                    <SPLIT distance="150" swimtime="00:01:57.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46310" points="366" reactiontime="+74" swimtime="00:00:33.53" resultid="48465" heatid="50860" lane="2" entrytime="00:00:33.56" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patryk" lastname="Podgórski" birthdate="2003-03-11" gender="M" nation="POL" license="101507700004" swrid="4947386" athleteid="48469">
              <RESULTS>
                <RESULT eventid="44394" points="544" reactiontime="+61" swimtime="00:01:03.50" resultid="48470" heatid="50723" lane="6" entrytime="00:01:03.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="521" reactiontime="+60" swimtime="00:02:19.02" resultid="48471" heatid="50784" lane="6" entrytime="00:02:15.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                    <SPLIT distance="100" swimtime="00:01:07.39" />
                    <SPLIT distance="150" swimtime="00:01:43.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="524" reactiontime="+71" swimtime="00:00:25.92" resultid="48472" heatid="50817" lane="5" entrytime="00:00:27.83" entrycourse="LCM" />
                <RESULT eventid="46310" points="514" reactiontime="+61" swimtime="00:00:29.95" resultid="48473" heatid="50862" lane="2" entrytime="00:00:29.26" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Gucwa" birthdate="2007-08-16" gender="M" nation="POL" license="101507700032" swrid="4995598" athleteid="48412">
              <RESULTS>
                <RESULT eventid="44378" points="349" reactiontime="+77" swimtime="00:01:06.59" resultid="48413" heatid="50669" lane="3" entrytime="00:01:05.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="330" reactiontime="+67" swimtime="00:00:32.20" resultid="48414" heatid="50763" lane="6" entrytime="00:00:33.38" entrycourse="LCM" />
                <RESULT eventid="46298" points="359" reactiontime="+61" swimtime="00:00:29.40" resultid="48415" heatid="50808" lane="1" />
                <RESULT eventid="46310" points="287" reactiontime="+70" swimtime="00:00:36.37" resultid="48416" heatid="50858" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Chłąd" birthdate="2006-05-22" gender="F" nation="POL" license="101507600039" swrid="5165387" athleteid="48426">
              <RESULTS>
                <RESULT eventid="44380" points="578" reactiontime="+81" swimtime="00:01:02.07" resultid="48427" heatid="50688" lane="0" entrytime="00:01:01.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="619" reactiontime="+77" swimtime="00:02:12.53" resultid="48428" heatid="50744" lane="1" entrytime="00:02:13.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                    <SPLIT distance="100" swimtime="00:01:05.25" />
                    <SPLIT distance="150" swimtime="00:01:39.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="552" reactiontime="+76" swimtime="00:04:48.24" resultid="48429" heatid="50805" lane="2" entrytime="00:04:43.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                    <SPLIT distance="100" swimtime="00:01:08.07" />
                    <SPLIT distance="150" swimtime="00:01:44.33" />
                    <SPLIT distance="200" swimtime="00:02:21.14" />
                    <SPLIT distance="250" swimtime="00:02:57.37" />
                    <SPLIT distance="300" swimtime="00:03:34.22" />
                    <SPLIT distance="350" swimtime="00:04:11.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="539" reactiontime="+80" swimtime="00:00:29.08" resultid="48430" heatid="50833" lane="6" entrytime="00:00:29.10" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jagoda" lastname="Justyńska" birthdate="2007-08-14" gender="F" nation="POL" license="101507600093" swrid="4918049" athleteid="48417">
              <RESULTS>
                <RESULT eventid="44380" points="467" reactiontime="+78" swimtime="00:01:06.62" resultid="48418" heatid="50684" lane="3" entrytime="00:01:06.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="472" reactiontime="+80" swimtime="00:02:25.05" resultid="48419" heatid="50742" lane="9" entrytime="00:02:29.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="100" swimtime="00:01:09.82" />
                    <SPLIT distance="150" swimtime="00:01:48.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46287" points="397" reactiontime="+79" swimtime="00:10:59.47" resultid="48420" heatid="50791" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.01" />
                    <SPLIT distance="100" swimtime="00:01:12.77" />
                    <SPLIT distance="150" swimtime="00:01:53.10" />
                    <SPLIT distance="200" swimtime="00:02:34.76" />
                    <SPLIT distance="250" swimtime="00:03:16.64" />
                    <SPLIT distance="300" swimtime="00:03:58.76" />
                    <SPLIT distance="350" swimtime="00:04:40.76" />
                    <SPLIT distance="400" swimtime="00:05:22.97" />
                    <SPLIT distance="450" swimtime="00:06:05.49" />
                    <SPLIT distance="500" swimtime="00:06:48.38" />
                    <SPLIT distance="550" swimtime="00:07:31.06" />
                    <SPLIT distance="600" swimtime="00:08:13.55" />
                    <SPLIT distance="650" swimtime="00:08:55.41" />
                    <SPLIT distance="700" swimtime="00:09:37.60" />
                    <SPLIT distance="750" swimtime="00:10:19.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="514" reactiontime="+75" swimtime="00:00:29.53" resultid="48421" heatid="50829" lane="5" entrytime="00:00:33.07" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Iga" lastname="Kosacka" birthdate="2003-11-21" gender="F" nation="POL" license="101507600017" swrid="5013984" athleteid="48422">
              <RESULTS>
                <RESULT eventid="44380" status="DNS" swimtime="00:00:00.00" resultid="48423" heatid="50685" lane="0" entrytime="00:01:06.02" entrycourse="LCM" />
                <RESULT eventid="44413" status="DNS" swimtime="00:00:00.00" resultid="48424" heatid="50778" lane="6" entrytime="00:00:30.96" entrycourse="LCM" />
                <RESULT eventid="46300" status="DNS" swimtime="00:00:00.00" resultid="48425" heatid="50832" lane="5" entrytime="00:00:29.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hanna" lastname="Mielnik" birthdate="2007-05-01" gender="F" nation="POL" license="101507600065" swrid="4918007" athleteid="48445">
              <RESULTS>
                <RESULT eventid="44388" points="545" reactiontime="+70" swimtime="00:02:29.12" resultid="48446" heatid="50706" lane="4" entrytime="00:02:35.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.84" />
                    <SPLIT distance="100" swimtime="00:01:11.00" />
                    <SPLIT distance="150" swimtime="00:01:49.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44409" points="629" reactiontime="+74" swimtime="00:01:14.82" resultid="48447" heatid="50756" lane="6" entrytime="00:01:16.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46304" points="589" reactiontime="+74" swimtime="00:02:45.86" resultid="48448" heatid="50843" lane="2" entrytime="00:02:47.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.73" />
                    <SPLIT distance="100" swimtime="00:01:21.19" />
                    <SPLIT distance="150" swimtime="00:02:05.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Polok" birthdate="2007-08-29" gender="F" nation="POL" license="101507600066" swrid="4918052" athleteid="48435">
              <RESULTS>
                <RESULT eventid="44384" points="435" reactiontime="+68" swimtime="00:00:38.80" resultid="48436" heatid="50701" lane="6" entrytime="00:00:39.30" entrycourse="LCM" />
                <RESULT eventid="44392" points="437" reactiontime="+58" swimtime="00:02:46.08" resultid="48437" heatid="50712" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                    <SPLIT distance="100" swimtime="00:01:23.88" />
                    <SPLIT distance="150" swimtime="00:02:08.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44409" points="444" reactiontime="+68" swimtime="00:01:24.02" resultid="48438" heatid="50752" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="333" reactiontime="+67" swimtime="00:00:35.24" resultid="48439" heatid="50770" lane="5" />
                <RESULT eventid="46304" points="452" reactiontime="+67" swimtime="00:03:01.26" resultid="48440" heatid="50843" lane="9" entrytime="00:03:00.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.76" />
                    <SPLIT distance="100" swimtime="00:01:26.47" />
                    <SPLIT distance="150" swimtime="00:02:14.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zofia" lastname="Bobrowska" birthdate="2007-09-24" gender="F" nation="POL" license="101507600014" swrid="4133153" athleteid="48485">
              <RESULTS>
                <RESULT eventid="44413" points="380" reactiontime="+70" swimtime="00:00:33.70" resultid="48486" heatid="50776" lane="5" entrytime="00:00:33.68" entrycourse="LCM" />
                <RESULT eventid="46287" points="423" reactiontime="+73" swimtime="00:10:45.45" resultid="48487" heatid="50792" lane="7" entrytime="00:12:18.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.15" />
                    <SPLIT distance="100" swimtime="00:01:17.25" />
                    <SPLIT distance="150" swimtime="00:01:57.95" />
                    <SPLIT distance="200" swimtime="00:02:39.19" />
                    <SPLIT distance="250" swimtime="00:03:19.63" />
                    <SPLIT distance="300" swimtime="00:04:01.10" />
                    <SPLIT distance="350" swimtime="00:04:42.32" />
                    <SPLIT distance="400" swimtime="00:05:24.02" />
                    <SPLIT distance="450" swimtime="00:06:04.89" />
                    <SPLIT distance="500" swimtime="00:06:45.72" />
                    <SPLIT distance="550" swimtime="00:07:26.74" />
                    <SPLIT distance="600" swimtime="00:08:07.63" />
                    <SPLIT distance="650" swimtime="00:08:47.59" />
                    <SPLIT distance="700" swimtime="00:09:27.61" />
                    <SPLIT distance="750" swimtime="00:10:07.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46308" points="328" reactiontime="+76" swimtime="00:01:20.44" resultid="48488" heatid="50900" lane="0" entrytime="00:01:16.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Baranek" birthdate="2004-10-24" gender="M" nation="POL" license="101507700001" swrid="5097697" athleteid="48398">
              <RESULTS>
                <RESULT eventid="44378" points="636" reactiontime="+72" swimtime="00:00:54.53" resultid="48399" heatid="50676" lane="5" entrytime="00:00:54.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="556" reactiontime="+75" swimtime="00:02:04.02" resultid="48400" heatid="50739" lane="8" entrytime="00:02:02.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.36" />
                    <SPLIT distance="100" swimtime="00:00:59.83" />
                    <SPLIT distance="150" swimtime="00:01:32.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="541" reactiontime="+71" swimtime="00:00:27.33" resultid="48401" heatid="50766" lane="6" entrytime="00:00:29.23" entrycourse="LCM" />
                <RESULT eventid="46298" points="576" reactiontime="+72" swimtime="00:00:25.13" resultid="48402" heatid="50820" lane="5" entrytime="00:00:25.97" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Korpacki" birthdate="2006-09-20" gender="M" nation="POL" license="101507700029" swrid="5250927" athleteid="48386">
              <RESULTS>
                <RESULT eventid="44378" points="519" reactiontime="+63" swimtime="00:00:58.34" resultid="48387" heatid="50670" lane="6" entrytime="00:01:03.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="475" reactiontime="+62" swimtime="00:00:28.54" resultid="48388" heatid="50763" lane="5" entrytime="00:00:32.99" entrycourse="LCM" />
                <RESULT eventid="46306" points="458" reactiontime="+63" swimtime="00:01:04.19" resultid="48389" heatid="50847" lane="2" entrytime="00:01:10.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03801" nation="POL" region="01" clubid="48103" name="UKS Delfinek Legnica">
          <ATHLETES>
            <ATHLETE firstname="Dominik" lastname="Kuleta" birthdate="2008-08-05" gender="M" nation="POL" license="103801700081" swrid="5250892" athleteid="48145">
              <RESULTS>
                <RESULT eventid="44394" status="DNS" swimtime="00:00:00.00" resultid="48146" heatid="50720" lane="9" entrytime="00:01:21.22" entrycourse="LCM" />
                <RESULT eventid="44415" status="DNS" swimtime="00:00:00.00" resultid="48147" heatid="50781" lane="5" />
                <RESULT eventid="46310" status="DNS" swimtime="00:00:00.00" resultid="48148" heatid="50859" lane="1" entrytime="00:00:42.72" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Konarska" birthdate="2005-07-28" gender="F" nation="POL" license="103801600074" swrid="5250941" athleteid="48154">
              <RESULTS>
                <RESULT eventid="44396" points="353" reactiontime="+65" swimtime="00:01:21.40" resultid="48155" heatid="50726" lane="8" entrytime="00:01:22.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="310" reactiontime="+73" swimtime="00:00:36.06" resultid="48156" heatid="50776" lane="1" entrytime="00:00:34.93" entrycourse="LCM" />
                <RESULT eventid="44417" points="299" reactiontime="+63" swimtime="00:03:04.30" resultid="48157" heatid="50787" lane="4" entrytime="00:03:03.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.16" />
                    <SPLIT distance="100" swimtime="00:01:29.09" />
                    <SPLIT distance="150" swimtime="00:02:17.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="318" reactiontime="+77" swimtime="00:05:46.29" resultid="48158" heatid="50801" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.39" />
                    <SPLIT distance="100" swimtime="00:01:18.28" />
                    <SPLIT distance="150" swimtime="00:02:03.01" />
                    <SPLIT distance="200" swimtime="00:02:47.69" />
                    <SPLIT distance="250" swimtime="00:03:33.33" />
                    <SPLIT distance="300" swimtime="00:04:18.34" />
                    <SPLIT distance="350" swimtime="00:05:03.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="406" reactiontime="+59" swimtime="00:00:36.41" resultid="48159" heatid="50906" lane="8" entrytime="00:00:41.04" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Drożdż" birthdate="2005-08-03" gender="F" nation="POL" license="103801600042" swrid="5071690" athleteid="48133">
              <RESULTS>
                <RESULT eventid="44388" points="263" reactiontime="+68" swimtime="00:03:09.95" resultid="48134" heatid="50706" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.38" />
                    <SPLIT distance="100" swimtime="00:01:27.00" />
                    <SPLIT distance="150" swimtime="00:02:19.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="404" reactiontime="+65" swimtime="00:00:33.04" resultid="48135" heatid="50777" lane="7" entrytime="00:00:33.15" entrycourse="LCM" />
                <RESULT eventid="46300" points="460" reactiontime="+62" swimtime="00:00:30.65" resultid="48136" heatid="50831" lane="9" entrytime="00:00:31.05" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Wiśniewska" birthdate="2007-06-23" gender="F" nation="POL" license="103801600085" swrid="5001949" athleteid="48104">
              <RESULTS>
                <RESULT eventid="44380" points="366" reactiontime="+82" swimtime="00:01:12.26" resultid="48105" heatid="50682" lane="3" entrytime="00:01:10.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="381" reactiontime="+79" swimtime="00:00:33.68" resultid="48106" heatid="50776" lane="2" entrytime="00:00:34.36" entrycourse="LCM" />
                <RESULT eventid="44417" points="235" reactiontime="+74" swimtime="00:03:19.61" resultid="48107" heatid="50787" lane="3" entrytime="00:03:17.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.56" />
                    <SPLIT distance="100" swimtime="00:01:39.23" />
                    <SPLIT distance="150" swimtime="00:02:30.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46308" points="339" reactiontime="+78" swimtime="00:01:19.54" resultid="48108" heatid="50898" lane="7" entrytime="00:01:27.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Hoszowska" birthdate="2007-01-14" gender="F" nation="POL" license="103801600064" swrid="5166039" athleteid="48109">
              <RESULTS>
                <RESULT eventid="44380" points="269" reactiontime="+66" swimtime="00:01:20.05" resultid="48110" heatid="50680" lane="7" entrytime="00:01:20.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="244" reactiontime="+69" swimtime="00:00:39.08" resultid="48111" heatid="50773" lane="8" />
                <RESULT eventid="46300" points="315" reactiontime="+70" swimtime="00:00:34.76" resultid="48112" heatid="50824" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Parszeniew" birthdate="2007-09-18" gender="M" nation="POL" license="103801700087" swrid="5193000" athleteid="48117">
              <RESULTS>
                <RESULT eventid="44382" points="253" reactiontime="+73" swimtime="00:00:41.02" resultid="48118" heatid="50693" lane="8" entrytime="00:00:42.30" entrycourse="LCM" />
                <RESULT eventid="44411" points="283" reactiontime="+75" swimtime="00:00:33.92" resultid="48119" heatid="50763" lane="1" entrytime="00:00:34.42" entrycourse="LCM" />
                <RESULT eventid="46298" points="293" reactiontime="+75" swimtime="00:00:31.48" resultid="48120" heatid="50814" lane="3" entrytime="00:00:31.87" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Skowron" birthdate="2007-08-10" gender="M" nation="POL" license="103801700090" swrid="4834347" athleteid="48141">
              <RESULTS>
                <RESULT eventid="44394" points="389" reactiontime="+69" swimtime="00:01:10.97" resultid="48142" heatid="50721" lane="2" entrytime="00:01:15.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="325" reactiontime="+70" swimtime="00:02:42.66" resultid="48143" heatid="50783" lane="2" entrytime="00:02:40.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.25" />
                    <SPLIT distance="100" swimtime="00:01:18.12" />
                    <SPLIT distance="150" swimtime="00:02:01.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46310" points="392" reactiontime="+60" swimtime="00:00:32.79" resultid="48144" heatid="50860" lane="7" entrytime="00:00:35.04" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Chrenowski" birthdate="2004-03-11" gender="M" nation="POL" license="103801700040" swrid="4858830" athleteid="48137">
              <RESULTS>
                <RESULT eventid="44390" points="439" reactiontime="+66" swimtime="00:02:29.96" resultid="48138" heatid="50709" lane="3" entrytime="00:02:46.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.89" />
                    <SPLIT distance="100" swimtime="00:01:06.95" />
                    <SPLIT distance="150" swimtime="00:01:54.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="407" reactiontime="+68" swimtime="00:01:16.75" resultid="48139" heatid="50745" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="541" reactiontime="+64" swimtime="00:00:25.65" resultid="48140" heatid="50818" lane="3" entrytime="00:00:26.78" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrianna" lastname="Radziwon" birthdate="2006-02-24" gender="F" nation="POL" license="103801600054" swrid="5173448" athleteid="48121">
              <RESULTS>
                <RESULT eventid="44384" points="544" reactiontime="+64" swimtime="00:00:36.01" resultid="48122" heatid="50702" lane="7" entrytime="00:00:36.53" entrycourse="LCM" />
                <RESULT eventid="44409" points="463" reactiontime="+65" swimtime="00:01:22.85" resultid="48123" heatid="50755" lane="9" entrytime="00:01:23.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46304" points="457" reactiontime="+66" swimtime="00:03:00.58" resultid="48124" heatid="50842" lane="6" entrytime="00:03:09.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.26" />
                    <SPLIT distance="100" swimtime="00:01:25.46" />
                    <SPLIT distance="150" swimtime="00:02:12.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Gałęza" birthdate="2004-01-23" gender="F" nation="POL" license="103801600092" swrid="4858766" athleteid="48149">
              <RESULTS>
                <RESULT eventid="44396" points="518" reactiontime="+67" swimtime="00:01:11.67" resultid="48150" heatid="50727" lane="3" entrytime="00:01:14.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44417" points="466" reactiontime="+72" swimtime="00:02:38.99" resultid="48151" heatid="50788" lane="1" entrytime="00:02:38.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                    <SPLIT distance="100" swimtime="00:01:18.01" />
                    <SPLIT distance="150" swimtime="00:01:59.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="530" reactiontime="+68" swimtime="00:00:29.24" resultid="48152" heatid="50832" lane="6" entrytime="00:00:29.90" entrycourse="LCM" />
                <RESULT eventid="46312" points="547" reactiontime="+63" swimtime="00:00:32.97" resultid="48153" heatid="50908" lane="5" entrytime="00:00:32.89" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Wołczak" birthdate="2004-02-10" gender="M" nation="POL" license="103801700039" swrid="4858855" athleteid="48129">
              <RESULTS>
                <RESULT eventid="44386" points="250" reactiontime="+59" swimtime="00:02:55.62" resultid="48130" heatid="50704" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                    <SPLIT distance="100" swimtime="00:01:15.71" />
                    <SPLIT distance="150" swimtime="00:02:04.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="391" reactiontime="+66" swimtime="00:00:30.44" resultid="48131" heatid="50765" lane="1" entrytime="00:00:30.87" entrycourse="LCM" />
                <RESULT eventid="46294" points="277" reactiontime="+68" swimtime="00:05:37.22" resultid="48132" heatid="50798" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.67" />
                    <SPLIT distance="100" swimtime="00:01:13.26" />
                    <SPLIT distance="150" swimtime="00:01:55.98" />
                    <SPLIT distance="200" swimtime="00:02:40.48" />
                    <SPLIT distance="250" swimtime="00:03:25.03" />
                    <SPLIT distance="300" swimtime="00:04:10.25" />
                    <SPLIT distance="350" swimtime="00:04:54.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aniela" lastname="Pietrukiewicz" birthdate="2005-07-14" gender="F" nation="POL" license="103801600137" swrid="4858847" athleteid="48125">
              <RESULTS>
                <RESULT eventid="44384" points="275" reactiontime="+93" swimtime="00:00:45.19" resultid="48126" heatid="50698" lane="5" />
                <RESULT eventid="44417" points="239" reactiontime="+81" swimtime="00:03:18.63" resultid="48127" heatid="50785" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.54" />
                    <SPLIT distance="150" swimtime="00:02:28.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" status="DNS" swimtime="00:00:00.00" resultid="48128" heatid="50904" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Pawlik" birthdate="2004-10-04" gender="M" nation="POL" license="103801700096" swrid="4858859" athleteid="48113">
              <RESULTS>
                <RESULT eventid="44382" points="290" reactiontime="+66" swimtime="00:00:39.18" resultid="48114" heatid="50693" lane="7" entrytime="00:00:39.19" entrycourse="LCM" />
                <RESULT eventid="44415" points="240" reactiontime="+63" swimtime="00:03:00.00" resultid="48115" heatid="50783" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.47" />
                    <SPLIT distance="100" swimtime="00:01:27.41" />
                    <SPLIT distance="150" swimtime="00:02:15.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="362" reactiontime="+61" swimtime="00:00:29.32" resultid="48116" heatid="50815" lane="5" entrytime="00:00:29.81" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04901" nation="POL" region="01" clubid="46715" name="KS Neptun Świdnica">
          <ATHLETES>
            <ATHLETE firstname="Kinga" lastname="Kamieniarz" birthdate="2005-04-09" gender="F" nation="POL" license="104901600046" swrid="5166049" athleteid="46756">
              <RESULTS>
                <RESULT eventid="44384" points="597" reactiontime="+69" swimtime="00:00:34.91" resultid="46757" heatid="50702" lane="3" entrytime="00:00:35.79" entrycourse="LCM" />
                <RESULT eventid="44409" points="574" reactiontime="+61" swimtime="00:01:17.15" resultid="46758" heatid="50756" lane="7" entrytime="00:01:17.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46304" points="609" reactiontime="+64" swimtime="00:02:44.03" resultid="46759" heatid="50843" lane="3" entrytime="00:02:45.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.72" />
                    <SPLIT distance="100" swimtime="00:01:18.27" />
                    <SPLIT distance="150" swimtime="00:02:01.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Lęga" birthdate="2005-04-20" gender="F" nation="POL" license="104901600009" swrid="4995402" athleteid="46732">
              <RESULTS>
                <RESULT eventid="44380" points="550" reactiontime="+72" swimtime="00:01:03.11" resultid="46733" heatid="50686" lane="1" entrytime="00:01:04.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="528" reactiontime="+75" swimtime="00:02:19.72" resultid="46734" heatid="50743" lane="2" entrytime="00:02:18.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                    <SPLIT distance="100" swimtime="00:01:07.55" />
                    <SPLIT distance="150" swimtime="00:01:44.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46287" points="515" reactiontime="+74" swimtime="00:10:04.44" resultid="46735" heatid="50792" lane="6" entrytime="00:10:16.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.63" />
                    <SPLIT distance="100" swimtime="00:01:09.46" />
                    <SPLIT distance="150" swimtime="00:01:47.16" />
                    <SPLIT distance="200" swimtime="00:02:25.47" />
                    <SPLIT distance="250" swimtime="00:03:04.05" />
                    <SPLIT distance="300" swimtime="00:03:42.36" />
                    <SPLIT distance="350" swimtime="00:04:20.99" />
                    <SPLIT distance="400" swimtime="00:04:59.43" />
                    <SPLIT distance="450" swimtime="00:05:37.81" />
                    <SPLIT distance="500" swimtime="00:06:16.33" />
                    <SPLIT distance="550" swimtime="00:06:54.18" />
                    <SPLIT distance="600" swimtime="00:07:32.92" />
                    <SPLIT distance="650" swimtime="00:08:11.48" />
                    <SPLIT distance="700" swimtime="00:08:50.08" />
                    <SPLIT distance="750" swimtime="00:09:27.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="502" reactiontime="+71" swimtime="00:04:57.34" resultid="46736" heatid="50805" lane="9" entrytime="00:04:56.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="100" swimtime="00:01:08.95" />
                    <SPLIT distance="150" swimtime="00:01:46.60" />
                    <SPLIT distance="200" swimtime="00:02:25.17" />
                    <SPLIT distance="250" swimtime="00:03:03.61" />
                    <SPLIT distance="300" swimtime="00:03:41.86" />
                    <SPLIT distance="350" swimtime="00:04:20.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="513" reactiontime="+66" swimtime="00:00:29.56" resultid="46737" heatid="50833" lane="0" entrytime="00:00:29.47" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kamila" lastname="Świdnicka" birthdate="2006-06-07" gender="F" nation="POL" license="104901600068" swrid="4995331" athleteid="46738">
              <RESULTS>
                <RESULT eventid="44380" points="539" reactiontime="+80" swimtime="00:01:03.52" resultid="46739" heatid="50686" lane="6" entrytime="00:01:04.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="507" reactiontime="+76" swimtime="00:02:21.60" resultid="46740" heatid="50743" lane="7" entrytime="00:02:19.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                    <SPLIT distance="100" swimtime="00:01:08.27" />
                    <SPLIT distance="150" swimtime="00:01:45.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46287" status="DNS" swimtime="00:00:00.00" resultid="46741" heatid="50792" lane="1" entrytime="00:12:27.26" entrycourse="LCM" />
                <RESULT eventid="46296" points="497" reactiontime="+76" swimtime="00:04:58.38" resultid="46742" heatid="50804" lane="5" entrytime="00:05:01.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                    <SPLIT distance="100" swimtime="00:01:09.85" />
                    <SPLIT distance="150" swimtime="00:01:48.32" />
                    <SPLIT distance="200" swimtime="00:02:27.02" />
                    <SPLIT distance="250" swimtime="00:03:05.75" />
                    <SPLIT distance="300" swimtime="00:03:44.19" />
                    <SPLIT distance="350" swimtime="00:04:23.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="508" reactiontime="+77" swimtime="00:00:29.66" resultid="46743" heatid="50831" lane="5" entrytime="00:00:30.16" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hubert" lastname="Hołdys" birthdate="2007-04-06" gender="M" nation="POL" license="104901700038" swrid="5341352" athleteid="46716">
              <RESULTS>
                <RESULT eventid="44378" points="339" reactiontime="+69" swimtime="00:01:07.25" resultid="46717" heatid="50668" lane="8" entrytime="00:01:07.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="274" reactiontime="+70" swimtime="00:00:39.92" resultid="46718" heatid="50693" lane="1" entrytime="00:00:41.28" entrycourse="LCM" />
                <RESULT eventid="44403" points="331" reactiontime="+51" swimtime="00:02:27.41" resultid="46719" heatid="50734" lane="4" entrytime="00:02:29.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.93" />
                    <SPLIT distance="100" swimtime="00:01:11.39" />
                    <SPLIT distance="150" swimtime="00:01:49.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="323" reactiontime="+50" swimtime="00:00:30.47" resultid="46720" heatid="50814" lane="4" entrytime="00:00:31.11" entrycourse="LCM" />
                <RESULT eventid="46306" points="235" reactiontime="+63" swimtime="00:01:20.14" resultid="46721" heatid="50846" lane="8" entrytime="00:01:21.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Florczak" birthdate="2007-03-02" gender="M" nation="POL" license="104901700026" swrid="5194172" athleteid="46750">
              <RESULTS>
                <RESULT eventid="44382" points="458" reactiontime="+63" swimtime="00:00:33.65" resultid="46751" heatid="50695" lane="9" entrytime="00:00:33.02" entrycourse="LCM" />
                <RESULT eventid="44407" points="410" reactiontime="+66" swimtime="00:01:16.51" resultid="46752" heatid="50749" lane="4" entrytime="00:01:13.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="445" reactiontime="+66" swimtime="00:00:29.15" resultid="46753" heatid="50766" lane="8" entrytime="00:00:29.77" entrycourse="LCM" />
                <RESULT eventid="46298" points="444" reactiontime="+64" swimtime="00:00:27.39" resultid="46754" heatid="50815" lane="0" entrytime="00:00:30.42" entrycourse="LCM" />
                <RESULT eventid="46302" points="394" reactiontime="+68" swimtime="00:02:52.00" resultid="46755" heatid="50839" lane="0" entrytime="00:02:40.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.96" />
                    <SPLIT distance="100" swimtime="00:01:21.86" />
                    <SPLIT distance="150" swimtime="00:02:07.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Kowalik" birthdate="2006-06-07" gender="M" nation="POL" license="104901700016" swrid="5165949" athleteid="46722">
              <RESULTS>
                <RESULT eventid="44378" points="418" reactiontime="+71" swimtime="00:01:02.73" resultid="46723" heatid="50671" lane="7" entrytime="00:01:03.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="394" reactiontime="+58" swimtime="00:02:19.03" resultid="46724" heatid="50735" lane="4" entrytime="00:02:22.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                    <SPLIT distance="100" swimtime="00:01:06.13" />
                    <SPLIT distance="150" swimtime="00:01:42.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="295" reactiontime="+71" swimtime="00:00:33.45" resultid="46725" heatid="50762" lane="1" entrytime="00:00:41.00" entrycourse="LCM" />
                <RESULT eventid="46294" points="418" reactiontime="+55" swimtime="00:04:54.12" resultid="46726" heatid="50798" lane="4" entrytime="00:05:03.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                    <SPLIT distance="100" swimtime="00:01:07.00" />
                    <SPLIT distance="150" swimtime="00:01:44.12" />
                    <SPLIT distance="200" swimtime="00:02:21.84" />
                    <SPLIT distance="250" swimtime="00:03:00.19" />
                    <SPLIT distance="300" swimtime="00:03:38.91" />
                    <SPLIT distance="350" swimtime="00:04:17.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="353" reactiontime="+70" swimtime="00:00:29.57" resultid="46727" heatid="50813" lane="7" entrytime="00:00:33.40" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcel" lastname="Borkowski" birthdate="2007-02-06" gender="M" nation="POL" license="104901700035" swrid="5353542" athleteid="46775">
              <RESULTS>
                <RESULT eventid="44386" points="446" reactiontime="+69" swimtime="00:02:24.89" resultid="46776" heatid="50705" lane="2" entrytime="00:02:29.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.75" />
                    <SPLIT distance="100" swimtime="00:01:07.70" />
                    <SPLIT distance="150" swimtime="00:01:45.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46285" points="457" reactiontime="+70" swimtime="00:18:50.66" resultid="46778" heatid="50790" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.30" />
                    <SPLIT distance="100" swimtime="00:01:11.25" />
                    <SPLIT distance="150" swimtime="00:01:49.04" />
                    <SPLIT distance="200" swimtime="00:02:26.63" />
                    <SPLIT distance="250" swimtime="00:03:04.37" />
                    <SPLIT distance="300" swimtime="00:03:41.87" />
                    <SPLIT distance="350" swimtime="00:04:19.37" />
                    <SPLIT distance="400" swimtime="00:04:57.21" />
                    <SPLIT distance="450" swimtime="00:05:34.73" />
                    <SPLIT distance="500" swimtime="00:06:12.45" />
                    <SPLIT distance="550" swimtime="00:06:50.19" />
                    <SPLIT distance="600" swimtime="00:07:27.85" />
                    <SPLIT distance="650" swimtime="00:08:05.76" />
                    <SPLIT distance="700" swimtime="00:08:43.40" />
                    <SPLIT distance="750" swimtime="00:09:21.61" />
                    <SPLIT distance="800" swimtime="00:09:59.72" />
                    <SPLIT distance="850" swimtime="00:10:38.00" />
                    <SPLIT distance="900" swimtime="00:11:16.43" />
                    <SPLIT distance="950" swimtime="00:11:54.79" />
                    <SPLIT distance="1000" swimtime="00:12:33.12" />
                    <SPLIT distance="1050" swimtime="00:13:11.76" />
                    <SPLIT distance="1100" swimtime="00:13:49.77" />
                    <SPLIT distance="1150" swimtime="00:14:27.75" />
                    <SPLIT distance="1200" swimtime="00:15:06.13" />
                    <SPLIT distance="1250" swimtime="00:15:43.86" />
                    <SPLIT distance="1300" swimtime="00:16:21.76" />
                    <SPLIT distance="1350" swimtime="00:16:59.87" />
                    <SPLIT distance="1400" swimtime="00:17:37.78" />
                    <SPLIT distance="1450" swimtime="00:18:14.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="458" reactiontime="+57" swimtime="00:04:45.37" resultid="46779" heatid="50799" lane="7" entrytime="00:04:49.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.59" />
                    <SPLIT distance="100" swimtime="00:01:05.22" />
                    <SPLIT distance="150" swimtime="00:01:41.18" />
                    <SPLIT distance="200" swimtime="00:02:17.60" />
                    <SPLIT distance="250" swimtime="00:02:55.02" />
                    <SPLIT distance="300" swimtime="00:03:31.99" />
                    <SPLIT distance="350" swimtime="00:04:09.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46306" points="385" reactiontime="+61" swimtime="00:01:08.02" resultid="50896" heatid="50844" lane="9" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Jaros" birthdate="2007-05-17" gender="F" nation="POL" license="104901600024" swrid="5088569" athleteid="46781">
              <RESULTS>
                <RESULT eventid="44388" points="448" reactiontime="+69" swimtime="00:02:39.14" resultid="46782" heatid="50706" lane="3" entrytime="00:02:44.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                    <SPLIT distance="100" swimtime="00:01:14.92" />
                    <SPLIT distance="150" swimtime="00:01:56.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46287" points="472" reactiontime="+72" swimtime="00:10:22.40" resultid="46785" heatid="50792" lane="2" entrytime="00:10:33.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="100" swimtime="00:01:13.14" />
                    <SPLIT distance="150" swimtime="00:01:52.69" />
                    <SPLIT distance="200" swimtime="00:02:31.73" />
                    <SPLIT distance="250" swimtime="00:03:10.94" />
                    <SPLIT distance="300" swimtime="00:03:49.84" />
                    <SPLIT distance="350" swimtime="00:04:28.93" />
                    <SPLIT distance="400" swimtime="00:05:08.30" />
                    <SPLIT distance="450" swimtime="00:05:46.34" />
                    <SPLIT distance="500" swimtime="00:06:25.60" />
                    <SPLIT distance="550" swimtime="00:07:05.66" />
                    <SPLIT distance="600" swimtime="00:07:45.67" />
                    <SPLIT distance="650" swimtime="00:08:25.68" />
                    <SPLIT distance="700" swimtime="00:09:05.44" />
                    <SPLIT distance="750" swimtime="00:09:44.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="480" reactiontime="+69" swimtime="00:05:01.82" resultid="46786" heatid="50804" lane="2" entrytime="00:05:04.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                    <SPLIT distance="100" swimtime="00:01:11.42" />
                    <SPLIT distance="150" swimtime="00:01:49.28" />
                    <SPLIT distance="200" swimtime="00:02:28.02" />
                    <SPLIT distance="250" swimtime="00:03:07.51" />
                    <SPLIT distance="300" swimtime="00:03:46.67" />
                    <SPLIT distance="350" swimtime="00:04:25.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46308" points="460" reactiontime="+71" swimtime="00:01:11.82" resultid="46787" heatid="50900" lane="7" entrytime="00:01:12.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Lęga" birthdate="2007-01-30" gender="F" nation="POL" license="104901600023" swrid="5088558" athleteid="46788">
              <RESULTS>
                <RESULT eventid="44396" points="431" reactiontime="+73" swimtime="00:01:16.18" resultid="46789" heatid="50727" lane="6" entrytime="00:01:14.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44417" points="434" reactiontime="+74" swimtime="00:02:42.83" resultid="46790" heatid="50788" lane="8" entrytime="00:02:41.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.67" />
                    <SPLIT distance="100" swimtime="00:01:20.25" />
                    <SPLIT distance="150" swimtime="00:02:02.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46308" points="321" reactiontime="+77" swimtime="00:01:21.02" resultid="46791" heatid="50900" lane="9" entrytime="00:01:17.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="430" reactiontime="+67" swimtime="00:00:35.73" resultid="46792" heatid="50907" lane="4" entrytime="00:00:35.45" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Gut" birthdate="2008-09-12" gender="M" nation="POL" license="104901700039" swrid="5341349" athleteid="46728">
              <RESULTS>
                <RESULT eventid="44378" points="286" reactiontime="+73" swimtime="00:01:11.18" resultid="46729" heatid="50666" lane="1" entrytime="00:01:23.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="279" reactiontime="+77" swimtime="00:02:36.06" resultid="46730" heatid="50733" lane="7" entrytime="00:02:41.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                    <SPLIT distance="100" swimtime="00:01:16.41" />
                    <SPLIT distance="150" swimtime="00:01:57.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="287" reactiontime="+67" swimtime="00:00:31.69" resultid="46731" heatid="50812" lane="6" entrytime="00:00:36.07" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kinga" lastname="Ścisłowicz" birthdate="2007-04-16" gender="F" nation="POL" license="104901600025" swrid="5165935" athleteid="46766">
              <RESULTS>
                <RESULT eventid="44384" points="441" reactiontime="+74" swimtime="00:00:38.60" resultid="46767" heatid="50701" lane="2" entrytime="00:00:39.59" entrycourse="LCM" />
                <RESULT eventid="44392" points="422" reactiontime="+82" swimtime="00:02:48.13" resultid="46768" heatid="50714" lane="6" entrytime="00:02:51.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                    <SPLIT distance="100" swimtime="00:01:25.17" />
                    <SPLIT distance="150" swimtime="00:02:09.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44409" points="456" reactiontime="+74" swimtime="00:01:23.26" resultid="46769" heatid="50755" lane="1" entrytime="00:01:22.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46304" points="456" reactiontime="+53" swimtime="00:03:00.65" resultid="46770" heatid="50842" lane="4" entrytime="00:03:00.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.99" />
                    <SPLIT distance="100" swimtime="00:01:28.40" />
                    <SPLIT distance="150" swimtime="00:02:14.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martyna" lastname="Kuśnierz" birthdate="2006-02-11" gender="F" nation="POL" license="104901600029" swrid="5165939" athleteid="46760">
              <RESULTS>
                <RESULT eventid="44384" points="472" reactiontime="+77" swimtime="00:00:37.76" resultid="46761" heatid="50702" lane="0" entrytime="00:00:37.68" entrycourse="LCM" />
                <RESULT eventid="44409" points="439" reactiontime="+68" swimtime="00:01:24.37" resultid="46762" heatid="50754" lane="5" entrytime="00:01:24.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="399" reactiontime="+72" swimtime="00:00:33.17" resultid="46763" heatid="50777" lane="8" entrytime="00:00:33.35" entrycourse="LCM" />
                <RESULT eventid="46300" points="436" reactiontime="+67" swimtime="00:00:31.20" resultid="46764" heatid="50830" lane="1" entrytime="00:00:31.95" entrycourse="LCM" />
                <RESULT eventid="46304" points="412" reactiontime="+74" swimtime="00:03:06.88" resultid="46765" heatid="50842" lane="3" entrytime="00:03:05.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.61" />
                    <SPLIT distance="100" swimtime="00:01:30.57" />
                    <SPLIT distance="150" swimtime="00:02:19.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Wrona" birthdate="2008-09-03" gender="F" nation="POL" license="104901600034" swrid="5272089" athleteid="46771">
              <RESULTS>
                <RESULT eventid="44384" points="205" reactiontime="+75" swimtime="00:00:49.84" resultid="46772" heatid="50699" lane="6" entrytime="00:00:55.18" entrycourse="LCM" />
                <RESULT eventid="44409" points="192" reactiontime="+75" swimtime="00:01:51.12" resultid="46773" heatid="50752" lane="3" entrytime="00:01:53.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="280" reactiontime="+65" swimtime="00:00:36.14" resultid="46774" heatid="50828" lane="8" entrytime="00:00:38.61" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04601" nation="POL" region="01" clubid="47957" name="UKS ,,SZAFIR&apos;&apos; Wałbrzych">
          <ATHLETES>
            <ATHLETE firstname="Mateusz" lastname="Dębski" birthdate="2004-03-16" gender="M" nation="POL" license="104601700041" swrid="5028296" athleteid="48009">
              <RESULTS>
                <RESULT eventid="44382" points="298" reactiontime="+78" swimtime="00:00:38.82" resultid="48010" heatid="50691" lane="1" />
                <RESULT eventid="44407" points="286" reactiontime="+76" swimtime="00:01:26.25" resultid="48011" heatid="50745" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="402" reactiontime="+80" swimtime="00:00:28.33" resultid="48012" heatid="50811" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Draus" birthdate="2007-03-19" gender="M" nation="POL" license="104601700024" swrid="5260095" athleteid="47958">
              <RESULTS>
                <RESULT eventid="44378" points="393" reactiontime="+73" swimtime="00:01:04.00" resultid="47959" heatid="50670" lane="2" entrytime="00:01:03.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="253" reactiontime="+72" swimtime="00:00:41.02" resultid="47960" heatid="50690" lane="8" />
                <RESULT eventid="44403" points="344" reactiontime="+71" swimtime="00:02:25.54" resultid="47961" heatid="50735" lane="6" entrytime="00:02:25.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.20" />
                    <SPLIT distance="100" swimtime="00:01:11.26" />
                    <SPLIT distance="150" swimtime="00:01:48.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="302" reactiontime="+69" swimtime="00:00:33.18" resultid="47962" heatid="50758" lane="2" />
                <RESULT eventid="46298" points="370" reactiontime="+69" swimtime="00:00:29.11" resultid="47963" heatid="50806" lane="5" />
                <RESULT eventid="46306" points="228" reactiontime="+78" swimtime="00:01:20.97" resultid="47964" heatid="50846" lane="7" entrytime="00:01:18.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Łąpieś" birthdate="2004-09-05" gender="F" nation="POL" license="104601600015" swrid="5194146" athleteid="48031">
              <RESULTS>
                <RESULT eventid="44396" points="492" reactiontime="+71" swimtime="00:01:12.91" resultid="48032" heatid="50727" lane="8" entrytime="00:01:16.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44417" points="439" reactiontime="+89" swimtime="00:02:42.19" resultid="48033" heatid="50787" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.71" />
                    <SPLIT distance="100" swimtime="00:01:19.78" />
                    <SPLIT distance="150" swimtime="00:02:02.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="529" reactiontime="+79" swimtime="00:00:29.25" resultid="48034" heatid="50830" lane="5" entrytime="00:00:31.14" entrycourse="LCM" />
                <RESULT eventid="46312" points="520" reactiontime="+79" swimtime="00:00:33.53" resultid="48035" heatid="50907" lane="2" entrytime="00:00:35.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miłosz" lastname="Kowalski" birthdate="2008-01-19" gender="M" nation="POL" license="104601700033" swrid="5296038" athleteid="47984">
              <RESULTS>
                <RESULT eventid="44378" points="297" reactiontime="+72" swimtime="00:01:10.26" resultid="47985" heatid="50666" lane="7" entrytime="00:01:21.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="295" reactiontime="+83" swimtime="00:01:17.88" resultid="47986" heatid="50719" lane="5" entrytime="00:01:21.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="223" reactiontime="+76" swimtime="00:01:33.75" resultid="47987" heatid="50747" lane="9" entrytime="00:01:42.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="289" reactiontime="+74" swimtime="00:00:31.60" resultid="47988" heatid="50810" lane="3" />
                <RESULT eventid="46310" points="270" reactiontime="+77" swimtime="00:00:37.12" resultid="47989" heatid="50859" lane="2" entrytime="00:00:41.10" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Kaszuba" birthdate="2008-02-21" gender="M" nation="POL" license="104601700076" swrid="5296035" athleteid="47990">
              <RESULTS>
                <RESULT eventid="44378" points="249" reactiontime="+72" swimtime="00:01:14.55" resultid="47991" heatid="50667" lane="0" entrytime="00:01:12.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="161" reactiontime="+65" swimtime="00:01:35.12" resultid="47992" heatid="50719" lane="1" entrytime="00:01:28.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="228" reactiontime="+68" swimtime="00:00:36.42" resultid="47993" heatid="50761" lane="7" />
                <RESULT eventid="46298" points="238" reactiontime="+72" swimtime="00:00:33.73" resultid="47994" heatid="50811" lane="1" />
                <RESULT eventid="46310" points="169" reactiontime="+84" swimtime="00:00:43.33" resultid="47995" heatid="50857" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Klaudia" lastname="Żurawska" birthdate="2002-10-19" gender="F" nation="POL" license="104601600016" swrid="5108824" athleteid="48017">
              <RESULTS>
                <RESULT eventid="44396" points="441" reactiontime="+71" swimtime="00:01:15.59" resultid="48019" heatid="50727" lane="1" entrytime="00:01:16.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="447" reactiontime="+62" swimtime="00:00:31.94" resultid="48020" heatid="50777" lane="5" entrytime="00:00:32.52" entrycourse="LCM" />
                <RESULT eventid="44417" points="388" reactiontime="+81" swimtime="00:02:49.06" resultid="48021" heatid="50786" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.40" />
                    <SPLIT distance="100" swimtime="00:01:21.82" />
                    <SPLIT distance="150" swimtime="00:02:05.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="467" reactiontime="+70" swimtime="00:00:30.50" resultid="48023" heatid="50831" lane="8" entrytime="00:00:30.84" entrycourse="LCM" />
                <RESULT eventid="46312" points="439" reactiontime="+83" swimtime="00:00:35.48" resultid="48025" heatid="50907" lane="7" entrytime="00:00:35.92" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Mrzygłód" birthdate="2005-03-05" gender="M" nation="POL" license="104601700020" swrid="5083100" athleteid="47979">
              <RESULTS>
                <RESULT eventid="44378" points="556" reactiontime="+67" swimtime="00:00:57.02" resultid="47980" heatid="50675" lane="0" entrytime="00:00:57.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="516" reactiontime="+67" swimtime="00:02:07.14" resultid="47981" heatid="50738" lane="1" entrytime="00:02:08.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.80" />
                    <SPLIT distance="100" swimtime="00:01:01.30" />
                    <SPLIT distance="150" swimtime="00:01:35.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="472" reactiontime="+68" swimtime="00:00:26.84" resultid="47982" heatid="50818" lane="6" entrytime="00:00:26.84" entrycourse="LCM" />
                <RESULT eventid="46306" status="DNS" swimtime="00:00:00.00" resultid="47983" heatid="50848" lane="8" entrytime="00:01:07.34" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Dębska" birthdate="2007-07-10" gender="F" nation="POL" license="104601600058" swrid="5296046" athleteid="48026">
              <RESULTS>
                <RESULT eventid="44396" points="305" reactiontime="+73" swimtime="00:01:25.45" resultid="48027" heatid="50725" lane="0" entrytime="00:01:27.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="252" reactiontime="+60" swimtime="00:00:38.65" resultid="48028" heatid="50772" lane="2" />
                <RESULT eventid="46300" points="393" reactiontime="+45" swimtime="00:00:32.29" resultid="48029" heatid="50826" lane="0" />
                <RESULT eventid="46312" points="316" reactiontime="+70" swimtime="00:00:39.59" resultid="48030" heatid="50905" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Kołomańska" birthdate="2008-09-20" gender="F" nation="POL" license="104601600030" swrid="5166070" athleteid="47996">
              <RESULTS>
                <RESULT eventid="44380" points="439" reactiontime="+56" swimtime="00:01:08.01" resultid="47997" heatid="50683" lane="5" entrytime="00:01:08.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="399" reactiontime="+66" swimtime="00:02:33.35" resultid="47998" heatid="50741" lane="7" entrytime="00:02:34.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.11" />
                    <SPLIT distance="100" swimtime="00:01:14.54" />
                    <SPLIT distance="150" swimtime="00:01:54.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="450" reactiontime="+55" swimtime="00:00:30.88" resultid="47999" heatid="50827" lane="9" />
                <RESULT eventid="46308" points="231" reactiontime="+61" swimtime="00:01:30.30" resultid="48000" heatid="50898" lane="8" entrytime="00:01:29.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Róża" lastname="Garba" birthdate="2008-11-30" gender="F" nation="POL" license="104601600031" swrid="5244075" athleteid="48001">
              <RESULTS>
                <RESULT eventid="44380" points="395" reactiontime="+75" swimtime="00:01:10.47" resultid="48002" heatid="50682" lane="6" entrytime="00:01:10.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44396" points="341" reactiontime="+87" swimtime="00:01:22.34" resultid="48003" heatid="50726" lane="7" entrytime="00:01:21.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="400" reactiontime="+71" swimtime="00:00:33.15" resultid="48004" heatid="50776" lane="7" entrytime="00:00:34.68" entrycourse="LCM" />
                <RESULT eventid="44417" points="324" reactiontime="+67" swimtime="00:02:59.53" resultid="48005" heatid="50787" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.82" />
                    <SPLIT distance="100" swimtime="00:01:30.18" />
                    <SPLIT distance="150" swimtime="00:02:16.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="419" reactiontime="+61" swimtime="00:00:31.62" resultid="48006" heatid="50826" lane="2" />
                <RESULT eventid="46308" points="350" reactiontime="+63" swimtime="00:01:18.66" resultid="48007" heatid="50899" lane="5" entrytime="00:01:17.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="371" reactiontime="+76" swimtime="00:00:37.54" resultid="48008" heatid="50906" lane="3" entrytime="00:00:39.38" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antoni" lastname="Laszkiewicz" birthdate="2007-02-01" gender="M" nation="POL" license="104601700006" swrid="5200973" athleteid="47971">
              <RESULTS>
                <RESULT eventid="44378" points="362" reactiontime="+67" swimtime="00:01:05.78" resultid="47972" heatid="50669" lane="7" entrytime="00:01:05.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="275" reactiontime="+60" swimtime="00:00:39.87" resultid="47973" heatid="50689" lane="4" />
                <RESULT eventid="44403" points="332" reactiontime="+68" swimtime="00:02:27.16" resultid="47974" heatid="50734" lane="2" entrytime="00:02:30.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.51" />
                    <SPLIT distance="100" swimtime="00:01:13.66" />
                    <SPLIT distance="150" swimtime="00:01:52.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="275" reactiontime="+63" swimtime="00:01:27.38" resultid="47975" heatid="50747" lane="5" entrytime="00:01:31.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="331" reactiontime="+66" swimtime="00:00:32.17" resultid="47976" heatid="50760" lane="1" />
                <RESULT eventid="46298" points="351" reactiontime="+67" swimtime="00:00:29.62" resultid="47977" heatid="50813" lane="6" entrytime="00:00:33.34" entrycourse="LCM" />
                <RESULT eventid="46306" points="200" reactiontime="+70" swimtime="00:01:24.60" resultid="47978" heatid="50845" lane="3" entrytime="00:01:24.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Król" birthdate="2005-06-16" gender="M" nation="POL" license="104601700047" swrid="5190446" athleteid="47965">
              <RESULTS>
                <RESULT eventid="44378" points="438" reactiontime="+75" swimtime="00:01:01.74" resultid="47966" heatid="50665" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="401" reactiontime="+71" swimtime="00:00:35.18" resultid="47967" heatid="50690" lane="9" />
                <RESULT eventid="44394" points="330" reactiontime="+70" swimtime="00:01:14.98" resultid="47968" heatid="50719" lane="6" entrytime="00:01:23.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="377" reactiontime="+75" swimtime="00:01:18.71" resultid="47969" heatid="50746" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="417" reactiontime="+78" swimtime="00:00:27.97" resultid="47970" heatid="50810" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06414" nation="POL" region="14" clubid="47543" name="MKS Piaseczno">
          <ATHLETES>
            <ATHLETE firstname="Krzysztof" lastname="Kasprzak" birthdate="2005-04-21" gender="M" nation="POL" license="106414700217" swrid="5006560" athleteid="47544">
              <RESULTS>
                <RESULT eventid="44378" points="558" reactiontime="+64" swimtime="00:00:56.95" resultid="47545" heatid="50675" lane="5" entrytime="00:00:56.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="494" reactiontime="+60" swimtime="00:01:05.55" resultid="47546" heatid="50723" lane="7" entrytime="00:01:05.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="508" reactiontime="+64" swimtime="00:02:07.82" resultid="47547" heatid="50738" lane="7" entrytime="00:02:06.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.88" />
                    <SPLIT distance="100" swimtime="00:01:02.04" />
                    <SPLIT distance="150" swimtime="00:01:36.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="509" swimtime="00:00:27.88" resultid="47548" heatid="50767" lane="7" entrytime="00:00:28.73" entrycourse="LCM" />
                <RESULT eventid="46294" points="503" reactiontime="+67" swimtime="00:04:36.62" resultid="47549" heatid="50800" lane="1" entrytime="00:04:34.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.73" />
                    <SPLIT distance="100" swimtime="00:01:04.87" />
                    <SPLIT distance="150" swimtime="00:01:39.78" />
                    <SPLIT distance="200" swimtime="00:02:15.81" />
                    <SPLIT distance="250" swimtime="00:02:51.38" />
                    <SPLIT distance="300" swimtime="00:03:26.96" />
                    <SPLIT distance="350" swimtime="00:04:02.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="565" reactiontime="+64" swimtime="00:00:25.29" resultid="47550" heatid="50821" lane="6" entrytime="00:00:25.22" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zofia" lastname="Har" birthdate="2004-09-14" gender="F" nation="POL" license="106414600132" swrid="4980369" athleteid="47577">
              <RESULTS>
                <RESULT eventid="44384" points="602" reactiontime="+75" swimtime="00:00:34.80" resultid="47578" heatid="50702" lane="6" entrytime="00:00:36.07" entrycourse="LCM" />
                <RESULT eventid="44409" points="554" reactiontime="+64" swimtime="00:01:18.05" resultid="47579" heatid="50756" lane="9" entrytime="00:01:18.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="537" reactiontime="+74" swimtime="00:00:29.12" resultid="47580" heatid="50825" lane="7" />
                <RESULT eventid="46304" points="599" reactiontime="+72" swimtime="00:02:45.01" resultid="47581" heatid="50843" lane="7" entrytime="00:02:47.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                    <SPLIT distance="100" swimtime="00:01:18.89" />
                    <SPLIT distance="150" swimtime="00:02:01.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwia" lastname="Samoraj" birthdate="2005-02-25" gender="F" nation="POL" license="106414600107" swrid="5036197" athleteid="47565">
              <RESULTS>
                <RESULT eventid="44380" points="582" reactiontime="+68" swimtime="00:01:01.93" resultid="47566" heatid="50688" lane="9" entrytime="00:01:01.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="640" reactiontime="+72" swimtime="00:02:11.05" resultid="47567" heatid="50744" lane="6" entrytime="00:02:11.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                    <SPLIT distance="100" swimtime="00:01:03.63" />
                    <SPLIT distance="150" swimtime="00:01:37.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46287" points="594" reactiontime="+74" swimtime="00:09:36.62" resultid="47568" heatid="50792" lane="5" entrytime="00:09:41.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                    <SPLIT distance="100" swimtime="00:01:07.96" />
                    <SPLIT distance="150" swimtime="00:01:43.73" />
                    <SPLIT distance="200" swimtime="00:02:19.58" />
                    <SPLIT distance="250" swimtime="00:02:55.24" />
                    <SPLIT distance="300" swimtime="00:03:31.38" />
                    <SPLIT distance="350" swimtime="00:04:07.62" />
                    <SPLIT distance="400" swimtime="00:04:44.32" />
                    <SPLIT distance="450" swimtime="00:05:20.62" />
                    <SPLIT distance="500" swimtime="00:05:57.55" />
                    <SPLIT distance="550" swimtime="00:06:34.41" />
                    <SPLIT distance="600" swimtime="00:07:10.67" />
                    <SPLIT distance="650" swimtime="00:07:48.10" />
                    <SPLIT distance="700" swimtime="00:08:25.00" />
                    <SPLIT distance="750" swimtime="00:09:01.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="591" reactiontime="+74" swimtime="00:04:41.76" resultid="47569" heatid="50805" lane="3" entrytime="00:04:41.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.66" />
                    <SPLIT distance="100" swimtime="00:01:06.31" />
                    <SPLIT distance="150" swimtime="00:01:41.80" />
                    <SPLIT distance="200" swimtime="00:02:17.73" />
                    <SPLIT distance="250" swimtime="00:02:53.67" />
                    <SPLIT distance="300" swimtime="00:03:30.44" />
                    <SPLIT distance="350" swimtime="00:04:07.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46308" points="489" reactiontime="+71" swimtime="00:01:10.38" resultid="47570" heatid="50901" lane="9" entrytime="00:01:09.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Tkacz" birthdate="2005-05-09" gender="M" nation="POL" license="106414700071" swrid="5020373" athleteid="47558">
              <RESULTS>
                <RESULT eventid="44378" points="646" reactiontime="+71" swimtime="00:00:54.26" resultid="47559" heatid="50676" lane="6" entrytime="00:00:55.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="549" reactiontime="+70" swimtime="00:00:31.69" resultid="47560" heatid="50695" lane="2" entrytime="00:00:31.79" entrycourse="LCM" />
                <RESULT eventid="44407" points="524" reactiontime="+69" swimtime="00:01:10.52" resultid="47561" heatid="50749" lane="8" entrytime="00:01:20.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="589" reactiontime="+67" swimtime="00:00:26.56" resultid="47562" heatid="50768" lane="5" entrytime="00:00:26.71" entrycourse="LCM" />
                <RESULT eventid="46298" points="634" reactiontime="+67" swimtime="00:00:24.34" resultid="47563" heatid="50822" lane="9" entrytime="00:00:24.86" entrycourse="LCM" />
                <RESULT eventid="46306" points="539" reactiontime="+68" swimtime="00:01:00.82" resultid="47564" heatid="50849" lane="6" entrytime="00:00:59.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Franciszek" lastname="Sobieszek" birthdate="2005-07-07" gender="M" nation="POL" license="106414700129" swrid="4899850" athleteid="47551">
              <RESULTS>
                <RESULT eventid="44378" points="599" reactiontime="+62" swimtime="00:00:55.62" resultid="47552" heatid="50676" lane="1" entrytime="00:00:55.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="588" reactiontime="+56" swimtime="00:01:01.86" resultid="47553" heatid="50723" lane="5" entrytime="00:01:00.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="539" reactiontime="+65" swimtime="00:02:05.30" resultid="47554" heatid="50739" lane="0" entrytime="00:02:03.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.97" />
                    <SPLIT distance="100" swimtime="00:01:00.69" />
                    <SPLIT distance="150" swimtime="00:01:33.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="559" reactiontime="+55" swimtime="00:02:15.86" resultid="47555" heatid="50784" lane="3" entrytime="00:02:12.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                    <SPLIT distance="100" swimtime="00:01:07.04" />
                    <SPLIT distance="150" swimtime="00:01:42.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="568" reactiontime="+67" swimtime="00:04:25.60" resultid="47556" heatid="50799" lane="5" entrytime="00:04:45.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.67" />
                    <SPLIT distance="100" swimtime="00:01:01.98" />
                    <SPLIT distance="150" swimtime="00:01:35.84" />
                    <SPLIT distance="200" swimtime="00:02:10.15" />
                    <SPLIT distance="250" swimtime="00:02:44.17" />
                    <SPLIT distance="300" swimtime="00:03:18.99" />
                    <SPLIT distance="350" swimtime="00:03:53.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46310" points="628" reactiontime="+54" swimtime="00:00:28.02" resultid="47557" heatid="50862" lane="3" entrytime="00:00:27.65" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Bałda" birthdate="2005-03-25" gender="F" nation="POL" license="106414600130" swrid="5088737" athleteid="47571">
              <RESULTS>
                <RESULT eventid="44384" points="663" reactiontime="+72" swimtime="00:00:33.71" resultid="47572" heatid="50703" lane="5" entrytime="00:00:33.59" entrycourse="LCM" />
                <RESULT eventid="44409" points="658" reactiontime="+62" swimtime="00:01:13.73" resultid="47573" heatid="50756" lane="4" entrytime="00:01:13.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="514" reactiontime="+64" swimtime="00:00:30.49" resultid="47574" heatid="50778" lane="4" entrytime="00:00:30.49" entrycourse="LCM" />
                <RESULT eventid="46300" points="538" reactiontime="+74" swimtime="00:00:29.09" resultid="47575" heatid="50830" lane="3" entrytime="00:00:31.57" entrycourse="LCM" />
                <RESULT eventid="46304" points="634" reactiontime="+71" swimtime="00:02:41.93" resultid="47576" heatid="50843" lane="5" entrytime="00:02:42.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                    <SPLIT distance="100" swimtime="00:01:18.02" />
                    <SPLIT distance="150" swimtime="00:02:00.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00515" nation="POL" region="15" clubid="46793" name="KS Posnania Poznań">
          <ATHLETES>
            <ATHLETE firstname="Jan" lastname="Pawlak" birthdate="2005-04-15" gender="M" nation="POL" license="100515700211" swrid="5117073" athleteid="46822">
              <RESULTS>
                <RESULT eventid="44382" points="527" reactiontime="+69" swimtime="00:00:32.11" resultid="46823" heatid="50694" lane="0" entrytime="00:00:34.66" entrycourse="LCM" />
                <RESULT eventid="44407" points="508" reactiontime="+68" swimtime="00:01:11.27" resultid="46824" heatid="50750" lane="5" entrytime="00:01:10.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46302" points="500" reactiontime="+64" swimtime="00:02:38.82" resultid="46825" heatid="50838" lane="4" entrytime="00:02:42.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                    <SPLIT distance="100" swimtime="00:01:16.24" />
                    <SPLIT distance="150" swimtime="00:01:58.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Wielgus" birthdate="2001-03-29" gender="M" nation="POL" license="100515700203" swrid="4905538" athleteid="46835">
              <RESULTS>
                <RESULT eventid="44390" points="516" reactiontime="+64" swimtime="00:02:22.09" resultid="46836" heatid="50710" lane="2" entrytime="00:02:32.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.16" />
                    <SPLIT distance="100" swimtime="00:01:05.91" />
                    <SPLIT distance="150" swimtime="00:01:48.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="464" reactiontime="+64" swimtime="00:00:28.75" resultid="46837" heatid="50760" lane="3" />
                <RESULT eventid="46298" points="505" reactiontime="+65" swimtime="00:00:26.25" resultid="46838" heatid="50819" lane="4" entrytime="00:00:26.31" entrycourse="LCM" />
                <RESULT eventid="46310" points="532" reactiontime="+59" swimtime="00:00:29.61" resultid="46839" heatid="50861" lane="5" entrytime="00:00:30.71" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tymoteusz" lastname="Tomczak" birthdate="2002-05-02" gender="M" nation="POL" license="100515700236" swrid="5071598" athleteid="46826">
              <RESULTS>
                <RESULT eventid="44382" points="622" reactiontime="+69" swimtime="00:00:30.39" resultid="46827" heatid="50695" lane="6" entrytime="00:00:31.77" entrycourse="LCM" />
                <RESULT eventid="46302" points="629" reactiontime="+68" swimtime="00:02:27.19" resultid="46828" heatid="50839" lane="5" entrytime="00:02:26.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                    <SPLIT distance="100" swimtime="00:01:09.61" />
                    <SPLIT distance="150" swimtime="00:01:48.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="458" reactiontime="+65" swimtime="00:02:25.16" resultid="49071" heatid="50780" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                    <SPLIT distance="100" swimtime="00:01:10.21" />
                    <SPLIT distance="150" swimtime="00:01:47.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Apolonia" lastname="Popławska" birthdate="2002-06-01" gender="F" nation="POL" license="100515600277" swrid="4946114" athleteid="46816">
              <RESULTS>
                <RESULT eventid="44380" points="537" reactiontime="+68" swimtime="00:01:03.58" resultid="46817" heatid="50687" lane="0" entrytime="00:01:03.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44384" points="550" reactiontime="+65" swimtime="00:00:35.87" resultid="46818" heatid="50702" lane="2" entrytime="00:00:36.29" entrycourse="LCM" />
                <RESULT eventid="44405" points="506" reactiontime="+55" swimtime="00:02:21.70" resultid="46819" heatid="50741" lane="4" entrytime="00:02:30.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                    <SPLIT distance="100" swimtime="00:01:09.29" />
                    <SPLIT distance="150" swimtime="00:01:46.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="490" reactiontime="+70" swimtime="00:00:30.97" resultid="46820" heatid="50778" lane="2" entrytime="00:00:31.09" entrycourse="LCM" />
                <RESULT eventid="46300" points="552" reactiontime="+66" swimtime="00:00:28.84" resultid="46821" heatid="50834" lane="0" entrytime="00:00:28.69" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kamil" lastname="Cempura" birthdate="2005-04-29" gender="M" nation="POL" license="100515700213" swrid="5117079" athleteid="46803">
              <RESULTS>
                <RESULT eventid="44378" points="424" reactiontime="+68" swimtime="00:01:02.41" resultid="46804" heatid="50672" lane="7" entrytime="00:01:01.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44390" points="399" reactiontime="+65" swimtime="00:02:34.84" resultid="46805" heatid="50710" lane="6" entrytime="00:02:32.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                    <SPLIT distance="100" swimtime="00:01:13.66" />
                    <SPLIT distance="150" swimtime="00:01:58.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="400" reactiontime="+72" swimtime="00:00:28.37" resultid="49072" heatid="50817" lane="6" entrytime="00:00:28.05" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcel" lastname="Wojtyniak" birthdate="2005-06-16" gender="M" nation="POL" license="100515700217" swrid="5117075" athleteid="46794">
              <RESULTS>
                <RESULT eventid="44378" points="497" reactiontime="+66" swimtime="00:00:59.22" resultid="46795" heatid="50668" lane="9" entrytime="00:01:07.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="407" reactiontime="+59" swimtime="00:02:31.01" resultid="46796" heatid="50783" lane="6" entrytime="00:02:39.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                    <SPLIT distance="100" swimtime="00:01:10.87" />
                    <SPLIT distance="150" swimtime="00:01:50.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="478" reactiontime="+67" swimtime="00:00:26.73" resultid="46797" heatid="50819" lane="2" entrytime="00:00:26.46" entrycourse="LCM" />
                <RESULT eventid="46310" points="473" reactiontime="+56" swimtime="00:00:30.79" resultid="46798" heatid="50862" lane="9" entrytime="00:00:30.55" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Zawieja" birthdate="2005-06-25" gender="M" nation="POL" license="100515700218" swrid="5117081" athleteid="46799">
              <RESULTS>
                <RESULT eventid="44378" points="422" reactiontime="+61" swimtime="00:01:02.52" resultid="46800" heatid="50667" lane="6" entrytime="00:01:09.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="395" reactiontime="+62" swimtime="00:02:18.92" resultid="46801" heatid="50733" lane="1" entrytime="00:02:42.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                    <SPLIT distance="100" swimtime="00:01:07.14" />
                    <SPLIT distance="150" swimtime="00:01:43.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="442" reactiontime="+60" swimtime="00:04:48.74" resultid="46802" heatid="50798" lane="2" entrytime="00:05:21.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                    <SPLIT distance="100" swimtime="00:01:07.70" />
                    <SPLIT distance="150" swimtime="00:01:45.05" />
                    <SPLIT distance="200" swimtime="00:02:22.61" />
                    <SPLIT distance="250" swimtime="00:03:00.15" />
                    <SPLIT distance="300" swimtime="00:03:38.19" />
                    <SPLIT distance="350" swimtime="00:04:15.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maksymilian" lastname="Kaczmarek" birthdate="2006-04-17" gender="M" nation="POL" license="100515700239" swrid="5227565" athleteid="46807">
              <RESULTS>
                <RESULT eventid="44378" points="488" reactiontime="+70" swimtime="00:00:59.58" resultid="46808" heatid="50673" lane="1" entrytime="00:01:00.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="480" reactiontime="+70" swimtime="00:02:10.20" resultid="46809" heatid="50736" lane="5" entrytime="00:02:16.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                    <SPLIT distance="100" swimtime="00:01:03.28" />
                    <SPLIT distance="150" swimtime="00:01:37.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="447" reactiontime="+68" swimtime="00:00:27.34" resultid="46810" heatid="50818" lane="8" entrytime="00:00:27.20" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Bocheńska" birthdate="2005-07-22" gender="F" nation="POL" license="100515600255" swrid="5153525" athleteid="46811">
              <RESULTS>
                <RESULT eventid="44380" points="463" reactiontime="+80" swimtime="00:01:06.82" resultid="46812" heatid="50685" lane="1" entrytime="00:01:05.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="309" reactiontime="+78" swimtime="00:00:36.10" resultid="46813" heatid="50776" lane="6" entrytime="00:00:34.12" entrycourse="LCM" />
                <RESULT eventid="46296" points="399" reactiontime="+80" swimtime="00:05:21.13" resultid="46814" heatid="50804" lane="8" entrytime="00:05:36.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.36" />
                    <SPLIT distance="100" swimtime="00:01:13.61" />
                    <SPLIT distance="150" swimtime="00:01:54.37" />
                    <SPLIT distance="200" swimtime="00:02:36.23" />
                    <SPLIT distance="250" swimtime="00:03:18.35" />
                    <SPLIT distance="300" swimtime="00:03:59.95" />
                    <SPLIT distance="350" swimtime="00:04:40.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="448" reactiontime="+77" swimtime="00:00:30.92" resultid="46815" heatid="50831" lane="3" entrytime="00:00:30.44" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olga" lastname="Zarzeczna" birthdate="2005-10-01" gender="F" nation="POL" license="100515600224" swrid="5117085" athleteid="46840">
              <RESULTS>
                <RESULT eventid="44392" points="425" reactiontime="+73" swimtime="00:02:47.64" resultid="46841" heatid="50715" lane="8" entrytime="00:02:43.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                    <SPLIT distance="100" swimtime="00:01:19.91" />
                    <SPLIT distance="150" swimtime="00:02:06.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="278" reactiontime="+73" swimtime="00:00:37.40" resultid="46842" heatid="50776" lane="0" entrytime="00:00:34.99" entrycourse="LCM" />
                <RESULT eventid="46296" points="415" reactiontime="+73" swimtime="00:05:16.86" resultid="46843" heatid="50803" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                    <SPLIT distance="100" swimtime="00:01:13.50" />
                    <SPLIT distance="150" swimtime="00:01:54.25" />
                    <SPLIT distance="200" swimtime="00:02:35.21" />
                    <SPLIT distance="250" swimtime="00:03:15.59" />
                    <SPLIT distance="300" swimtime="00:03:56.34" />
                    <SPLIT distance="350" swimtime="00:04:37.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Wnuk" birthdate="2001-10-29" gender="M" nation="POL" license="100515700150" swrid="4749884" athleteid="46844">
              <RESULTS>
                <RESULT eventid="44394" points="546" reactiontime="+64" swimtime="00:01:03.41" resultid="46845" heatid="50723" lane="0" entrytime="00:01:06.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="509" reactiontime="+68" swimtime="00:02:20.12" resultid="46846" heatid="50784" lane="8" entrytime="00:02:23.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                    <SPLIT distance="100" swimtime="00:01:08.89" />
                    <SPLIT distance="150" swimtime="00:01:45.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46306" points="564" reactiontime="+65" swimtime="00:00:59.90" resultid="46847" heatid="50849" lane="7" entrytime="00:01:00.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46310" points="564" reactiontime="+64" swimtime="00:00:29.04" resultid="46848" heatid="50862" lane="1" entrytime="00:00:29.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patrycja" lastname="Brdęk" birthdate="2005-08-23" gender="F" nation="POL" license="100515600221" swrid="5117086" athleteid="46830">
              <RESULTS>
                <RESULT eventid="44384" points="466" reactiontime="+66" swimtime="00:00:37.92" resultid="46831" heatid="50702" lane="8" entrytime="00:00:37.65" entrycourse="LCM" />
                <RESULT eventid="44409" points="422" reactiontime="+67" swimtime="00:01:25.47" resultid="46832" heatid="50755" lane="0" entrytime="00:01:22.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="354" reactiontime="+68" swimtime="00:00:34.51" resultid="46833" heatid="50777" lane="1" entrytime="00:00:33.24" entrycourse="LCM" />
                <RESULT eventid="46300" points="479" reactiontime="+67" swimtime="00:00:30.25" resultid="46834" heatid="50831" lane="6" entrytime="00:00:30.60" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="95" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="44399" points="587" reactiontime="+62" swimtime="00:04:07.50" resultid="46849" heatid="50730" lane="4" entrytime="00:04:00.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.83" />
                    <SPLIT distance="100" swimtime="00:01:06.04" />
                    <SPLIT distance="150" swimtime="00:01:35.69" />
                    <SPLIT distance="200" swimtime="00:02:11.05" />
                    <SPLIT distance="250" swimtime="00:02:38.36" />
                    <SPLIT distance="300" swimtime="00:03:10.97" />
                    <SPLIT distance="350" swimtime="00:03:37.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="46794" number="1" reactiontime="+62" />
                    <RELAYPOSITION athleteid="46826" number="2" reactiontime="+7" />
                    <RELAYPOSITION athleteid="46844" number="3" reactiontime="+22" />
                    <RELAYPOSITION athleteid="46835" number="4" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46289" points="560" reactiontime="+71" swimtime="00:03:48.35" resultid="46852" heatid="50794" lane="6" entrytime="00:03:47.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.29" />
                    <SPLIT distance="100" swimtime="00:00:57.84" />
                    <SPLIT distance="150" swimtime="00:01:24.99" />
                    <SPLIT distance="200" swimtime="00:01:55.31" />
                    <SPLIT distance="250" swimtime="00:02:22.29" />
                    <SPLIT distance="300" swimtime="00:02:52.46" />
                    <SPLIT distance="350" swimtime="00:03:18.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="46822" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="46844" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="46835" number="3" reactiontime="+29" />
                    <RELAYPOSITION athleteid="46826" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="95" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="44399" points="429" reactiontime="+75" swimtime="00:04:34.72" resultid="46850" heatid="50730" lane="2" entrytime="00:04:32.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                    <SPLIT distance="100" swimtime="00:01:12.24" />
                    <SPLIT distance="150" swimtime="00:01:47.78" />
                    <SPLIT distance="200" swimtime="00:02:28.64" />
                    <SPLIT distance="250" swimtime="00:02:57.88" />
                    <SPLIT distance="300" swimtime="00:03:32.60" />
                    <SPLIT distance="350" swimtime="00:04:01.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="46803" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="46807" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="46822" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="46799" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46289" points="454" reactiontime="+74" swimtime="00:04:04.90" resultid="46853" heatid="50794" lane="7" entrytime="00:03:52.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.56" />
                    <SPLIT distance="100" swimtime="00:00:59.56" />
                    <SPLIT distance="150" swimtime="00:01:29.51" />
                    <SPLIT distance="200" swimtime="00:02:02.67" />
                    <SPLIT distance="250" swimtime="00:02:31.78" />
                    <SPLIT distance="300" swimtime="00:03:03.01" />
                    <SPLIT distance="350" swimtime="00:03:32.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="46807" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="46803" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="46794" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="46799" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="95" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="44401" points="411" reactiontime="+73" swimtime="00:05:09.85" resultid="46851" heatid="50887" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.10" />
                    <SPLIT distance="100" swimtime="00:01:14.65" />
                    <SPLIT distance="150" swimtime="00:01:52.59" />
                    <SPLIT distance="200" swimtime="00:02:39.09" />
                    <SPLIT distance="250" swimtime="00:03:16.71" />
                    <SPLIT distance="300" swimtime="00:04:03.82" />
                    <SPLIT distance="350" swimtime="00:04:33.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="46816" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="46830" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="46840" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="46811" number="4" reactiontime="-7" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46291" points="487" reactiontime="+68" swimtime="00:04:26.92" resultid="46854" heatid="50795" lane="6" entrytime="00:04:19.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                    <SPLIT distance="100" swimtime="00:01:07.68" />
                    <SPLIT distance="150" swimtime="00:01:40.31" />
                    <SPLIT distance="200" swimtime="00:02:16.45" />
                    <SPLIT distance="250" swimtime="00:02:46.83" />
                    <SPLIT distance="300" swimtime="00:03:20.43" />
                    <SPLIT distance="350" swimtime="00:03:51.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="46830" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="46840" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="46816" number="3" reactiontime="+28" />
                    <RELAYPOSITION athleteid="46811" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00601" nation="POL" region="01" clubid="48675" name="WKS Śląsk">
          <ATHLETES>
            <ATHLETE firstname="Adrian" lastname="Worobij" birthdate="2006-03-28" gender="M" nation="POL" license="100601700499" swrid="5223332" athleteid="48692">
              <RESULTS>
                <RESULT eventid="44378" points="527" reactiontime="+66" swimtime="00:00:58.05" resultid="48693" heatid="50675" lane="1" entrytime="00:00:57.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="340" reactiontime="+70" swimtime="00:00:37.17" resultid="48694" heatid="50693" lane="3" entrytime="00:00:37.44" entrycourse="LCM" />
                <RESULT eventid="44403" points="430" reactiontime="+69" swimtime="00:02:15.04" resultid="48695" heatid="50737" lane="8" entrytime="00:02:15.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                    <SPLIT distance="100" swimtime="00:01:06.65" />
                    <SPLIT distance="150" swimtime="00:01:42.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="474" swimtime="00:00:28.56" resultid="48696" heatid="50767" lane="6" entrytime="00:00:28.63" entrycourse="LCM" />
                <RESULT eventid="46294" points="460" reactiontime="+65" swimtime="00:04:44.96" resultid="48697" heatid="50799" lane="2" entrytime="00:04:49.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.29" />
                    <SPLIT distance="100" swimtime="00:01:07.39" />
                    <SPLIT distance="150" swimtime="00:01:44.51" />
                    <SPLIT distance="200" swimtime="00:02:21.60" />
                    <SPLIT distance="250" swimtime="00:02:58.28" />
                    <SPLIT distance="300" swimtime="00:03:35.50" />
                    <SPLIT distance="350" swimtime="00:04:11.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="490" reactiontime="+64" swimtime="00:00:26.51" resultid="48698" heatid="50808" lane="6" />
                <RESULT eventid="46306" points="432" reactiontime="+68" swimtime="00:01:05.48" resultid="48699" heatid="50848" lane="7" entrytime="00:01:07.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maksymilian" lastname="Adamczyk" birthdate="2003-06-02" gender="M" nation="POL" license="100601700376" swrid="5023601" athleteid="48710">
              <RESULTS>
                <RESULT eventid="44378" points="540" reactiontime="+59" swimtime="00:00:57.60" resultid="48711" heatid="50674" lane="2" entrytime="00:00:58.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="528" reactiontime="+51" swimtime="00:01:04.13" resultid="48712" heatid="50723" lane="2" entrytime="00:01:03.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="489" reactiontime="+51" swimtime="00:02:22.00" resultid="48713" heatid="50784" lane="2" entrytime="00:02:15.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                    <SPLIT distance="100" swimtime="00:01:08.99" />
                    <SPLIT distance="150" swimtime="00:01:46.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="507" reactiontime="+59" swimtime="00:00:26.21" resultid="48714" heatid="50820" lane="7" entrytime="00:00:26.14" entrycourse="LCM" />
                <RESULT eventid="46310" points="537" reactiontime="+47" swimtime="00:00:29.52" resultid="48715" heatid="50862" lane="7" entrytime="00:00:29.74" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patryk" lastname="Dąbrowski" birthdate="2000-09-09" gender="M" nation="POL" license="100601700344" swrid="4359249" athleteid="48753">
              <RESULTS>
                <RESULT eventid="44378" points="716" reactiontime="+74" swimtime="00:00:52.42" resultid="48754" heatid="50677" lane="2" entrytime="00:00:52.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="683" reactiontime="+71" swimtime="00:01:55.81" resultid="48755" heatid="50739" lane="5" entrytime="00:01:54.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.14" />
                    <SPLIT distance="100" swimtime="00:00:56.97" />
                    <SPLIT distance="150" swimtime="00:01:26.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="626" reactiontime="+74" swimtime="00:00:26.03" resultid="48756" heatid="50769" lane="7" entrytime="00:00:25.77" entrycourse="LCM" />
                <RESULT eventid="46298" points="659" reactiontime="+70" swimtime="00:00:24.02" resultid="48757" heatid="50822" lane="6" entrytime="00:00:23.90" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Marzec" birthdate="2007-06-24" gender="M" nation="POL" license="100601700557" swrid="5266460" athleteid="48736">
              <RESULTS>
                <RESULT eventid="44378" points="299" reactiontime="+76" swimtime="00:01:10.13" resultid="48737" heatid="50667" lane="2" entrytime="00:01:09.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="278" reactiontime="+66" swimtime="00:01:19.37" resultid="48738" heatid="50720" lane="8" entrytime="00:01:20.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="209" reactiontime="+72" swimtime="00:01:35.70" resultid="48739" heatid="50746" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46310" points="320" reactiontime="+62" swimtime="00:00:35.06" resultid="48740" heatid="50859" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Szeląg" birthdate="2003-03-24" gender="M" nation="POL" license="100601700616" swrid="5105235" athleteid="48758">
              <RESULTS>
                <RESULT eventid="44378" points="607" reactiontime="+68" swimtime="00:00:55.39" resultid="48759" heatid="50676" lane="2" entrytime="00:00:55.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="561" reactiontime="+66" swimtime="00:00:26.99" resultid="48760" heatid="50768" lane="8" entrytime="00:00:27.55" entrycourse="LCM" />
                <RESULT eventid="46298" points="513" reactiontime="+66" swimtime="00:00:26.11" resultid="48761" heatid="50821" lane="0" entrytime="00:00:25.76" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Goczling" birthdate="2008-02-19" gender="M" nation="POL" license="100601700588" swrid="5266500" athleteid="48775">
              <RESULTS>
                <RESULT eventid="44382" points="313" reactiontime="+51" swimtime="00:00:38.20" resultid="48776" heatid="50692" lane="4" entrytime="00:00:44.01" entrycourse="LCM" />
                <RESULT eventid="44407" points="283" reactiontime="+68" swimtime="00:01:26.55" resultid="48777" heatid="50747" lane="3" entrytime="00:01:31.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="283" swimtime="00:00:33.91" resultid="48778" heatid="50762" lane="4" entrytime="00:00:35.44" entrycourse="LCM" />
                <RESULT eventid="46306" points="235" reactiontime="+53" swimtime="00:01:20.20" resultid="48779" heatid="50845" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Bieroński" birthdate="1999-03-23" gender="M" nation="POL" license="100601700350" swrid="4639547" athleteid="48676">
              <RESULTS>
                <RESULT eventid="44378" points="692" reactiontime="+72" swimtime="00:00:53.02" resultid="48677" heatid="50677" lane="6" entrytime="00:00:52.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="673" reactiontime="+74" swimtime="00:01:56.35" resultid="48678" heatid="50739" lane="3" entrytime="00:01:57.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.32" />
                    <SPLIT distance="100" swimtime="00:00:56.94" />
                    <SPLIT distance="150" swimtime="00:01:27.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="632" reactiontime="+71" swimtime="00:00:25.95" resultid="48679" heatid="50769" lane="3" entrytime="00:00:25.37" entrycourse="LCM" />
                <RESULT eventid="46298" points="688" reactiontime="+72" swimtime="00:00:23.68" resultid="48680" heatid="50822" lane="3" entrytime="00:00:23.46" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Bednarczyk" birthdate="1994-01-06" gender="M" nation="POL" license="500601700657" swrid="4114570" athleteid="48746">
              <RESULTS>
                <RESULT eventid="44378" points="530" reactiontime="+70" swimtime="00:00:57.93" resultid="48747" heatid="50663" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44390" status="DNS" swimtime="00:00:00.00" resultid="48748" heatid="50708" lane="6" />
                <RESULT eventid="44403" points="418" reactiontime="+79" swimtime="00:02:16.36" resultid="48749" heatid="50732" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.85" />
                    <SPLIT distance="100" swimtime="00:01:03.85" />
                    <SPLIT distance="150" swimtime="00:01:39.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="577" reactiontime="+72" swimtime="00:00:26.75" resultid="48750" heatid="50761" lane="1" />
                <RESULT eventid="46298" points="541" reactiontime="+72" swimtime="00:00:25.65" resultid="48751" heatid="50808" lane="0" />
                <RESULT eventid="46306" points="500" reactiontime="+73" swimtime="00:01:02.33" resultid="48752" heatid="50845" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Szarek" birthdate="2006-06-27" gender="M" nation="POL" license="100601700498" swrid="5166099" athleteid="48681">
              <RESULTS>
                <RESULT eventid="44378" points="565" reactiontime="+77" swimtime="00:00:56.72" resultid="48682" heatid="50675" lane="6" entrytime="00:00:56.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="466" reactiontime="+75" swimtime="00:00:33.47" resultid="48683" heatid="50694" lane="6" entrytime="00:00:33.20" entrycourse="LCM" />
                <RESULT eventid="44390" points="480" reactiontime="+77" swimtime="00:02:25.51" resultid="48684" heatid="50711" lane="7" entrytime="00:02:24.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                    <SPLIT distance="100" swimtime="00:01:10.15" />
                    <SPLIT distance="150" swimtime="00:01:52.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="509" reactiontime="+73" swimtime="00:02:07.69" resultid="48685" heatid="50738" lane="6" entrytime="00:02:05.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.25" />
                    <SPLIT distance="100" swimtime="00:01:01.72" />
                    <SPLIT distance="150" swimtime="00:01:35.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="371" reactiontime="+71" swimtime="00:01:19.11" resultid="48686" heatid="50749" lane="3" entrytime="00:01:16.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="414" reactiontime="+75" swimtime="00:00:29.87" resultid="48687" heatid="50759" lane="7" />
                <RESULT eventid="46294" points="552" reactiontime="+66" swimtime="00:04:28.12" resultid="48688" heatid="50800" lane="9" entrytime="00:04:37.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.88" />
                    <SPLIT distance="100" swimtime="00:01:03.91" />
                    <SPLIT distance="150" swimtime="00:01:38.53" />
                    <SPLIT distance="200" swimtime="00:02:13.76" />
                    <SPLIT distance="250" swimtime="00:02:48.73" />
                    <SPLIT distance="300" swimtime="00:03:23.79" />
                    <SPLIT distance="350" swimtime="00:03:57.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="460" reactiontime="+75" swimtime="00:00:27.07" resultid="48689" heatid="50807" lane="3" />
                <RESULT eventid="46302" points="419" reactiontime="+68" swimtime="00:02:48.46" resultid="48690" heatid="50838" lane="5" entrytime="00:02:45.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.03" />
                    <SPLIT distance="100" swimtime="00:01:22.43" />
                    <SPLIT distance="150" swimtime="00:02:06.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46306" points="387" reactiontime="+68" swimtime="00:01:07.90" resultid="48691" heatid="50848" lane="2" entrytime="00:01:06.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maksymilian" lastname="Sypko" birthdate="2005-06-05" gender="M" nation="POL" license="100601700445" swrid="5198189" athleteid="49070">
              <RESULTS>
                <RESULT eventid="44407" points="467" reactiontime="+71" swimtime="00:01:13.29" resultid="49197" heatid="50749" lane="1" entrytime="00:01:18.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44378" points="511" reactiontime="+72" swimtime="00:00:58.65" resultid="49198" heatid="50674" lane="0" entrytime="00:00:58.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44390" points="504" reactiontime="+72" swimtime="00:02:23.16" resultid="49199" heatid="50711" lane="2" entrytime="00:02:24.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.21" />
                    <SPLIT distance="100" swimtime="00:01:07.81" />
                    <SPLIT distance="150" swimtime="00:01:50.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="471" reactiontime="+68" swimtime="00:04:42.72" resultid="49200" heatid="50800" lane="8" entrytime="00:04:36.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.56" />
                    <SPLIT distance="100" swimtime="00:01:01.83" />
                    <SPLIT distance="150" swimtime="00:01:36.88" />
                    <SPLIT distance="200" swimtime="00:02:12.35" />
                    <SPLIT distance="250" swimtime="00:02:47.94" />
                    <SPLIT distance="300" swimtime="00:03:24.81" />
                    <SPLIT distance="350" swimtime="00:04:03.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Cyrek" birthdate="2007-02-21" gender="M" nation="POL" license="100601700563" swrid="5226962" athleteid="48726">
              <RESULTS>
                <RESULT eventid="44378" points="445" reactiontime="+73" swimtime="00:01:01.42" resultid="48727" heatid="50671" lane="8" entrytime="00:01:03.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="407" reactiontime="+78" swimtime="00:00:30.04" resultid="48728" heatid="50758" lane="3" />
                <RESULT eventid="46298" points="422" reactiontime="+75" swimtime="00:00:27.86" resultid="48729" heatid="50808" lane="3" />
                <RESULT eventid="46310" points="420" reactiontime="+66" swimtime="00:00:32.03" resultid="48730" heatid="50858" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hanna" lastname="Prętkowska" birthdate="2007-08-17" gender="F" nation="POL" license="100601600564" swrid="5354932" athleteid="48810">
              <RESULTS>
                <RESULT eventid="44384" points="171" swimtime="00:00:52.93" resultid="48811" heatid="50699" lane="0" />
                <RESULT eventid="44396" points="303" reactiontime="+87" swimtime="00:01:25.65" resultid="48812" heatid="50725" lane="3" entrytime="00:01:25.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44409" points="192" reactiontime="+77" swimtime="00:01:51.03" resultid="48813" heatid="50753" lane="1" entrytime="00:01:38.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="301" reactiontime="+77" swimtime="00:00:40.23" resultid="48814" heatid="50904" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Kiszczak" birthdate="2000-04-23" gender="M" nation="POL" license="100601700467" swrid="4705231" athleteid="48722">
              <RESULTS>
                <RESULT eventid="44378" status="DNS" swimtime="00:00:00.00" resultid="48723" heatid="50677" lane="3" entrytime="00:00:51.09" entrycourse="LCM" />
                <RESULT eventid="44411" status="DNS" swimtime="00:00:00.00" resultid="48724" heatid="50769" lane="5" entrytime="00:00:25.04" entrycourse="LCM" />
                <RESULT eventid="46310" status="DNS" swimtime="00:00:00.00" resultid="48725" heatid="50862" lane="4" entrytime="00:00:26.55" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Konrad" lastname="Powroźnik" birthdate="1997-05-30" gender="M" nation="POL" license="100601700513" swrid="4369083" athleteid="48820">
              <RESULTS>
                <RESULT eventid="44386" points="628" reactiontime="+82" swimtime="00:02:09.27" resultid="48821" heatid="50705" lane="5" entrytime="00:02:08.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.38" />
                    <SPLIT distance="100" swimtime="00:01:00.67" />
                    <SPLIT distance="150" swimtime="00:01:34.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44390" points="599" reactiontime="+72" swimtime="00:02:15.17" resultid="48822" heatid="50711" lane="4" entrytime="00:02:08.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.41" />
                    <SPLIT distance="100" swimtime="00:01:04.48" />
                    <SPLIT distance="150" swimtime="00:01:43.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Dudek" birthdate="2008-01-07" gender="M" nation="POL" license="100601700653" swrid="4989146" athleteid="48770">
              <RESULTS>
                <RESULT eventid="44382" points="209" reactiontime="+72" swimtime="00:00:43.72" resultid="48771" heatid="50692" lane="8" />
                <RESULT eventid="44411" points="288" reactiontime="+68" swimtime="00:00:33.70" resultid="48772" heatid="50759" lane="4" />
                <RESULT eventid="46298" points="297" reactiontime="+80" swimtime="00:00:31.31" resultid="48773" heatid="50807" lane="0" />
                <RESULT eventid="46310" points="221" reactiontime="+79" swimtime="00:00:39.67" resultid="48774" heatid="50856" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Dziemieszkiewicz" birthdate="2008-03-18" gender="M" nation="POL" license="100601700654" swrid="4989150" athleteid="48731">
              <RESULTS>
                <RESULT eventid="44378" status="DNS" swimtime="00:00:00.00" resultid="48732" heatid="50667" lane="4" entrytime="00:01:07.88" entrycourse="LCM" />
                <RESULT eventid="44382" status="DNS" swimtime="00:00:00.00" resultid="48733" heatid="50689" lane="5" />
                <RESULT eventid="44403" status="DNS" swimtime="00:00:00.00" resultid="48734" heatid="50734" lane="0" entrytime="00:02:32.69" entrycourse="LCM" />
                <RESULT eventid="46298" status="DNS" swimtime="00:00:00.00" resultid="48735" heatid="50810" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maksymilian" lastname="Pruszyński" birthdate="2007-03-28" gender="M" nation="POL" license="100601700559" swrid="5266447" athleteid="48842">
              <RESULTS>
                <RESULT eventid="44394" status="DNS" swimtime="00:00:00.00" resultid="48843" heatid="50718" lane="5" />
                <RESULT eventid="44411" status="DNS" swimtime="00:00:00.00" resultid="48844" heatid="50759" lane="5" />
                <RESULT eventid="46298" status="DNS" swimtime="00:00:00.00" resultid="48845" heatid="50809" lane="4" />
                <RESULT eventid="46310" status="DNS" swimtime="00:00:00.00" resultid="48846" heatid="50855" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Poręba" birthdate="2007-01-11" gender="M" nation="POL" license="100601700528" swrid="5266480" athleteid="48741">
              <RESULTS>
                <RESULT eventid="44378" points="426" reactiontime="+70" swimtime="00:01:02.32" resultid="48742" heatid="50672" lane="2" entrytime="00:01:01.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="451" reactiontime="+71" swimtime="00:00:29.03" resultid="48743" heatid="50765" lane="5" entrytime="00:00:30.19" entrycourse="LCM" />
                <RESULT eventid="46298" points="452" reactiontime="+72" swimtime="00:00:27.23" resultid="48744" heatid="50812" lane="2" entrytime="00:00:36.38" entrycourse="LCM" />
                <RESULT eventid="46306" points="411" reactiontime="+74" swimtime="00:01:06.53" resultid="48745" heatid="50848" lane="0" entrytime="00:01:08.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Weronika" lastname="Fursewicz" birthdate="2007-08-04" gender="F" nation="POL" license="100601600556" swrid="5266456" athleteid="48800">
              <RESULTS>
                <RESULT eventid="44384" points="308" reactiontime="+64" swimtime="00:00:43.52" resultid="48801" heatid="50697" lane="6" />
                <RESULT eventid="44396" points="314" reactiontime="+71" swimtime="00:01:24.62" resultid="48802" heatid="50725" lane="2" entrytime="00:01:25.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44409" points="296" reactiontime="+49" swimtime="00:01:36.16" resultid="48803" heatid="50752" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" status="DNS" swimtime="00:00:00.00" resultid="48804" heatid="50903" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Ostaszewski" birthdate="2007-12-17" gender="M" nation="POL" license="100601700527" swrid="4005351" athleteid="48837">
              <RESULTS>
                <RESULT eventid="44394" points="364" reactiontime="+73" swimtime="00:01:12.56" resultid="48838" heatid="50721" lane="0" entrytime="00:01:15.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="339" reactiontime="+70" swimtime="00:02:40.48" resultid="48839" heatid="50781" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.09" />
                    <SPLIT distance="100" swimtime="00:01:19.27" />
                    <SPLIT distance="150" swimtime="00:02:00.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="375" reactiontime="+64" swimtime="00:05:04.99" resultid="48840" heatid="50796" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                    <SPLIT distance="100" swimtime="00:01:09.86" />
                    <SPLIT distance="150" swimtime="00:01:48.51" />
                    <SPLIT distance="200" swimtime="00:02:27.77" />
                    <SPLIT distance="250" swimtime="00:03:08.01" />
                    <SPLIT distance="300" swimtime="00:03:48.14" />
                    <SPLIT distance="350" swimtime="00:04:27.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46310" points="353" reactiontime="+69" swimtime="00:00:33.93" resultid="48841" heatid="50856" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Kozdrowski" birthdate="2007-01-28" gender="M" nation="POL" license="100601700589" swrid="5341438" athleteid="48785">
              <RESULTS>
                <RESULT eventid="44382" points="212" reactiontime="+50" swimtime="00:00:43.48" resultid="48786" heatid="50691" lane="2" />
                <RESULT eventid="44390" points="279" reactiontime="+71" swimtime="00:02:54.44" resultid="48787" heatid="50709" lane="8" entrytime="00:02:50.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.06" />
                    <SPLIT distance="100" swimtime="00:01:23.11" />
                    <SPLIT distance="150" swimtime="00:02:15.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="207" reactiontime="+69" swimtime="00:01:36.13" resultid="48788" heatid="50747" lane="7" entrytime="00:01:38.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46306" points="210" reactiontime="+47" swimtime="00:01:23.19" resultid="48789" heatid="50846" lane="0" entrytime="00:01:21.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Matysiak" birthdate="2007-07-21" gender="M" nation="POL" license="100601700524" swrid="5266498" athleteid="48790">
              <RESULTS>
                <RESULT eventid="44382" points="272" reactiontime="+68" swimtime="00:00:40.04" resultid="48791" heatid="50692" lane="7" />
                <RESULT eventid="44390" points="326" reactiontime="+65" swimtime="00:02:45.58" resultid="48792" heatid="50709" lane="6" entrytime="00:02:46.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                    <SPLIT distance="100" swimtime="00:01:20.07" />
                    <SPLIT distance="150" swimtime="00:02:08.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="279" reactiontime="+55" swimtime="00:01:26.99" resultid="48793" heatid="50747" lane="4" entrytime="00:01:30.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46302" points="297" reactiontime="+67" swimtime="00:03:08.97" resultid="48794" heatid="50838" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.12" />
                    <SPLIT distance="100" swimtime="00:01:31.92" />
                    <SPLIT distance="150" swimtime="00:02:20.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Radzikowski" birthdate="2008-04-17" gender="M" nation="POL" license="100601700529" swrid="5166095" athleteid="48795">
              <RESULTS>
                <RESULT eventid="44382" points="402" reactiontime="+59" swimtime="00:00:35.15" resultid="48796" heatid="50691" lane="0" />
                <RESULT eventid="44390" points="433" reactiontime="+63" swimtime="00:02:30.62" resultid="48797" heatid="50710" lane="5" entrytime="00:02:28.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.49" />
                    <SPLIT distance="100" swimtime="00:01:12.56" />
                    <SPLIT distance="150" swimtime="00:01:56.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="417" reactiontime="+64" swimtime="00:01:16.11" resultid="48798" heatid="50749" lane="2" entrytime="00:01:18.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46302" points="454" reactiontime="+64" swimtime="00:02:44.07" resultid="48799" heatid="50837" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                    <SPLIT distance="100" swimtime="00:01:19.68" />
                    <SPLIT distance="150" swimtime="00:02:02.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mikołaj" lastname="Kopacz" birthdate="2007-10-22" gender="M" nation="POL" license="100601700621" swrid="4978571" athleteid="48780">
              <RESULTS>
                <RESULT eventid="44382" points="257" reactiontime="+75" swimtime="00:00:40.77" resultid="48781" heatid="50689" lane="3" />
                <RESULT eventid="44411" points="209" reactiontime="+79" swimtime="00:00:37.51" resultid="48782" heatid="50758" lane="6" />
                <RESULT eventid="46298" points="279" reactiontime="+71" swimtime="00:00:31.99" resultid="48783" heatid="50809" lane="5" />
                <RESULT eventid="46310" points="206" reactiontime="+71" swimtime="00:00:40.60" resultid="48784" heatid="50857" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Turbańska" birthdate="2007-08-03" gender="F" nation="POL" license="100601600554" swrid="5266449" athleteid="48815">
              <RESULTS>
                <RESULT eventid="44384" points="539" reactiontime="+77" swimtime="00:00:36.12" resultid="48816" heatid="50699" lane="7" />
                <RESULT eventid="44392" points="375" reactiontime="+78" swimtime="00:02:54.81" resultid="48817" heatid="50713" lane="4" entrytime="00:02:56.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.16" />
                    <SPLIT distance="100" swimtime="00:01:23.37" />
                    <SPLIT distance="150" swimtime="00:02:13.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44409" points="464" reactiontime="+82" swimtime="00:01:22.78" resultid="48818" heatid="50754" lane="7" entrytime="00:01:27.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46304" points="301" reactiontime="+57" swimtime="00:03:27.41" resultid="48819" heatid="50840" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.09" />
                    <SPLIT distance="100" swimtime="00:01:38.84" />
                    <SPLIT distance="150" swimtime="00:02:33.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Pluta" birthdate="2007-04-05" gender="F" nation="POL" license="100601600647" swrid="5266494" athleteid="48847">
              <RESULTS>
                <RESULT eventid="44396" points="440" reactiontime="+84" swimtime="00:01:15.69" resultid="48848" heatid="50727" lane="2" entrytime="00:01:15.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="411" reactiontime="+58" swimtime="00:00:32.84" resultid="48849" heatid="50770" lane="4" />
                <RESULT eventid="44417" points="418" reactiontime="+80" swimtime="00:02:44.90" resultid="48850" heatid="50787" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.38" />
                    <SPLIT distance="100" swimtime="00:01:22.14" />
                    <SPLIT distance="150" swimtime="00:02:04.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46308" points="332" reactiontime="+57" swimtime="00:01:20.09" resultid="48851" heatid="50899" lane="4" entrytime="00:01:17.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martyna" lastname="Napieralczyk" birthdate="2008-06-16" gender="F" nation="POL" license="100601600525" swrid="5266472" athleteid="48832">
              <RESULTS>
                <RESULT eventid="44392" points="412" reactiontime="+79" swimtime="00:02:49.49" resultid="48833" heatid="50714" lane="3" entrytime="00:02:50.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.87" />
                    <SPLIT distance="100" swimtime="00:01:18.75" />
                    <SPLIT distance="150" swimtime="00:02:10.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44417" points="428" reactiontime="+62" swimtime="00:02:43.63" resultid="48834" heatid="50787" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.40" />
                    <SPLIT distance="100" swimtime="00:01:21.22" />
                    <SPLIT distance="150" swimtime="00:02:02.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="408" reactiontime="+55" swimtime="00:05:18.58" resultid="48835" heatid="50801" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                    <SPLIT distance="100" swimtime="00:01:13.92" />
                    <SPLIT distance="150" swimtime="00:01:53.88" />
                    <SPLIT distance="200" swimtime="00:02:34.88" />
                    <SPLIT distance="250" swimtime="00:03:16.58" />
                    <SPLIT distance="300" swimtime="00:03:58.52" />
                    <SPLIT distance="350" swimtime="00:04:39.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="414" reactiontime="+57" swimtime="00:00:36.19" resultid="48836" heatid="50907" lane="0" entrytime="00:00:37.30" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Modlińska" birthdate="2005-06-30" gender="F" nation="POL" license="100601600650" swrid="5147673" athleteid="48762">
              <RESULTS>
                <RESULT eventid="44380" points="527" reactiontime="+70" swimtime="00:01:03.99" resultid="48763" heatid="50686" lane="3" entrytime="00:01:04.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="455" reactiontime="+73" swimtime="00:00:31.75" resultid="48764" heatid="50778" lane="5" entrytime="00:00:30.69" entrycourse="LCM" />
                <RESULT eventid="46300" points="533" reactiontime="+66" swimtime="00:00:29.18" resultid="48765" heatid="50833" lane="4" entrytime="00:00:28.90" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Gałecki" birthdate="2006-01-03" gender="M" nation="POL" license="100601700553" swrid="5334389" athleteid="48700">
              <RESULTS>
                <RESULT eventid="44378" points="478" reactiontime="+72" swimtime="00:00:59.98" resultid="48701" heatid="50673" lane="7" entrytime="00:01:00.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="403" reactiontime="+74" swimtime="00:01:10.17" resultid="48702" heatid="50717" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="452" reactiontime="+73" swimtime="00:02:12.86" resultid="48703" heatid="50737" lane="3" entrytime="00:02:11.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                    <SPLIT distance="100" swimtime="00:01:06.09" />
                    <SPLIT distance="150" swimtime="00:01:40.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="423" reactiontime="+68" swimtime="00:00:29.66" resultid="48704" heatid="50759" lane="6" />
                <RESULT eventid="44415" points="422" reactiontime="+74" swimtime="00:02:29.16" resultid="48705" heatid="50782" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.37" />
                    <SPLIT distance="100" swimtime="00:01:13.61" />
                    <SPLIT distance="150" swimtime="00:01:51.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="445" reactiontime="+73" swimtime="00:04:48.24" resultid="48706" heatid="50797" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                    <SPLIT distance="100" swimtime="00:01:08.88" />
                    <SPLIT distance="150" swimtime="00:01:46.16" />
                    <SPLIT distance="200" swimtime="00:02:24.08" />
                    <SPLIT distance="250" swimtime="00:03:02.03" />
                    <SPLIT distance="300" swimtime="00:03:39.69" />
                    <SPLIT distance="350" swimtime="00:04:15.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="431" reactiontime="+73" swimtime="00:00:27.67" resultid="48707" heatid="50809" lane="7" />
                <RESULT eventid="46306" points="401" reactiontime="+73" swimtime="00:01:07.12" resultid="48708" heatid="50848" lane="1" entrytime="00:01:07.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46310" points="414" reactiontime="+70" swimtime="00:00:32.18" resultid="48709" heatid="50856" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwia" lastname="Grzesiak" birthdate="2007-11-16" gender="F" nation="POL" license="100601600530" swrid="5436179" athleteid="48827">
              <RESULTS>
                <RESULT eventid="44388" points="449" reactiontime="+73" swimtime="00:02:39.06" resultid="48828" heatid="50706" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.67" />
                    <SPLIT distance="100" swimtime="00:01:14.15" />
                    <SPLIT distance="150" swimtime="00:01:56.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="519" reactiontime="+73" swimtime="00:02:20.53" resultid="48829" heatid="50743" lane="1" entrytime="00:02:19.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                    <SPLIT distance="100" swimtime="00:01:08.27" />
                    <SPLIT distance="150" swimtime="00:01:45.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="433" reactiontime="+74" swimtime="00:00:32.29" resultid="48830" heatid="50771" lane="3" />
                <RESULT eventid="46308" points="500" reactiontime="+71" swimtime="00:01:09.89" resultid="48831" heatid="50901" lane="1" entrytime="00:01:08.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Szwedzki" birthdate="1994-04-18" gender="M" nation="POL" license="100601700371" swrid="4181303" athleteid="48823">
              <RESULTS>
                <RESULT eventid="44386" points="729" reactiontime="+69" swimtime="00:02:02.99" resultid="48824" heatid="50705" lane="4" entrytime="00:02:06.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.13" />
                    <SPLIT distance="100" swimtime="00:00:58.42" />
                    <SPLIT distance="150" swimtime="00:01:30.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="697" reactiontime="+60" swimtime="00:02:06.17" resultid="48826" heatid="50784" lane="4" entrytime="00:02:03.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                    <SPLIT distance="100" swimtime="00:01:02.08" />
                    <SPLIT distance="150" swimtime="00:01:34.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46302" points="784" reactiontime="+70" swimtime="00:02:16.74" resultid="49892" heatid="50839" lane="4" entrytime="00:02:08.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.03" />
                    <SPLIT distance="100" swimtime="00:01:05.97" />
                    <SPLIT distance="150" swimtime="00:01:41.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="44399" points="347" reactiontime="+70" swimtime="00:04:54.84" resultid="48852" heatid="50730" lane="9" entrytime="00:04:55.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                    <SPLIT distance="100" swimtime="00:01:13.91" />
                    <SPLIT distance="150" swimtime="00:01:54.08" />
                    <SPLIT distance="200" swimtime="00:02:42.13" />
                    <SPLIT distance="250" swimtime="00:03:13.41" />
                    <SPLIT distance="300" swimtime="00:03:50.33" />
                    <SPLIT distance="350" swimtime="00:04:20.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="48726" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="48790" number="2" reactiontime="+3" />
                    <RELAYPOSITION athleteid="48741" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="48837" number="4" reactiontime="+17" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46289" points="387" reactiontime="+78" swimtime="00:04:18.26" resultid="48854" heatid="50793" lane="4" entrytime="00:04:13.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                    <SPLIT distance="100" swimtime="00:01:01.39" />
                    <SPLIT distance="150" swimtime="00:01:34.21" />
                    <SPLIT distance="200" swimtime="00:02:11.32" />
                    <SPLIT distance="250" swimtime="00:02:41.42" />
                    <SPLIT distance="300" swimtime="00:03:15.86" />
                    <SPLIT distance="350" swimtime="00:03:44.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="48726" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="48785" number="2" />
                    <RELAYPOSITION athleteid="48837" number="3" />
                    <RELAYPOSITION athleteid="48741" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46314" points="360" reactiontime="+67" swimtime="00:09:47.84" resultid="48856" heatid="50870" lane="6" entrytime="00:09:43.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.73" />
                    <SPLIT distance="100" swimtime="00:01:12.80" />
                    <SPLIT distance="150" swimtime="00:01:51.77" />
                    <SPLIT distance="200" swimtime="00:02:28.46" />
                    <SPLIT distance="250" swimtime="00:02:59.94" />
                    <SPLIT distance="300" swimtime="00:03:36.35" />
                    <SPLIT distance="350" swimtime="00:04:14.28" />
                    <SPLIT distance="400" swimtime="00:04:51.52" />
                    <SPLIT distance="450" swimtime="00:05:25.16" />
                    <SPLIT distance="500" swimtime="00:06:05.72" />
                    <SPLIT distance="550" swimtime="00:06:46.37" />
                    <SPLIT distance="600" swimtime="00:07:26.18" />
                    <SPLIT distance="650" swimtime="00:07:57.37" />
                    <SPLIT distance="700" swimtime="00:08:35.27" />
                    <SPLIT distance="750" swimtime="00:09:13.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="48785" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="48837" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="48790" number="3" reactiontime="+28" />
                    <RELAYPOSITION athleteid="48741" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="44401" points="364" reactiontime="+70" swimtime="00:05:22.41" resultid="48853" heatid="50731" lane="6" entrytime="00:04:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                    <SPLIT distance="100" swimtime="00:01:18.57" />
                    <SPLIT distance="150" swimtime="00:01:57.11" />
                    <SPLIT distance="200" swimtime="00:02:43.54" />
                    <SPLIT distance="250" swimtime="00:03:20.10" />
                    <SPLIT distance="300" swimtime="00:04:06.24" />
                    <SPLIT distance="350" swimtime="00:04:43.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="48815" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="48827" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="48847" number="4" reactiontime="+7" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46291" points="409" reactiontime="+69" swimtime="00:04:42.96" resultid="48855" heatid="50795" lane="7" entrytime="00:04:24.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.22" />
                    <SPLIT distance="100" swimtime="00:01:08.83" />
                    <SPLIT distance="150" swimtime="00:01:45.93" />
                    <SPLIT distance="200" swimtime="00:02:28.26" />
                    <SPLIT distance="250" swimtime="00:03:01.09" />
                    <SPLIT distance="300" swimtime="00:03:39.26" />
                    <SPLIT distance="350" swimtime="00:04:09.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="48847" number="1" reactiontime="+69" />
                    <RELAYPOSITION number="2" reactiontime="+19" />
                    <RELAYPOSITION athleteid="48815" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="48827" number="4" reactiontime="-8" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46316" points="359" reactiontime="+57" swimtime="00:10:48.84" resultid="48857" heatid="50871" lane="6" entrytime="00:10:08.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                    <SPLIT distance="100" swimtime="00:01:11.57" />
                    <SPLIT distance="150" swimtime="00:01:50.85" />
                    <SPLIT distance="200" swimtime="00:02:30.02" />
                    <SPLIT distance="250" swimtime="00:03:10.48" />
                    <SPLIT distance="300" swimtime="00:03:55.94" />
                    <SPLIT distance="350" swimtime="00:04:40.67" />
                    <SPLIT distance="400" swimtime="00:05:25.12" />
                    <SPLIT distance="450" swimtime="00:06:06.13" />
                    <SPLIT distance="500" swimtime="00:06:51.02" />
                    <SPLIT distance="550" swimtime="00:07:35.80" />
                    <SPLIT distance="600" swimtime="00:08:19.44" />
                    <SPLIT distance="650" swimtime="00:08:52.35" />
                    <SPLIT distance="700" swimtime="00:09:30.02" />
                    <SPLIT distance="750" swimtime="00:10:09.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="48847" number="1" reactiontime="+57" />
                    <RELAYPOSITION number="2" reactiontime="+12" />
                    <RELAYPOSITION athleteid="48815" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="48827" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="04001" nation="POL" region="01" clubid="46517" name="KS &quot;BALTI&quot; Bielawa">
          <ATHLETES>
            <ATHLETE firstname="Adrian" lastname="Zarzycki" birthdate="2006-05-13" gender="M" nation="POL" license="104001700003" swrid="5024249" athleteid="46518">
              <RESULTS>
                <RESULT eventid="44378" points="483" reactiontime="+68" swimtime="00:00:59.77" resultid="46519" heatid="50672" lane="9" entrytime="00:01:02.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="428" reactiontime="+72" swimtime="00:00:34.41" resultid="46520" heatid="50694" lane="8" entrytime="00:00:34.52" entrycourse="LCM" />
                <RESULT eventid="44411" points="423" reactiontime="+71" swimtime="00:00:29.66" resultid="46521" heatid="50759" lane="8" />
                <RESULT eventid="46298" points="456" reactiontime="+72" swimtime="00:00:27.16" resultid="46522" heatid="50817" lane="3" entrytime="00:00:27.90" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Kuleta" birthdate="2006-01-19" gender="F" nation="POL" license="104001600001" swrid="5024246" athleteid="46536">
              <RESULTS>
                <RESULT eventid="44413" points="452" reactiontime="+69" swimtime="00:00:31.82" resultid="46537" heatid="50778" lane="9" entrytime="00:00:32.12" entrycourse="LCM" />
                <RESULT eventid="46300" points="527" reactiontime="+51" swimtime="00:00:29.30" resultid="46538" heatid="50823" lane="4" />
                <RESULT eventid="46312" points="521" reactiontime="+62" swimtime="00:00:33.52" resultid="46539" heatid="50908" lane="6" entrytime="00:00:33.77" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olivier" lastname="Paprzycki" birthdate="2006-11-10" gender="M" nation="POL" license="104001700010" swrid="5186697" athleteid="46523">
              <RESULTS>
                <RESULT eventid="44378" points="407" reactiontime="+74" swimtime="00:01:03.28" resultid="46524" heatid="50663" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44386" points="236" reactiontime="+78" swimtime="00:02:59.16" resultid="46525" heatid="50705" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                    <SPLIT distance="100" swimtime="00:01:16.56" />
                    <SPLIT distance="150" swimtime="00:02:05.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="399" reactiontime="+75" swimtime="00:00:30.23" resultid="46526" heatid="50765" lane="2" entrytime="00:00:30.42" entrycourse="LCM" />
                <RESULT eventid="46298" points="426" reactiontime="+71" swimtime="00:00:27.78" resultid="46527" heatid="50817" lane="8" entrytime="00:00:28.37" entrycourse="LCM" />
                <RESULT eventid="46306" points="298" reactiontime="+73" swimtime="00:01:14.05" resultid="46528" heatid="50847" lane="9" entrytime="00:01:13.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Pliszka" birthdate="2006-05-16" gender="M" nation="POL" license="104001700007" swrid="5043178" athleteid="46529">
              <RESULTS>
                <RESULT eventid="44378" points="538" reactiontime="+69" swimtime="00:00:57.65" resultid="46530" heatid="50674" lane="5" entrytime="00:00:58.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44390" points="473" reactiontime="+68" swimtime="00:02:26.30" resultid="46531" heatid="50711" lane="9" entrytime="00:02:27.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.54" />
                    <SPLIT distance="100" swimtime="00:01:09.04" />
                    <SPLIT distance="150" swimtime="00:01:53.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="490" reactiontime="+70" swimtime="00:02:09.35" resultid="46532" heatid="50738" lane="9" entrytime="00:02:10.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.77" />
                    <SPLIT distance="100" swimtime="00:01:02.08" />
                    <SPLIT distance="150" swimtime="00:01:36.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="460" reactiontime="+71" swimtime="00:00:28.84" resultid="46533" heatid="50765" lane="4" entrytime="00:00:30.17" entrycourse="LCM" />
                <RESULT eventid="46298" points="487" reactiontime="+77" swimtime="00:00:26.56" resultid="46534" heatid="50818" lane="0" entrytime="00:00:27.31" entrycourse="LCM" />
                <RESULT eventid="46306" points="434" reactiontime="+71" swimtime="00:01:05.33" resultid="46535" heatid="50845" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02401" nation="POL" region="01" clubid="47018" name="MKP ,,Atol&apos;&apos; Oleśnica">
          <ATHLETES>
            <ATHLETE firstname="Wiktor" lastname="Korzeniowski" birthdate="2003-11-04" gender="M" nation="POL" license="102401700076" swrid="5028293" athleteid="47068">
              <RESULTS>
                <RESULT eventid="44394" points="481" reactiontime="+63" swimtime="00:01:06.17" resultid="47069" heatid="50721" lane="8" entrytime="00:01:15.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="536" reactiontime="+76" swimtime="00:00:27.41" resultid="47070" heatid="50768" lane="7" entrytime="00:00:27.48" entrycourse="LCM" />
                <RESULT eventid="46298" points="568" reactiontime="+69" swimtime="00:00:25.24" resultid="47071" heatid="50820" lane="4" entrytime="00:00:25.87" entrycourse="LCM" />
                <RESULT eventid="46310" points="505" reactiontime="+60" swimtime="00:00:30.12" resultid="47072" heatid="50862" lane="0" entrytime="00:00:30.09" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Zdanowicz" birthdate="2005-11-25" gender="M" nation="POL" license="102401700017" swrid="5022561" athleteid="47054">
              <RESULTS>
                <RESULT eventid="44382" points="547" reactiontime="+63" swimtime="00:00:31.72" resultid="47055" heatid="50695" lane="7" entrytime="00:00:32.02" entrycourse="LCM" />
                <RESULT eventid="44407" points="520" reactiontime="+61" swimtime="00:01:10.72" resultid="47056" heatid="50750" lane="6" entrytime="00:01:11.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46302" points="489" reactiontime="+65" swimtime="00:02:40.04" resultid="47057" heatid="50839" lane="8" entrytime="00:02:39.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                    <SPLIT distance="100" swimtime="00:01:15.00" />
                    <SPLIT distance="150" swimtime="00:01:57.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karol" lastname="Słomski" birthdate="2003-03-07" gender="M" nation="POL" license="102401700023" swrid="4929873" athleteid="47058">
              <RESULTS>
                <RESULT eventid="44382" points="584" reactiontime="+67" swimtime="00:00:31.04" resultid="47059" heatid="50695" lane="3" entrytime="00:00:31.48" entrycourse="LCM" />
                <RESULT eventid="44411" points="535" reactiontime="+74" swimtime="00:00:27.43" resultid="47060" heatid="50894" lane="4" entrytime="00:00:28.34" entrycourse="LCM" />
                <RESULT eventid="46298" points="539" reactiontime="+70" swimtime="00:00:25.68" resultid="47061" heatid="50820" lane="6" entrytime="00:00:26.13" entrycourse="LCM" />
                <RESULT eventid="46310" points="462" reactiontime="+61" swimtime="00:00:31.03" resultid="47062" heatid="50861" lane="9" entrytime="00:00:32.36" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nina" lastname="Ganc" birthdate="2008-11-12" gender="F" nation="POL" license="102401600069" swrid="5354911" athleteid="47046">
              <RESULTS>
                <RESULT eventid="44380" points="434" reactiontime="+88" swimtime="00:01:08.29" resultid="47047" heatid="50680" lane="8" entrytime="00:01:25.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="389" reactiontime="+84" swimtime="00:02:34.64" resultid="47048" heatid="50741" lane="8" entrytime="00:02:35.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                    <SPLIT distance="100" swimtime="00:01:14.56" />
                    <SPLIT distance="150" swimtime="00:01:56.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="283" reactiontime="+75" swimtime="00:00:37.17" resultid="47049" heatid="50770" lane="8" />
                <RESULT eventid="46300" points="437" reactiontime="+74" swimtime="00:00:31.18" resultid="47050" heatid="50827" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patrycja" lastname="Stalska" birthdate="2008-05-31" gender="F" nation="POL" license="102401600080" swrid="5254261" athleteid="47063">
              <RESULTS>
                <RESULT eventid="44384" points="323" reactiontime="+78" swimtime="00:00:42.83" resultid="47064" heatid="50700" lane="1" entrytime="00:00:45.36" entrycourse="LCM" />
                <RESULT eventid="44396" points="290" reactiontime="+66" swimtime="00:01:26.88" resultid="47065" heatid="50725" lane="4" entrytime="00:01:24.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="357" reactiontime="+77" swimtime="00:00:33.35" resultid="47066" heatid="50829" lane="1" entrytime="00:00:33.76" entrycourse="LCM" />
                <RESULT eventid="46312" points="304" reactiontime="+63" swimtime="00:00:40.11" resultid="47067" heatid="50906" lane="0" entrytime="00:00:41.80" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Sieradzan" birthdate="2007-06-09" gender="M" nation="POL" license="102401700066" swrid="5220820" athleteid="47033">
              <RESULTS>
                <RESULT eventid="44378" points="375" reactiontime="+70" swimtime="00:01:05.03" resultid="47034" heatid="50668" lane="0" entrytime="00:01:07.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="291" reactiontime="+69" swimtime="00:00:33.57" resultid="47035" heatid="50763" lane="2" entrytime="00:00:33.85" entrycourse="LCM" />
                <RESULT eventid="46298" points="365" reactiontime="+59" swimtime="00:00:29.25" resultid="47036" heatid="50815" lane="4" entrytime="00:00:29.63" entrycourse="LCM" />
                <RESULT eventid="46310" points="248" reactiontime="+69" swimtime="00:00:38.15" resultid="47037" heatid="50857" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kornel" lastname="Pawłowski" birthdate="2008-06-05" gender="M" nation="POL" license="102401700052" swrid="5191077" athleteid="47019">
              <RESULTS>
                <RESULT eventid="44378" points="458" reactiontime="+74" swimtime="00:01:00.82" resultid="47020" heatid="50672" lane="8" entrytime="00:01:01.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="442" reactiontime="+71" swimtime="00:01:08.06" resultid="47021" heatid="50722" lane="3" entrytime="00:01:09.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="405" reactiontime="+73" swimtime="00:02:17.80" resultid="47022" heatid="50736" lane="3" entrytime="00:02:16.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.03" />
                    <SPLIT distance="100" swimtime="00:01:06.02" />
                    <SPLIT distance="150" swimtime="00:01:42.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="358" reactiontime="+71" swimtime="00:00:31.34" resultid="47023" heatid="50763" lane="4" entrytime="00:00:32.89" entrycourse="LCM" />
                <RESULT eventid="44415" points="396" reactiontime="+72" swimtime="00:02:32.39" resultid="47024" heatid="50783" lane="4" entrytime="00:02:32.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.05" />
                    <SPLIT distance="100" swimtime="00:01:14.93" />
                    <SPLIT distance="150" swimtime="00:01:54.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="397" reactiontime="+69" swimtime="00:00:28.43" resultid="47025" heatid="50817" lane="0" entrytime="00:00:28.40" entrycourse="LCM" />
                <RESULT eventid="46310" points="428" reactiontime="+72" swimtime="00:00:31.84" resultid="47026" heatid="50861" lane="7" entrytime="00:00:31.91" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Terka" birthdate="2006-05-25" gender="F" nation="POL" license="102401600035" swrid="5022556" athleteid="47038">
              <RESULTS>
                <RESULT eventid="44380" points="492" reactiontime="+75" swimtime="00:01:05.49" resultid="47039" heatid="50685" lane="2" entrytime="00:01:05.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="498" reactiontime="+49" swimtime="00:02:22.49" resultid="47040" heatid="50742" lane="4" entrytime="00:02:23.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                    <SPLIT distance="100" swimtime="00:01:09.58" />
                    <SPLIT distance="150" swimtime="00:01:47.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Bilski" birthdate="2002-08-09" gender="M" nation="POL" license="102401700057" swrid="5022574" athleteid="47073">
              <RESULTS>
                <RESULT eventid="44411" points="629" reactiontime="+62" swimtime="00:00:25.98" resultid="47074" heatid="50768" lane="2" entrytime="00:00:27.36" entrycourse="LCM" />
                <RESULT eventid="46298" points="580" reactiontime="+62" swimtime="00:00:25.06" resultid="47075" heatid="50821" lane="2" entrytime="00:00:25.42" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lena" lastname="Chodorowska" birthdate="2006-08-18" gender="F" nation="POL" license="102401600053" swrid="5113519" athleteid="47042">
              <RESULTS>
                <RESULT eventid="44380" points="589" reactiontime="+74" swimtime="00:01:01.66" resultid="47043" heatid="50687" lane="5" entrytime="00:01:01.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="615" reactiontime="+71" swimtime="00:00:27.82" resultid="47044" heatid="50835" lane="0" entrytime="00:00:27.95" entrycourse="LCM" />
                <RESULT eventid="46312" points="554" reactiontime="+80" swimtime="00:00:32.85" resultid="47045" heatid="50908" lane="2" entrytime="00:00:33.79" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mikołaj" lastname="Mosiak" birthdate="2003-01-02" gender="M" nation="POL" license="102401700015" swrid="4837654" athleteid="47027">
              <RESULTS>
                <RESULT eventid="44378" points="591" reactiontime="+63" swimtime="00:00:55.88" resultid="47028" heatid="50676" lane="9" entrytime="00:00:56.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="577" reactiontime="+64" swimtime="00:02:02.48" resultid="47029" heatid="50738" lane="5" entrytime="00:02:04.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.13" />
                    <SPLIT distance="100" swimtime="00:00:58.97" />
                    <SPLIT distance="150" swimtime="00:01:31.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="571" reactiontime="+64" swimtime="00:00:26.83" resultid="47030" heatid="50766" lane="0" entrytime="00:00:29.77" entrycourse="LCM" />
                <RESULT eventid="46298" points="571" reactiontime="+63" swimtime="00:00:25.20" resultid="47031" heatid="50819" lane="7" entrytime="00:00:26.51" entrycourse="LCM" />
                <RESULT eventid="46306" points="569" reactiontime="+65" swimtime="00:00:59.73" resultid="47032" heatid="50844" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jagoda" lastname="Reda" birthdate="2007-10-20" gender="F" nation="POL" license="102401600062" swrid="5220822" athleteid="47051">
              <RESULTS>
                <RESULT eventid="44380" points="415" reactiontime="+76" swimtime="00:01:09.27" resultid="47052" heatid="50682" lane="7" entrytime="00:01:10.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="431" reactiontime="+77" swimtime="00:00:31.32" resultid="47053" heatid="50830" lane="6" entrytime="00:00:31.60" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="95" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="44399" points="551" reactiontime="+62" swimtime="00:04:12.75" resultid="47076" heatid="50729" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                    <SPLIT distance="100" swimtime="00:01:05.15" />
                    <SPLIT distance="150" swimtime="00:01:37.06" />
                    <SPLIT distance="200" swimtime="00:02:15.71" />
                    <SPLIT distance="250" swimtime="00:02:43.92" />
                    <SPLIT distance="300" swimtime="00:03:16.33" />
                    <SPLIT distance="350" swimtime="00:03:42.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="47068" number="1" reactiontime="+62" />
                    <RELAYPOSITION athleteid="47054" number="2" reactiontime="+18" />
                    <RELAYPOSITION athleteid="47027" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="47073" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46289" points="584" reactiontime="+62" swimtime="00:03:45.15" resultid="47077" heatid="50794" lane="1" entrytime="00:03:53.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.24" />
                    <SPLIT distance="100" swimtime="00:00:56.90" />
                    <SPLIT distance="150" swimtime="00:01:23.00" />
                    <SPLIT distance="200" swimtime="00:01:51.74" />
                    <SPLIT distance="250" swimtime="00:02:18.57" />
                    <SPLIT distance="300" swimtime="00:02:47.93" />
                    <SPLIT distance="350" swimtime="00:03:14.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="47073" number="1" reactiontime="+62" />
                    <RELAYPOSITION athleteid="47027" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="47058" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="47068" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02201" nation="POL" region="01" clubid="49635" name="UKS Shark Rudna">
          <ATHLETES>
            <ATHLETE firstname="Weronika" lastname="Stembalska" birthdate="2007-01-15" gender="F" nation="POL" license="102201600096" swrid="5384598" athleteid="49651">
              <RESULTS>
                <RESULT eventid="44380" points="409" reactiontime="+74" swimtime="00:01:09.66" resultid="49652" heatid="50682" lane="9" entrytime="00:01:11.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="348" reactiontime="+75" swimtime="00:00:34.72" resultid="49653" heatid="50775" lane="5" entrytime="00:00:35.26" entrycourse="LCM" />
                <RESULT eventid="46300" points="467" reactiontime="+77" swimtime="00:00:30.50" resultid="49654" heatid="50831" lane="1" entrytime="00:00:30.77" entrycourse="LCM" />
                <RESULT eventid="46312" points="385" reactiontime="+66" swimtime="00:00:37.08" resultid="49655" heatid="50906" lane="4" entrytime="00:00:37.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Misiak" birthdate="2005-12-14" gender="M" nation="POL" license="102201700081" swrid="5135289" athleteid="49636">
              <RESULTS>
                <RESULT eventid="44378" points="650" reactiontime="+68" swimtime="00:00:54.14" resultid="49637" heatid="50676" lane="4" entrytime="00:00:54.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44390" points="549" reactiontime="+66" swimtime="00:02:19.16" resultid="49638" heatid="50707" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.83" />
                    <SPLIT distance="100" swimtime="00:01:06.39" />
                    <SPLIT distance="150" swimtime="00:01:46.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="566" reactiontime="+68" swimtime="00:02:03.30" resultid="49639" heatid="50738" lane="3" entrytime="00:02:05.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.68" />
                    <SPLIT distance="100" swimtime="00:00:58.97" />
                    <SPLIT distance="150" swimtime="00:01:31.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="655" reactiontime="+69" swimtime="00:00:25.64" resultid="49640" heatid="50769" lane="2" entrytime="00:00:25.61" entrycourse="LCM" />
                <RESULT eventid="46298" points="652" reactiontime="+56" swimtime="00:00:24.11" resultid="49641" heatid="50822" lane="2" entrytime="00:00:24.17" entrycourse="LCM" />
                <RESULT eventid="46306" points="617" reactiontime="+63" swimtime="00:00:58.13" resultid="49642" heatid="50849" lane="5" entrytime="00:00:58.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Adamczewska" birthdate="2004-04-06" gender="F" nation="POL" license="102201600092" swrid="5024285" athleteid="49662">
              <RESULTS>
                <RESULT eventid="44384" points="564" reactiontime="+67" swimtime="00:00:35.58" resultid="49663" heatid="50702" lane="4" entrytime="00:00:35.55" entrycourse="LCM" />
                <RESULT eventid="44409" points="521" reactiontime="+63" swimtime="00:01:19.68" resultid="49664" heatid="50755" lane="5" entrytime="00:01:18.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="523" reactiontime="+68" swimtime="00:00:30.31" resultid="49665" heatid="50779" lane="1" entrytime="00:00:29.95" entrycourse="LCM" />
                <RESULT eventid="46300" points="551" reactiontime="+69" swimtime="00:00:28.87" resultid="49666" heatid="50833" lane="2" entrytime="00:00:29.10" entrycourse="LCM" />
                <RESULT eventid="46308" points="528" reactiontime="+65" swimtime="00:01:08.63" resultid="49667" heatid="50900" lane="5" entrytime="00:01:10.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adela" lastname="Piskorska" birthdate="2003-11-16" gender="F" nation="POL" license="102201600099" swrid="4931147" athleteid="49675">
              <RESULTS>
                <RESULT eventid="44396" points="796" reactiontime="+57" swimtime="00:01:02.10" resultid="49676" heatid="50728" lane="4" entrytime="00:01:01.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44417" points="747" reactiontime="+57" swimtime="00:02:15.92" resultid="49677" heatid="50788" lane="4" entrytime="00:02:16.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                    <SPLIT distance="100" swimtime="00:01:05.45" />
                    <SPLIT distance="150" swimtime="00:01:40.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="791" reactiontime="+57" swimtime="00:00:29.17" resultid="49678" heatid="50909" lane="5" entrytime="00:00:28.78" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Trzpil" birthdate="2005-03-17" gender="M" nation="POL" license="102201700084" swrid="5148198" athleteid="49643">
              <RESULTS>
                <RESULT eventid="44378" points="554" reactiontime="+74" swimtime="00:00:57.09" resultid="49644" heatid="50675" lane="9" entrytime="00:00:57.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="476" reactiontime="+73" swimtime="00:00:33.23" resultid="49645" heatid="50695" lane="8" entrytime="00:00:32.42" entrycourse="LCM" />
                <RESULT eventid="44390" points="474" reactiontime="+78" swimtime="00:02:26.16" resultid="49646" heatid="50708" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.28" />
                    <SPLIT distance="100" swimtime="00:01:11.41" />
                    <SPLIT distance="150" swimtime="00:01:52.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="466" reactiontime="+75" swimtime="00:01:13.32" resultid="49647" heatid="50750" lane="1" entrytime="00:01:11.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="539" reactiontime="+75" swimtime="00:00:27.36" resultid="49648" heatid="50894" lane="3" entrytime="00:00:28.54" entrycourse="LCM" />
                <RESULT eventid="46298" points="546" reactiontime="+74" swimtime="00:00:25.58" resultid="49649" heatid="50820" lane="8" entrytime="00:00:26.20" entrycourse="LCM" />
                <RESULT eventid="46302" points="485" reactiontime="+75" swimtime="00:02:40.48" resultid="49650" heatid="50839" lane="7" entrytime="00:02:37.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                    <SPLIT distance="100" swimtime="00:01:17.43" />
                    <SPLIT distance="150" swimtime="00:01:59.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Kościelniak" birthdate="2002-06-07" gender="F" nation="POL" license="102201600063" swrid="4892800" athleteid="49668">
              <RESULTS>
                <RESULT eventid="44396" points="626" reactiontime="+63" swimtime="00:01:07.28" resultid="49669" heatid="50728" lane="6" entrytime="00:01:06.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="655" reactiontime="+64" swimtime="00:00:28.12" resultid="49670" heatid="50779" lane="4" entrytime="00:00:28.59" entrycourse="LCM" />
                <RESULT eventid="44417" points="632" reactiontime="+65" swimtime="00:02:23.67" resultid="49671" heatid="50788" lane="5" entrytime="00:02:22.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.03" />
                    <SPLIT distance="100" swimtime="00:01:11.36" />
                    <SPLIT distance="150" swimtime="00:01:48.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="604" reactiontime="+68" swimtime="00:00:28.00" resultid="49672" heatid="50835" lane="8" entrytime="00:00:27.93" entrycourse="LCM" />
                <RESULT eventid="46308" points="595" reactiontime="+70" swimtime="00:01:05.95" resultid="49673" heatid="50900" lane="4" entrytime="00:01:10.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="661" reactiontime="+62" swimtime="00:00:30.96" resultid="49674" heatid="50909" lane="6" entrytime="00:00:30.55" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Rybicka" birthdate="2006-04-09" gender="F" nation="POL" license="102201600097" swrid="5384596" athleteid="49656">
              <RESULTS>
                <RESULT eventid="44380" status="DNS" swimtime="00:00:00.00" resultid="49657" heatid="50679" lane="5" />
                <RESULT eventid="44384" status="DNS" swimtime="00:00:00.00" resultid="49658" heatid="50697" lane="5" />
                <RESULT eventid="44409" status="DNS" swimtime="00:00:00.00" resultid="49659" heatid="50753" lane="6" entrytime="00:01:36.95" entrycourse="LCM" />
                <RESULT eventid="46300" status="DNS" swimtime="00:00:00.00" resultid="49660" heatid="50825" lane="6" />
                <RESULT eventid="46304" status="DNS" swimtime="00:00:00.00" resultid="49661" heatid="50841" lane="8" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01713" nation="POL" region="13" clubid="46459">
          <ATHLETES>
            <ATHLETE firstname="Jacek" lastname="Sokulski" birthdate="1991-02-10" gender="M" nation="POL" license="101713700005" swrid="4062177" athleteid="46460">
              <RESULTS>
                <RESULT eventid="44378" status="DNS" swimtime="00:00:00.00" resultid="46461" heatid="50676" lane="3" entrytime="00:00:54.89" entrycourse="LCM" />
                <RESULT eventid="44411" points="701" reactiontime="+67" swimtime="00:00:25.06" resultid="46462" heatid="50769" lane="4" entrytime="00:00:24.82" entrycourse="LCM" />
                <RESULT eventid="46298" points="662" reactiontime="+65" swimtime="00:00:23.99" resultid="46463" heatid="50822" lane="7" entrytime="00:00:24.40" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01201" nation="POL" region="01" clubid="47582" name="MKS Piast Głogów">
          <ATHLETES>
            <ATHLETE firstname="Piotr" lastname="Musielak" birthdate="2006-07-13" gender="M" nation="POL" license="101201700260" swrid="5024279" athleteid="47625">
              <RESULTS>
                <RESULT eventid="44382" points="338" reactiontime="+53" swimtime="00:00:37.22" resultid="47626" heatid="50693" lane="9" entrytime="00:00:43.48" entrycourse="LCM" />
                <RESULT eventid="44407" points="314" reactiontime="+65" swimtime="00:01:23.66" resultid="47627" heatid="50747" lane="6" entrytime="00:01:33.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46302" status="DNS" swimtime="00:00:00.00" resultid="47628" heatid="50838" lane="6" entrytime="00:03:20.23" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Skokowski" birthdate="2005-01-13" gender="M" nation="POL" license="101201700239" swrid="5148191" athleteid="47583">
              <RESULTS>
                <RESULT eventid="44378" points="425" reactiontime="+78" swimtime="00:01:02.39" resultid="47584" heatid="50669" lane="9" entrytime="00:01:06.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="364" reactiontime="+76" swimtime="00:02:22.76" resultid="47585" heatid="50734" lane="5" entrytime="00:02:30.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                    <SPLIT distance="100" swimtime="00:01:09.21" />
                    <SPLIT distance="150" swimtime="00:01:47.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="348" reactiontime="+84" swimtime="00:00:31.65" resultid="47586" heatid="50763" lane="7" entrytime="00:00:34.29" entrycourse="LCM" />
                <RESULT eventid="46298" points="377" reactiontime="+88" swimtime="00:00:28.94" resultid="47587" heatid="50815" lane="6" entrytime="00:00:30.02" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Tywoniuk" birthdate="2008-06-10" gender="M" nation="POL" license="101201700357" swrid="5421084" athleteid="47593">
              <RESULTS>
                <RESULT eventid="44378" points="308" reactiontime="+74" swimtime="00:01:09.41" resultid="47594" heatid="50664" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="262" reactiontime="+85" swimtime="00:01:21.03" resultid="47595" heatid="50717" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="310" reactiontime="+73" swimtime="00:00:30.88" resultid="47596" heatid="50808" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Białas" birthdate="2006-03-08" gender="M" nation="POL" license="101201700252" swrid="4951837" athleteid="47637">
              <RESULTS>
                <RESULT eventid="44394" points="365" reactiontime="+73" swimtime="00:01:12.49" resultid="47638" heatid="50718" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="284" reactiontime="+66" swimtime="00:02:50.11" resultid="47639" heatid="50781" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.16" />
                    <SPLIT distance="150" swimtime="00:02:07.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="394" reactiontime="+71" swimtime="00:00:28.51" resultid="47640" heatid="50813" lane="5" entrytime="00:00:32.96" entrycourse="LCM" />
                <RESULT eventid="46310" points="392" reactiontime="+72" swimtime="00:00:32.77" resultid="47641" heatid="50859" lane="3" entrytime="00:00:39.74" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Klaudia" lastname="Wątroba" birthdate="2006-03-05" gender="F" nation="POL" license="101201600268" swrid="4901145" athleteid="47612">
              <RESULTS>
                <RESULT eventid="44380" points="387" reactiontime="+86" swimtime="00:01:10.93" resultid="47613" heatid="50681" lane="5" entrytime="00:01:12.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="289" reactiontime="+72" swimtime="00:00:36.92" resultid="47614" heatid="50774" lane="8" entrytime="00:00:40.39" entrycourse="LCM" />
                <RESULT eventid="46300" points="406" reactiontime="+67" swimtime="00:00:31.95" resultid="47615" heatid="50830" lane="9" entrytime="00:00:32.49" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcel" lastname="Piotrowski" birthdate="2007-03-24" gender="M" nation="POL" license="101201700278" swrid="5214663" athleteid="47620">
              <RESULTS>
                <RESULT eventid="44382" points="398" reactiontime="+80" swimtime="00:00:35.25" resultid="47621" heatid="50690" lane="3" />
                <RESULT eventid="44407" points="371" reactiontime="+78" swimtime="00:01:19.13" resultid="47622" heatid="50746" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="417" reactiontime="+80" swimtime="00:04:54.43" resultid="47623" heatid="50798" lane="7" entrytime="00:05:30.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                    <SPLIT distance="100" swimtime="00:01:08.55" />
                    <SPLIT distance="150" swimtime="00:01:46.72" />
                    <SPLIT distance="200" swimtime="00:02:24.93" />
                    <SPLIT distance="250" swimtime="00:03:03.78" />
                    <SPLIT distance="300" swimtime="00:03:41.77" />
                    <SPLIT distance="350" swimtime="00:04:19.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46302" points="347" reactiontime="+77" swimtime="00:02:59.33" resultid="47624" heatid="50837" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                    <SPLIT distance="100" swimtime="00:01:25.95" />
                    <SPLIT distance="150" swimtime="00:02:13.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Raś" birthdate="2007-02-17" gender="M" nation="POL" license="101201700279" swrid="5108615" athleteid="47602">
              <RESULTS>
                <RESULT eventid="44378" points="331" reactiontime="+70" swimtime="00:01:07.81" resultid="47603" heatid="50665" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="273" reactiontime="+82" swimtime="00:02:37.16" resultid="47604" heatid="50733" lane="2" entrytime="00:02:41.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.49" />
                    <SPLIT distance="100" swimtime="00:01:15.29" />
                    <SPLIT distance="150" swimtime="00:01:55.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="328" reactiontime="+78" swimtime="00:00:30.32" resultid="47605" heatid="50812" lane="1" entrytime="00:00:36.71" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartłomiej" lastname="Włodarczyk" birthdate="2005-02-05" gender="M" nation="POL" license="101201700248" swrid="5108614" athleteid="47588">
              <RESULTS>
                <RESULT eventid="44378" points="437" reactiontime="+71" swimtime="00:01:01.77" resultid="47589" heatid="50671" lane="9" entrytime="00:01:03.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="426" reactiontime="+83" swimtime="00:02:15.49" resultid="47590" heatid="50736" lane="2" entrytime="00:02:16.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                    <SPLIT distance="100" swimtime="00:01:05.30" />
                    <SPLIT distance="150" swimtime="00:01:40.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="390" reactiontime="+81" swimtime="00:00:30.46" resultid="47591" heatid="50765" lane="0" entrytime="00:00:31.24" entrycourse="LCM" />
                <RESULT eventid="46306" points="322" reactiontime="+73" swimtime="00:01:12.19" resultid="47592" heatid="50845" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Heiduk" birthdate="2005-04-05" gender="M" nation="POL" license="101201700222" swrid="5148189" athleteid="47633">
              <RESULTS>
                <RESULT eventid="44394" points="478" reactiontime="+71" swimtime="00:01:06.30" resultid="47634" heatid="50722" lane="5" entrytime="00:01:07.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="453" reactiontime="+75" swimtime="00:02:25.67" resultid="47635" heatid="50784" lane="9" entrytime="00:02:29.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                    <SPLIT distance="100" swimtime="00:01:09.16" />
                    <SPLIT distance="150" swimtime="00:01:47.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46310" points="494" reactiontime="+67" swimtime="00:00:30.35" resultid="47636" heatid="50861" lane="6" entrytime="00:00:31.35" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alicja" lastname="Musiał" birthdate="2005-03-30" gender="F" nation="POL" license="101201600229" swrid="5153489" athleteid="47629">
              <RESULTS>
                <RESULT eventid="44384" points="408" reactiontime="+80" swimtime="00:00:39.63" resultid="47630" heatid="50697" lane="3" />
                <RESULT eventid="44409" points="370" reactiontime="+78" swimtime="00:01:29.28" resultid="47631" heatid="50752" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46304" points="342" reactiontime="+77" swimtime="00:03:18.82" resultid="47632" heatid="50842" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.24" />
                    <SPLIT distance="100" swimtime="00:01:33.95" />
                    <SPLIT distance="150" swimtime="00:02:27.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Mita" birthdate="2006-07-06" gender="M" nation="POL" license="101201700259" swrid="4901150" athleteid="47597">
              <RESULTS>
                <RESULT eventid="44378" points="428" reactiontime="+73" swimtime="00:01:02.21" resultid="47598" heatid="50666" lane="3" entrytime="00:01:14.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="473" reactiontime="+69" swimtime="00:00:28.57" resultid="47599" heatid="50763" lane="8" entrytime="00:00:34.43" entrycourse="LCM" />
                <RESULT eventid="46298" points="423" reactiontime="+63" swimtime="00:00:27.84" resultid="47600" heatid="50813" lane="4" entrytime="00:00:32.88" entrycourse="LCM" />
                <RESULT eventid="46306" points="380" reactiontime="+52" swimtime="00:01:08.29" resultid="47601" heatid="50845" lane="4" entrytime="00:01:23.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT comment="-1" eventid="44399" reactiontime="+73" status="DSQ" swimtime="00:04:48.01" resultid="47642" heatid="50730" lane="8" entrytime="00:04:50.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                    <SPLIT distance="100" swimtime="00:01:12.24" />
                    <SPLIT distance="150" swimtime="00:01:49.29" />
                    <SPLIT distance="200" swimtime="00:02:34.40" />
                    <SPLIT distance="250" swimtime="00:03:04.54" />
                    <SPLIT distance="300" swimtime="00:03:42.40" />
                    <SPLIT distance="350" swimtime="00:04:12.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="47637" number="1" reactiontime="+73" status="DSQ" />
                    <RELAYPOSITION athleteid="47620" number="2" reactiontime="+67" status="DSQ" />
                    <RELAYPOSITION athleteid="47597" number="3" reactiontime="+54" status="DSQ" />
                    <RELAYPOSITION athleteid="47602" number="4" reactiontime="-17" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="S-3" eventid="46289" reactiontime="+73" status="DSQ" swimtime="00:00:00.00" resultid="47643" heatid="50794" lane="8" entrytime="00:04:08.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.26" />
                    <SPLIT distance="100" swimtime="00:01:03.26" />
                    <SPLIT distance="150" swimtime="00:01:32.20" />
                    <SPLIT distance="200" swimtime="00:02:04.70" />
                    <SPLIT distance="250" swimtime="00:02:35.96" />
                    <SPLIT distance="300" swimtime="00:03:12.34" />
                    <SPLIT distance="350" swimtime="00:03:41.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="47637" number="1" reactiontime="+73" status="DSQ" />
                    <RELAYPOSITION athleteid="47620" number="2" reactiontime="+43" status="DSQ" />
                    <RELAYPOSITION athleteid="47597" number="3" reactiontime="+27" status="DSQ" />
                    <RELAYPOSITION athleteid="47602" number="4" reactiontime="+63" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="95" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="46314" points="458" reactiontime="+78" swimtime="00:09:02.86" resultid="47644" heatid="50870" lane="5" entrytime="00:08:57.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                    <SPLIT distance="100" swimtime="00:01:03.70" />
                    <SPLIT distance="150" swimtime="00:01:40.25" />
                    <SPLIT distance="200" swimtime="00:02:17.24" />
                    <SPLIT distance="250" swimtime="00:02:46.80" />
                    <SPLIT distance="300" swimtime="00:03:20.73" />
                    <SPLIT distance="350" swimtime="00:03:57.03" />
                    <SPLIT distance="400" swimtime="00:04:33.56" />
                    <SPLIT distance="450" swimtime="00:05:02.32" />
                    <SPLIT distance="500" swimtime="00:05:35.24" />
                    <SPLIT distance="550" swimtime="00:06:10.10" />
                    <SPLIT distance="600" swimtime="00:06:44.88" />
                    <SPLIT distance="650" swimtime="00:07:15.45" />
                    <SPLIT distance="700" swimtime="00:07:51.32" />
                    <SPLIT distance="750" swimtime="00:08:28.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="47583" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="47588" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="47633" number="3" reactiontime="+60" />
                    <RELAYPOSITION athleteid="47620" number="4" reactiontime="+65" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="08114" nation="POL" region="14" clubid="49413" name="AZS  KU Uniwersytetu Warszawskiego">
          <ATHLETES>
            <ATHLETE firstname="Igor" lastname="Rębas" birthdate="1989-12-11" gender="M" nation="POL" license="508114700069" swrid="4251117" athleteid="49417">
              <RESULTS>
                <RESULT eventid="44378" points="634" reactiontime="+76" swimtime="00:00:54.60" resultid="49418" heatid="50677" lane="1" entrytime="00:00:53.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="508" reactiontime="+72" swimtime="00:02:07.76" resultid="49419" heatid="50739" lane="6" entrytime="00:01:59.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.44" />
                    <SPLIT distance="100" swimtime="00:01:00.70" />
                    <SPLIT distance="150" swimtime="00:01:34.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Micorek" birthdate="1993-08-25" gender="M" nation="POL" license="108114700041" swrid="4086676" athleteid="49414">
              <RESULTS>
                <RESULT eventid="44378" points="575" reactiontime="+69" swimtime="00:00:56.39" resultid="49415" heatid="50677" lane="9" entrytime="00:00:53.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="561" reactiontime="+75" swimtime="00:00:27.00" resultid="49416" heatid="50769" lane="8" entrytime="00:00:26.13" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Godlewski" birthdate="1996-05-26" gender="M" nation="POL" license="108114700059" swrid="4285522" athleteid="49420">
              <RESULTS>
                <RESULT eventid="44382" points="534" reactiontime="+71" swimtime="00:00:31.97" resultid="49421" heatid="50695" lane="1" entrytime="00:00:32.18" entrycourse="LCM" />
                <RESULT eventid="44407" points="463" reactiontime="+76" swimtime="00:01:13.48" resultid="49422" heatid="50745" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00901" nation="POL" region="01" clubid="48608" name="ULKS ,,Wodny Świat&apos;&apos;">
          <ATHLETES>
            <ATHLETE firstname="Kinga" lastname="Zabrzeska" birthdate="2007-05-16" gender="F" nation="POL" license="100901600040" swrid="5204359" athleteid="48616">
              <RESULTS>
                <RESULT eventid="44380" points="418" reactiontime="+69" swimtime="00:01:09.15" resultid="48617" heatid="50684" lane="9" entrytime="00:01:07.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44392" points="379" reactiontime="+70" swimtime="00:02:54.16" resultid="48618" heatid="50714" lane="9" entrytime="00:02:53.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.13" />
                    <SPLIT distance="100" swimtime="00:01:23.59" />
                    <SPLIT distance="150" swimtime="00:02:14.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="384" reactiontime="+67" swimtime="00:02:35.33" resultid="48619" heatid="50741" lane="9" entrytime="00:02:37.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.12" />
                    <SPLIT distance="100" swimtime="00:01:14.94" />
                    <SPLIT distance="150" swimtime="00:01:56.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="311" reactiontime="+58" swimtime="00:00:36.03" resultid="48620" heatid="50775" lane="4" entrytime="00:00:35.20" entrycourse="LCM" />
                <RESULT eventid="46300" points="452" reactiontime="+60" swimtime="00:00:30.82" resultid="48621" heatid="50830" lane="4" entrytime="00:00:31.12" entrycourse="LCM" />
                <RESULT eventid="46312" points="370" reactiontime="+74" swimtime="00:00:37.57" resultid="48622" heatid="50905" lane="9" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06401" nation="POL" region="01" clubid="46540" name="KS &quot;Swimmers Centrum Ślęza&quot;">
          <ATHLETES>
            <ATHLETE firstname="Julian" lastname="Stefurak" birthdate="2008-05-02" gender="M" nation="POL" license="106401700004" swrid="5311183" athleteid="46541">
              <RESULTS>
                <RESULT eventid="44382" points="296" reactiontime="+56" swimtime="00:00:38.93" resultid="46542" heatid="50690" lane="5" />
                <RESULT eventid="44407" points="276" reactiontime="+69" swimtime="00:01:27.26" resultid="46543" heatid="50748" lane="8" entrytime="00:01:26.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="272" reactiontime="+64" swimtime="00:00:34.37" resultid="46544" heatid="50758" lane="4" />
                <RESULT eventid="46302" points="305" reactiontime="+58" swimtime="00:03:07.22" resultid="46545" heatid="50837" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.36" />
                    <SPLIT distance="100" swimtime="00:01:31.21" />
                    <SPLIT distance="150" swimtime="00:02:20.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pola" lastname="Pietryk" birthdate="2008-09-26" gender="F" nation="POL" license="106401600002" swrid="5354927" athleteid="46546">
              <RESULTS>
                <RESULT eventid="46287" points="382" reactiontime="+83" swimtime="00:11:07.77" resultid="46547" heatid="50791" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.19" />
                    <SPLIT distance="100" swimtime="00:01:16.73" />
                    <SPLIT distance="150" swimtime="00:01:57.76" />
                    <SPLIT distance="200" swimtime="00:02:40.13" />
                    <SPLIT distance="250" swimtime="00:03:22.06" />
                    <SPLIT distance="300" swimtime="00:04:04.34" />
                    <SPLIT distance="350" swimtime="00:04:47.05" />
                    <SPLIT distance="400" swimtime="00:05:30.77" />
                    <SPLIT distance="450" swimtime="00:06:13.91" />
                    <SPLIT distance="500" swimtime="00:06:57.20" />
                    <SPLIT distance="550" swimtime="00:07:41.55" />
                    <SPLIT distance="600" swimtime="00:08:23.80" />
                    <SPLIT distance="650" swimtime="00:09:06.08" />
                    <SPLIT distance="700" swimtime="00:09:47.67" />
                    <SPLIT distance="750" swimtime="00:10:28.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="381" reactiontime="+85" swimtime="00:05:25.89" resultid="46548" heatid="50802" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                    <SPLIT distance="100" swimtime="00:01:15.25" />
                    <SPLIT distance="150" swimtime="00:01:56.93" />
                    <SPLIT distance="200" swimtime="00:02:38.54" />
                    <SPLIT distance="250" swimtime="00:03:21.19" />
                    <SPLIT distance="300" swimtime="00:04:03.20" />
                    <SPLIT distance="350" swimtime="00:04:45.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46308" points="266" reactiontime="+79" swimtime="00:01:26.24" resultid="46549" heatid="50899" lane="9" entrytime="00:01:22.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="05901" nation="POL" region="01" clubid="47659" name="UKP &quot;Na Fali&quot;">
          <ATHLETES>
            <ATHLETE firstname="Alan" lastname="Wojtowicz" birthdate="2008-04-29" gender="M" nation="POL" license="105901700004" swrid="5260082" athleteid="47660">
              <RESULTS>
                <RESULT eventid="44378" points="388" reactiontime="+64" swimtime="00:01:04.30" resultid="47661" heatid="50670" lane="8" entrytime="00:01:04.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="370" reactiontime="+68" swimtime="00:02:22.06" resultid="47662" heatid="50733" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.70" />
                    <SPLIT distance="100" swimtime="00:01:08.00" />
                    <SPLIT distance="150" swimtime="00:01:46.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="397" reactiontime="+66" swimtime="00:00:28.44" resultid="47663" heatid="50816" lane="5" entrytime="00:00:28.74" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Kodlew" birthdate="2005-01-12" gender="M" nation="POL" license="105901700002" swrid="5260110" athleteid="47664">
              <RESULTS>
                <RESULT eventid="44382" points="392" reactiontime="+74" swimtime="00:00:35.44" resultid="47665" heatid="50693" lane="5" entrytime="00:00:37.12" entrycourse="LCM" />
                <RESULT eventid="44403" points="485" reactiontime="+75" swimtime="00:02:09.81" resultid="47666" heatid="50737" lane="6" entrytime="00:02:12.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                    <SPLIT distance="100" swimtime="00:01:02.21" />
                    <SPLIT distance="150" swimtime="00:01:35.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="457" reactiontime="+75" swimtime="00:04:45.65" resultid="47667" heatid="50799" lane="1" entrytime="00:04:52.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                    <SPLIT distance="100" swimtime="00:01:06.94" />
                    <SPLIT distance="150" swimtime="00:01:42.94" />
                    <SPLIT distance="200" swimtime="00:02:20.31" />
                    <SPLIT distance="250" swimtime="00:02:58.05" />
                    <SPLIT distance="300" swimtime="00:03:35.85" />
                    <SPLIT distance="350" swimtime="00:04:12.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01101" nation="POL" region="01" clubid="47693" name="UKP Manta Jelcz-Laskowice">
          <ATHLETES>
            <ATHLETE firstname="Anna" lastname="Kicińska" birthdate="2004-05-14" gender="F" nation="POL" license="101101600042" swrid="5022564" athleteid="49111">
              <RESULTS>
                <RESULT eventid="44380" points="581" reactiontime="+66" swimtime="00:01:01.95" resultid="49112" heatid="50687" lane="9" entrytime="00:01:03.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44396" points="562" reactiontime="+68" swimtime="00:01:09.73" resultid="49113" heatid="50728" lane="2" entrytime="00:01:08.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="499" reactiontime="+73" swimtime="00:00:30.78" resultid="49114" heatid="50778" lane="7" entrytime="00:00:31.73" entrycourse="LCM" />
                <RESULT eventid="44417" points="478" reactiontime="+75" swimtime="00:02:37.66" resultid="49115" heatid="50788" lane="6" entrytime="00:02:30.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                    <SPLIT distance="100" swimtime="00:01:15.63" />
                    <SPLIT distance="150" swimtime="00:01:57.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="568" reactiontime="+78" swimtime="00:00:28.58" resultid="49116" heatid="50834" lane="2" entrytime="00:00:28.51" entrycourse="LCM" />
                <RESULT eventid="46312" points="572" reactiontime="+70" swimtime="00:00:32.49" resultid="49117" heatid="50909" lane="0" entrytime="00:00:32.28" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Piskorska" birthdate="2007-06-21" gender="F" nation="POL" license="101101600069" swrid="5416713" athleteid="49146">
              <RESULTS>
                <RESULT eventid="44380" points="431" reactiontime="+68" swimtime="00:01:08.45" resultid="49147" heatid="50679" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.49" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O-1" eventid="44396" status="DSQ" swimtime="00:01:16.78" resultid="49148" heatid="50727" lane="9" entrytime="00:01:17.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="358" reactiontime="+65" swimtime="00:00:34.40" resultid="49149" heatid="50773" lane="0" />
                <RESULT eventid="44417" points="410" reactiontime="+71" swimtime="00:02:45.97" resultid="49150" heatid="50787" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.44" />
                    <SPLIT distance="100" swimtime="00:01:21.97" />
                    <SPLIT distance="150" swimtime="00:02:04.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" status="DNS" swimtime="00:00:00.00" resultid="49151" heatid="50803" lane="5" />
                <RESULT eventid="46312" status="DNS" swimtime="00:00:00.00" resultid="49152" heatid="50905" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Wilgosz" birthdate="2005-04-10" gender="F" nation="POL" license="101101600032" swrid="5088625" athleteid="49153">
              <RESULTS>
                <RESULT eventid="44380" status="DNS" swimtime="00:00:00.00" resultid="49154" heatid="50687" lane="6" entrytime="00:01:02.25" entrycourse="LCM" />
                <RESULT eventid="44405" points="523" reactiontime="+69" swimtime="00:02:20.17" resultid="49156" heatid="50744" lane="9" entrytime="00:02:16.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                    <SPLIT distance="100" swimtime="00:01:07.48" />
                    <SPLIT distance="150" swimtime="00:01:43.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" status="DNS" swimtime="00:00:00.00" resultid="49158" heatid="50805" lane="0" entrytime="00:04:54.91" entrycourse="LCM" />
                <RESULT eventid="46300" points="513" reactiontime="+71" swimtime="00:00:29.55" resultid="49159" heatid="50834" lane="8" entrytime="00:00:28.63" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Paprocki" birthdate="2008-05-19" gender="M" nation="POL" license="101101700077" swrid="5462493" athleteid="49094">
              <RESULTS>
                <RESULT eventid="44378" points="255" reactiontime="+78" swimtime="00:01:13.94" resultid="49095" heatid="50666" lane="6" entrytime="00:01:15.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="197" reactiontime="+93" swimtime="00:01:29.10" resultid="49096" heatid="50718" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="207" reactiontime="+82" swimtime="00:02:52.19" resultid="49097" heatid="50733" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.64" />
                    <SPLIT distance="100" swimtime="00:01:22.83" />
                    <SPLIT distance="150" swimtime="00:02:10.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="177" reactiontime="+81" swimtime="00:01:41.18" resultid="49098" heatid="50746" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="242" swimtime="00:00:33.53" resultid="49099" heatid="50807" lane="4" />
                <RESULT eventid="46310" points="205" reactiontime="+89" swimtime="00:00:40.69" resultid="49100" heatid="50857" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hanna" lastname="Misiewicz" birthdate="2008-05-11" gender="F" nation="POL" license="101101600066" swrid="5244049" athleteid="49132">
              <RESULTS>
                <RESULT eventid="44380" points="431" reactiontime="+80" swimtime="00:01:08.41" resultid="49133" heatid="50684" lane="8" entrytime="00:01:07.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44396" points="318" reactiontime="+88" swimtime="00:01:24.34" resultid="49134" heatid="50726" lane="1" entrytime="00:01:22.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="382" reactiontime="+84" swimtime="00:02:35.60" resultid="49135" heatid="50741" lane="2" entrytime="00:02:34.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                    <SPLIT distance="100" swimtime="00:01:17.02" />
                    <SPLIT distance="150" swimtime="00:01:58.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="328" reactiontime="+77" swimtime="00:00:35.41" resultid="49136" heatid="50774" lane="9" entrytime="00:00:42.51" entrycourse="LCM" />
                <RESULT eventid="46296" points="360" reactiontime="+59" swimtime="00:05:32.25" resultid="49137" heatid="50802" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                    <SPLIT distance="100" swimtime="00:01:18.24" />
                    <SPLIT distance="150" swimtime="00:02:00.83" />
                    <SPLIT distance="200" swimtime="00:02:44.46" />
                    <SPLIT distance="250" swimtime="00:03:27.79" />
                    <SPLIT distance="300" swimtime="00:04:10.11" />
                    <SPLIT distance="350" swimtime="00:04:52.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46308" status="DNS" swimtime="00:00:00.00" resultid="49138" heatid="50898" lane="5" entrytime="00:01:25.60" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Kobuszyński" birthdate="2006-02-22" gender="M" nation="POL" license="101101700049" swrid="5191089" athleteid="49080">
              <RESULTS>
                <RESULT eventid="44378" points="428" reactiontime="+48" swimtime="00:01:02.21" resultid="49081" heatid="50665" lane="4" entrytime="00:01:37.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="401" reactiontime="+58" swimtime="00:01:10.26" resultid="49082" heatid="50720" lane="7" entrytime="00:01:19.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="404" reactiontime="+60" swimtime="00:00:30.12" resultid="49083" heatid="50763" lane="0" entrytime="00:00:35.07" entrycourse="LCM" />
                <RESULT eventid="44415" points="360" reactiontime="+60" swimtime="00:02:37.26" resultid="49084" heatid="50782" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                    <SPLIT distance="100" swimtime="00:01:17.33" />
                    <SPLIT distance="150" swimtime="00:01:59.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="436" reactiontime="+60" swimtime="00:00:27.56" resultid="49085" heatid="50814" lane="1" entrytime="00:00:32.58" entrycourse="LCM" />
                <RESULT eventid="46310" points="399" reactiontime="+56" swimtime="00:00:32.58" resultid="49086" heatid="50859" lane="0" entrytime="00:00:51.24" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Kłak" birthdate="2006-11-11" gender="F" nation="POL" license="101101600067" swrid="5088628" athleteid="49118">
              <RESULTS>
                <RESULT eventid="44380" points="458" reactiontime="+76" swimtime="00:01:07.08" resultid="49119" heatid="50680" lane="9" entrytime="00:01:27.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44384" points="451" reactiontime="+77" swimtime="00:00:38.32" resultid="49120" heatid="50699" lane="3" entrytime="00:00:53.57" entrycourse="LCM" />
                <RESULT eventid="44413" status="DNS" swimtime="00:00:00.00" resultid="49121" heatid="50771" lane="2" />
                <RESULT eventid="46300" status="DNS" swimtime="00:00:00.00" resultid="49122" heatid="50828" lane="7" entrytime="00:00:38.16" entrycourse="LCM" />
                <RESULT eventid="46304" points="394" reactiontime="+74" swimtime="00:03:09.71" resultid="49123" heatid="50842" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.04" />
                    <SPLIT distance="100" swimtime="00:01:30.61" />
                    <SPLIT distance="150" swimtime="00:02:20.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="373" reactiontime="+89" swimtime="00:00:37.47" resultid="49124" heatid="50903" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olivia" lastname="Sławińska" birthdate="2006-04-28" gender="F" nation="POL" license="101101600057" swrid="5253970" athleteid="49181">
              <RESULTS>
                <RESULT eventid="44384" points="515" reactiontime="+72" swimtime="00:00:36.67" resultid="49182" heatid="50702" lane="1" entrytime="00:00:36.68" entrycourse="LCM" />
                <RESULT eventid="44392" points="469" reactiontime="+69" swimtime="00:02:42.25" resultid="49183" heatid="50715" lane="0" entrytime="00:02:44.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.60" />
                    <SPLIT distance="100" swimtime="00:01:18.82" />
                    <SPLIT distance="150" swimtime="00:02:04.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44409" points="489" reactiontime="+71" swimtime="00:01:21.35" resultid="49184" heatid="50755" lane="7" entrytime="00:01:22.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="410" reactiontime="+68" swimtime="00:00:32.87" resultid="49185" heatid="50776" lane="9" entrytime="00:00:35.14" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oskar" lastname="Wołodko" birthdate="2005-11-23" gender="M" nation="POL" license="101101700058" swrid="5160043" athleteid="49174">
              <RESULTS>
                <RESULT eventid="44382" points="489" reactiontime="+68" swimtime="00:00:32.93" resultid="49175" heatid="50693" lane="2" entrytime="00:00:38.86" entrycourse="LCM" />
                <RESULT eventid="44390" points="434" reactiontime="+72" swimtime="00:02:30.57" resultid="49176" heatid="50707" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.06" />
                    <SPLIT distance="100" swimtime="00:01:12.83" />
                    <SPLIT distance="150" swimtime="00:01:55.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="490" reactiontime="+70" swimtime="00:01:12.11" resultid="49177" heatid="50748" lane="7" entrytime="00:01:26.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="406" reactiontime="+64" swimtime="00:00:30.07" resultid="49178" heatid="50761" lane="2" />
                <RESULT eventid="46294" points="468" reactiontime="+67" swimtime="00:04:43.39" resultid="49179" heatid="50798" lane="5" entrytime="00:05:05.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.52" />
                    <SPLIT distance="100" swimtime="00:01:04.48" />
                    <SPLIT distance="150" swimtime="00:01:40.20" />
                    <SPLIT distance="200" swimtime="00:02:17.19" />
                    <SPLIT distance="250" swimtime="00:02:53.74" />
                    <SPLIT distance="300" swimtime="00:03:31.05" />
                    <SPLIT distance="350" swimtime="00:04:08.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46302" points="476" reactiontime="+67" swimtime="00:02:41.42" resultid="49180" heatid="50838" lane="3" entrytime="00:03:09.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="100" swimtime="00:01:16.49" />
                    <SPLIT distance="150" swimtime="00:01:58.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Drzycimski" birthdate="2007-12-07" gender="M" nation="POL" license="101101700070" swrid="5287801" athleteid="49073">
              <RESULTS>
                <RESULT eventid="44378" points="359" reactiontime="+88" swimtime="00:01:06.00" resultid="49074" heatid="50670" lane="0" entrytime="00:01:04.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="289" reactiontime="+95" swimtime="00:01:18.41" resultid="49075" heatid="50718" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="323" reactiontime="+87" swimtime="00:02:28.54" resultid="49076" heatid="50732" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                    <SPLIT distance="100" swimtime="00:01:13.07" />
                    <SPLIT distance="150" swimtime="00:01:51.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="309" reactiontime="+83" swimtime="00:00:32.91" resultid="49077" heatid="50759" lane="1" />
                <RESULT eventid="46298" points="348" reactiontime="+82" swimtime="00:00:29.72" resultid="49078" heatid="50810" lane="1" />
                <RESULT eventid="46310" points="276" reactiontime="+78" swimtime="00:00:36.83" resultid="49079" heatid="50857" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Cholewa" birthdate="2008-05-18" gender="F" nation="POL" license="101101600065" swrid="5287802" athleteid="49104">
              <RESULTS>
                <RESULT eventid="44380" points="336" reactiontime="+88" swimtime="00:01:14.35" resultid="49105" heatid="50681" lane="3" entrytime="00:01:13.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44396" points="291" reactiontime="+75" swimtime="00:01:26.85" resultid="49106" heatid="50724" lane="4" entrytime="00:01:29.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="291" reactiontime="+94" swimtime="00:02:50.39" resultid="49107" heatid="50740" lane="7" entrytime="00:02:44.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.43" />
                    <SPLIT distance="100" swimtime="00:01:22.27" />
                    <SPLIT distance="150" swimtime="00:02:08.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="331" reactiontime="+95" swimtime="00:00:35.30" resultid="49108" heatid="50773" lane="3" entrytime="00:00:46.96" entrycourse="LCM" />
                <RESULT eventid="46296" points="309" reactiontime="+92" swimtime="00:05:49.51" resultid="49109" heatid="50802" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.20" />
                    <SPLIT distance="100" swimtime="00:01:20.76" />
                    <SPLIT distance="150" swimtime="00:02:05.77" />
                    <SPLIT distance="200" swimtime="00:02:51.09" />
                    <SPLIT distance="250" swimtime="00:03:36.45" />
                    <SPLIT distance="300" swimtime="00:04:21.72" />
                    <SPLIT distance="350" swimtime="00:05:07.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="267" reactiontime="+70" swimtime="00:00:41.85" resultid="49110" heatid="50905" lane="6" entrytime="00:00:45.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Włodarczyk" birthdate="2008-03-03" gender="F" nation="POL" license="101101600064" swrid="5287617" athleteid="49160">
              <RESULTS>
                <RESULT eventid="44380" points="410" reactiontime="+67" swimtime="00:01:09.55" resultid="49161" heatid="50683" lane="1" entrytime="00:01:09.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44396" points="355" reactiontime="+77" swimtime="00:01:21.28" resultid="49162" heatid="50725" lane="6" entrytime="00:01:25.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="414" reactiontime="+56" swimtime="00:02:31.52" resultid="49163" heatid="50740" lane="4" entrytime="00:02:37.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.07" />
                    <SPLIT distance="100" swimtime="00:01:14.03" />
                    <SPLIT distance="150" swimtime="00:01:52.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="317" reactiontime="+53" swimtime="00:00:35.81" resultid="49164" heatid="50773" lane="4" entrytime="00:00:43.63" entrycourse="LCM" />
                <RESULT eventid="46296" points="402" reactiontime="+71" swimtime="00:05:20.23" resultid="49165" heatid="50803" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.82" />
                    <SPLIT distance="100" swimtime="00:01:17.10" />
                    <SPLIT distance="150" swimtime="00:01:58.70" />
                    <SPLIT distance="200" swimtime="00:02:39.78" />
                    <SPLIT distance="250" swimtime="00:03:21.45" />
                    <SPLIT distance="300" swimtime="00:04:02.68" />
                    <SPLIT distance="350" swimtime="00:04:43.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46308" points="308" reactiontime="+72" swimtime="00:01:22.15" resultid="49166" heatid="50898" lane="3" entrytime="00:01:26.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Laszczak" birthdate="2007-02-26" gender="F" nation="POL" license="101101600053" swrid="5191091" athleteid="49125">
              <RESULTS>
                <RESULT eventid="44380" points="470" reactiontime="+77" swimtime="00:01:06.47" resultid="49126" heatid="50683" lane="9" entrytime="00:01:09.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44396" points="481" reactiontime="+75" swimtime="00:01:13.47" resultid="49127" heatid="50727" lane="4" entrytime="00:01:13.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="469" reactiontime="+79" swimtime="00:02:25.33" resultid="49128" heatid="50742" lane="7" entrytime="00:02:26.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                    <SPLIT distance="100" swimtime="00:01:11.04" />
                    <SPLIT distance="150" swimtime="00:01:50.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44417" points="467" reactiontime="+76" swimtime="00:02:38.90" resultid="49129" heatid="50788" lane="0" entrytime="00:02:41.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.00" />
                    <SPLIT distance="100" swimtime="00:01:18.06" />
                    <SPLIT distance="150" swimtime="00:01:59.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="435" reactiontime="+79" swimtime="00:05:11.97" resultid="49130" heatid="50804" lane="1" entrytime="00:05:36.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                    <SPLIT distance="100" swimtime="00:01:11.55" />
                    <SPLIT distance="150" swimtime="00:01:50.84" />
                    <SPLIT distance="200" swimtime="00:02:30.64" />
                    <SPLIT distance="250" swimtime="00:03:11.01" />
                    <SPLIT distance="300" swimtime="00:03:51.93" />
                    <SPLIT distance="350" swimtime="00:04:33.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="499" reactiontime="+68" swimtime="00:00:34.00" resultid="49131" heatid="50908" lane="0" entrytime="00:00:35.31" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roman" lastname="Żerek" birthdate="1988-02-01" gender="M" nation="POL" license="101101700074" swrid="4072671" athleteid="49101">
              <RESULTS>
                <RESULT eventid="44378" points="435" reactiontime="+72" swimtime="00:01:01.88" resultid="49102" heatid="50665" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="492" reactiontime="+70" swimtime="00:00:26.47" resultid="49103" heatid="50818" lane="2" entrytime="00:00:27.04" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Wołodko" birthdate="2007-08-23" gender="M" nation="POL" license="101101700059" swrid="4917952" athleteid="49167">
              <RESULTS>
                <RESULT eventid="44382" points="368" reactiontime="+64" swimtime="00:00:36.21" resultid="49168" heatid="50693" lane="0" entrytime="00:00:43.03" entrycourse="LCM" />
                <RESULT eventid="44390" points="310" reactiontime="+66" swimtime="00:02:48.42" resultid="49169" heatid="50709" lane="7" entrytime="00:02:47.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                    <SPLIT distance="100" swimtime="00:01:22.28" />
                    <SPLIT distance="150" swimtime="00:02:09.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="299" reactiontime="+64" swimtime="00:01:24.99" resultid="49170" heatid="50747" lane="0" entrytime="00:01:42.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="287" reactiontime="+65" swimtime="00:00:33.76" resultid="49171" heatid="50758" lane="5" />
                <RESULT eventid="46298" points="311" reactiontime="+54" swimtime="00:00:30.83" resultid="49172" heatid="50812" lane="4" entrytime="00:00:35.63" entrycourse="LCM" />
                <RESULT eventid="46302" points="280" reactiontime="+68" swimtime="00:03:12.72" resultid="49173" heatid="50837" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.09" />
                    <SPLIT distance="100" swimtime="00:01:34.11" />
                    <SPLIT distance="150" swimtime="00:02:23.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwier" lastname="Pańka" birthdate="2007-05-23" gender="M" nation="POL" license="101101700056" swrid="5316786" athleteid="49087">
              <RESULTS>
                <RESULT eventid="44378" points="318" reactiontime="+66" swimtime="00:01:08.66" resultid="49088" heatid="50667" lane="3" entrytime="00:01:08.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="298" reactiontime="+62" swimtime="00:01:17.54" resultid="49089" heatid="50720" lane="3" entrytime="00:01:18.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="276" reactiontime="+67" swimtime="00:02:36.57" resultid="49090" heatid="50733" lane="3" entrytime="00:02:36.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                    <SPLIT distance="100" swimtime="00:01:16.01" />
                    <SPLIT distance="150" swimtime="00:01:58.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="314" reactiontime="+61" swimtime="00:02:44.52" resultid="49091" heatid="50782" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.77" />
                    <SPLIT distance="100" swimtime="00:01:21.75" />
                    <SPLIT distance="150" swimtime="00:02:04.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="301" reactiontime="+62" swimtime="00:00:31.17" resultid="49092" heatid="50812" lane="9" entrytime="00:00:38.29" entrycourse="LCM" />
                <RESULT eventid="46310" points="315" reactiontime="+60" swimtime="00:00:35.26" resultid="49093" heatid="50859" lane="6" entrytime="00:00:40.37" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicola" lastname="Piebiak" birthdate="2008-05-12" gender="F" nation="POL" license="101101600060" swrid="5212910" athleteid="49139">
              <RESULTS>
                <RESULT eventid="44380" points="563" reactiontime="+78" swimtime="00:01:02.59" resultid="49140" heatid="50687" lane="8" entrytime="00:01:02.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44392" points="463" reactiontime="+82" swimtime="00:02:43.00" resultid="49141" heatid="50715" lane="7" entrytime="00:02:41.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                    <SPLIT distance="100" swimtime="00:01:17.41" />
                    <SPLIT distance="150" swimtime="00:02:07.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="516" reactiontime="+80" swimtime="00:02:20.79" resultid="49142" heatid="50743" lane="9" entrytime="00:02:22.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.42" />
                    <SPLIT distance="100" swimtime="00:01:09.03" />
                    <SPLIT distance="150" swimtime="00:01:46.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44417" points="486" reactiontime="+71" swimtime="00:02:36.87" resultid="49143" heatid="50785" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.49" />
                    <SPLIT distance="100" swimtime="00:01:17.81" />
                    <SPLIT distance="150" swimtime="00:01:58.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="483" reactiontime="+83" swimtime="00:05:01.35" resultid="49144" heatid="50803" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                    <SPLIT distance="100" swimtime="00:01:11.81" />
                    <SPLIT distance="150" swimtime="00:01:51.80" />
                    <SPLIT distance="200" swimtime="00:02:31.31" />
                    <SPLIT distance="250" swimtime="00:03:09.49" />
                    <SPLIT distance="300" swimtime="00:03:48.04" />
                    <SPLIT distance="350" swimtime="00:04:26.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="535" reactiontime="+80" swimtime="00:00:29.15" resultid="49145" heatid="50831" lane="4" entrytime="00:00:30.11" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="95" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="44399" points="386" reactiontime="+66" swimtime="00:04:44.66" resultid="49188" heatid="50729" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="100" swimtime="00:01:15.49" />
                    <SPLIT distance="150" swimtime="00:01:49.66" />
                    <SPLIT distance="200" swimtime="00:02:28.08" />
                    <SPLIT distance="250" swimtime="00:02:59.38" />
                    <SPLIT distance="300" swimtime="00:03:38.05" />
                    <SPLIT distance="350" swimtime="00:04:11.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="49087" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="49174" number="2" reactiontime="+23" />
                    <RELAYPOSITION athleteid="49080" number="3" reactiontime="+14" />
                    <RELAYPOSITION athleteid="49073" number="4" reactiontime="+63" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46289" points="374" reactiontime="+70" swimtime="00:04:21.14" resultid="49191" heatid="50793" lane="6" entrytime="00:04:56.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.70" />
                    <SPLIT distance="100" swimtime="00:01:00.15" />
                    <SPLIT distance="150" swimtime="00:01:29.86" />
                    <SPLIT distance="200" swimtime="00:02:04.92" />
                    <SPLIT distance="250" swimtime="00:02:38.46" />
                    <SPLIT distance="300" swimtime="00:03:12.55" />
                    <SPLIT distance="350" swimtime="00:03:45.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="49174" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="49080" number="2" />
                    <RELAYPOSITION athleteid="49073" number="3" />
                    <RELAYPOSITION athleteid="49167" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46314" points="363" reactiontime="+73" swimtime="00:09:46.48" resultid="49194" heatid="50870" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.06" />
                    <SPLIT distance="100" swimtime="00:01:03.72" />
                    <SPLIT distance="150" swimtime="00:01:39.12" />
                    <SPLIT distance="200" swimtime="00:02:14.11" />
                    <SPLIT distance="250" swimtime="00:02:45.42" />
                    <SPLIT distance="300" swimtime="00:03:22.95" />
                    <SPLIT distance="350" swimtime="00:04:02.60" />
                    <SPLIT distance="400" swimtime="00:04:40.96" />
                    <SPLIT distance="450" swimtime="00:05:16.69" />
                    <SPLIT distance="500" swimtime="00:05:55.81" />
                    <SPLIT distance="550" swimtime="00:06:35.73" />
                    <SPLIT distance="600" swimtime="00:07:11.76" />
                    <SPLIT distance="650" swimtime="00:07:46.87" />
                    <SPLIT distance="700" swimtime="00:08:27.94" />
                    <SPLIT distance="750" swimtime="00:09:09.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="49174" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="49080" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="49073" number="3" reactiontime="+58" />
                    <RELAYPOSITION athleteid="49167" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="95" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="44401" points="496" reactiontime="+74" swimtime="00:04:50.97" resultid="49189" heatid="50887" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.91" />
                    <SPLIT distance="100" swimtime="00:01:13.82" />
                    <SPLIT distance="150" swimtime="00:01:50.70" />
                    <SPLIT distance="200" swimtime="00:02:34.71" />
                    <SPLIT distance="250" swimtime="00:03:07.43" />
                    <SPLIT distance="300" swimtime="00:03:48.08" />
                    <SPLIT distance="350" swimtime="00:04:17.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="49125" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="49181" number="2" reactiontime="+22" />
                    <RELAYPOSITION athleteid="49111" number="3" reactiontime="-1" />
                    <RELAYPOSITION athleteid="49153" number="4" reactiontime="-14" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46291" points="534" reactiontime="+76" swimtime="00:04:18.75" resultid="49192" heatid="50795" lane="2" entrytime="00:04:20.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.45" />
                    <SPLIT distance="100" swimtime="00:01:02.95" />
                    <SPLIT distance="150" swimtime="00:01:33.69" />
                    <SPLIT distance="200" swimtime="00:02:08.34" />
                    <SPLIT distance="250" swimtime="00:02:39.38" />
                    <SPLIT distance="300" swimtime="00:03:15.25" />
                    <SPLIT distance="350" swimtime="00:03:45.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="49153" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="49181" number="2" reactiontime="+25" />
                    <RELAYPOSITION athleteid="49125" number="3" reactiontime="+17" />
                    <RELAYPOSITION athleteid="49111" number="4" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46316" points="484" reactiontime="+73" swimtime="00:09:47.69" resultid="49195" heatid="50871" lane="5" entrytime="00:09:34.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                    <SPLIT distance="100" swimtime="00:01:08.71" />
                    <SPLIT distance="150" swimtime="00:01:46.78" />
                    <SPLIT distance="200" swimtime="00:02:23.71" />
                    <SPLIT distance="250" swimtime="00:02:55.85" />
                    <SPLIT distance="300" swimtime="00:03:32.74" />
                    <SPLIT distance="350" swimtime="00:04:10.40" />
                    <SPLIT distance="400" swimtime="00:04:46.00" />
                    <SPLIT distance="450" swimtime="00:05:21.70" />
                    <SPLIT distance="500" swimtime="00:06:00.96" />
                    <SPLIT distance="550" swimtime="00:06:40.84" />
                    <SPLIT distance="600" swimtime="00:07:18.81" />
                    <SPLIT distance="650" swimtime="00:07:51.98" />
                    <SPLIT distance="700" swimtime="00:08:30.35" />
                    <SPLIT distance="750" swimtime="00:09:10.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="49153" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="49111" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="49118" number="3" reactiontime="+26" />
                    <RELAYPOSITION athleteid="49125" number="4" reactiontime="+3" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="44401" points="373" reactiontime="+74" swimtime="00:05:19.82" resultid="49190" heatid="50731" lane="1" entrytime="00:05:27.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                    <SPLIT distance="100" swimtime="00:01:13.21" />
                    <SPLIT distance="150" swimtime="00:01:58.36" />
                    <SPLIT distance="200" swimtime="00:02:49.84" />
                    <SPLIT distance="250" swimtime="00:03:26.45" />
                    <SPLIT distance="300" swimtime="00:04:10.45" />
                    <SPLIT distance="350" swimtime="00:04:43.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="49139" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="49104" number="2" reactiontime="+76" />
                    <RELAYPOSITION athleteid="49160" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="49132" number="4" reactiontime="+11" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46291" points="427" reactiontime="+88" swimtime="00:04:38.80" resultid="49193" heatid="50795" lane="1" entrytime="00:04:32.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                    <SPLIT distance="100" swimtime="00:01:04.05" />
                    <SPLIT distance="150" swimtime="00:01:36.70" />
                    <SPLIT distance="200" swimtime="00:02:13.33" />
                    <SPLIT distance="250" swimtime="00:02:48.16" />
                    <SPLIT distance="300" swimtime="00:03:27.88" />
                    <SPLIT distance="350" swimtime="00:04:01.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="49139" number="1" reactiontime="+88" />
                    <RELAYPOSITION athleteid="49132" number="2" reactiontime="+29" />
                    <RELAYPOSITION athleteid="49104" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="49160" number="4" reactiontime="+7" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46316" points="405" reactiontime="+84" swimtime="00:10:23.28" resultid="49196" heatid="50871" lane="2" entrytime="00:10:17.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.75" />
                    <SPLIT distance="100" swimtime="00:01:07.66" />
                    <SPLIT distance="150" swimtime="00:01:45.63" />
                    <SPLIT distance="200" swimtime="00:02:20.78" />
                    <SPLIT distance="250" swimtime="00:02:55.14" />
                    <SPLIT distance="300" swimtime="00:03:36.13" />
                    <SPLIT distance="350" swimtime="00:04:18.36" />
                    <SPLIT distance="400" swimtime="00:04:57.02" />
                    <SPLIT distance="450" swimtime="00:05:32.47" />
                    <SPLIT distance="500" swimtime="00:06:12.65" />
                    <SPLIT distance="550" swimtime="00:06:53.40" />
                    <SPLIT distance="600" swimtime="00:07:33.44" />
                    <SPLIT distance="650" swimtime="00:08:11.26" />
                    <SPLIT distance="700" swimtime="00:08:55.62" />
                    <SPLIT distance="750" swimtime="00:09:41.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="49139" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="49132" number="2" reactiontime="+19" />
                    <RELAYPOSITION athleteid="49160" number="3" reactiontime="+25" />
                    <RELAYPOSITION athleteid="49104" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02101" nation="POL" region="01" clubid="47884" name="UKS &apos;&apos;ORKA&apos;&apos; Lubań">
          <ATHLETES>
            <ATHLETE firstname="Julita" lastname="Jośko" birthdate="2004-04-30" gender="F" nation="POL" license="102101600129" swrid="4910964" athleteid="47906">
              <RESULTS>
                <RESULT eventid="44380" points="408" reactiontime="+74" swimtime="00:01:09.71" resultid="47907" heatid="50679" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44396" points="406" reactiontime="+73" swimtime="00:01:17.72" resultid="47908" heatid="50724" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="272" reactiontime="+74" swimtime="00:00:37.66" resultid="47909" heatid="50774" lane="7" entrytime="00:00:39.80" entrycourse="LCM" />
                <RESULT eventid="46300" points="488" reactiontime="+75" swimtime="00:00:30.05" resultid="47910" heatid="50826" lane="4" />
                <RESULT eventid="46312" points="450" reactiontime="+79" swimtime="00:00:35.19" resultid="47911" heatid="50906" lane="2" entrytime="00:00:39.73" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Iga" lastname="Krasowska" birthdate="2006-04-23" gender="F" nation="POL" license="102101600054" swrid="5190400" athleteid="47912">
              <RESULTS>
                <RESULT eventid="44384" points="483" reactiontime="+63" swimtime="00:00:37.46" resultid="47913" heatid="50702" lane="9" entrytime="00:00:37.97" entrycourse="LCM" />
                <RESULT eventid="44392" points="451" reactiontime="+59" swimtime="00:02:44.36" resultid="47914" heatid="50714" lane="4" entrytime="00:02:47.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                    <SPLIT distance="100" swimtime="00:01:17.64" />
                    <SPLIT distance="150" swimtime="00:02:05.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44409" points="486" reactiontime="+55" swimtime="00:01:21.53" resultid="47915" heatid="50754" lane="4" entrytime="00:01:23.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46304" points="474" reactiontime="+63" swimtime="00:02:58.39" resultid="47916" heatid="50842" lane="5" entrytime="00:03:04.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.45" />
                    <SPLIT distance="100" swimtime="00:01:24.97" />
                    <SPLIT distance="150" swimtime="00:02:11.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Kozik" birthdate="2006-04-19" gender="M" nation="POL" license="102101700060" swrid="5024309" athleteid="47885">
              <RESULTS>
                <RESULT eventid="44378" points="543" reactiontime="+69" swimtime="00:00:57.47" resultid="47886" heatid="50675" lane="4" entrytime="00:00:56.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="498" reactiontime="+70" swimtime="00:00:28.08" resultid="47887" heatid="50768" lane="0" entrytime="00:00:27.62" entrycourse="LCM" />
                <RESULT eventid="46298" points="556" reactiontime="+72" swimtime="00:00:25.42" resultid="47888" heatid="50821" lane="7" entrytime="00:00:25.48" entrycourse="LCM" />
                <RESULT eventid="46306" points="381" reactiontime="+70" swimtime="00:01:08.24" resultid="47889" heatid="50846" lane="4" entrytime="00:01:15.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46310" points="456" reactiontime="+69" swimtime="00:00:31.17" resultid="47890" heatid="50860" lane="8" entrytime="00:00:36.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Konrad" lastname="Pawlewicz" birthdate="2003-12-26" gender="M" nation="POL" license="102101700041" swrid="4931114" athleteid="47896">
              <RESULTS>
                <RESULT eventid="44378" points="585" reactiontime="+67" swimtime="00:00:56.07" resultid="47897" heatid="50674" lane="4" entrytime="00:00:57.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="511" reactiontime="+71" swimtime="00:00:27.85" resultid="47898" heatid="50894" lane="2" entrytime="00:00:28.69" entrycourse="LCM" />
                <RESULT eventid="46298" points="523" reactiontime="+70" swimtime="00:00:25.94" resultid="47899" heatid="50819" lane="5" entrytime="00:00:26.32" entrycourse="LCM" />
                <RESULT eventid="46306" points="430" reactiontime="+73" swimtime="00:01:05.55" resultid="47900" heatid="50847" lane="3" entrytime="00:01:09.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Musiał" birthdate="2004-09-19" gender="M" nation="POL" license="102101700044" swrid="4931089" athleteid="47891">
              <RESULTS>
                <RESULT eventid="44378" points="460" reactiontime="+64" swimtime="00:01:00.73" resultid="47892" heatid="50673" lane="3" entrytime="00:00:59.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" status="DNS" swimtime="00:00:00.00" resultid="47893" heatid="50766" lane="4" entrytime="00:00:29.17" entrycourse="LCM" />
                <RESULT eventid="46298" points="445" reactiontime="+65" swimtime="00:00:27.37" resultid="47894" heatid="50818" lane="4" entrytime="00:00:26.68" entrycourse="LCM" />
                <RESULT eventid="46310" points="395" reactiontime="+58" swimtime="00:00:32.69" resultid="47895" heatid="50860" lane="4" entrytime="00:00:32.36" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Trefler" birthdate="2004-06-11" gender="F" nation="POL" license="102101600045" swrid="4931103" athleteid="47917">
              <RESULTS>
                <RESULT eventid="44392" points="525" reactiontime="+64" swimtime="00:02:36.33" resultid="47918" heatid="50716" lane="2" entrytime="00:02:30.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                    <SPLIT distance="100" swimtime="00:01:12.56" />
                    <SPLIT distance="150" swimtime="00:01:58.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44409" points="458" reactiontime="+61" swimtime="00:01:23.14" resultid="47919" heatid="50756" lane="8" entrytime="00:01:17.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="409" reactiontime="+64" swimtime="00:00:32.89" resultid="47920" heatid="50779" lane="7" entrytime="00:00:29.88" entrycourse="LCM" />
                <RESULT eventid="46308" points="448" reactiontime="+68" swimtime="00:01:12.49" resultid="47921" heatid="50901" lane="3" entrytime="00:01:06.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Abramowicz" birthdate="2005-02-15" gender="F" nation="POL" license="102101600059" swrid="5024238" athleteid="47901">
              <RESULTS>
                <RESULT eventid="44380" points="530" reactiontime="+77" swimtime="00:01:03.87" resultid="47902" heatid="50685" lane="7" entrytime="00:01:05.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="498" reactiontime="+80" swimtime="00:00:30.81" resultid="47903" heatid="50778" lane="3" entrytime="00:00:30.94" entrycourse="LCM" />
                <RESULT eventid="46300" points="526" reactiontime="+75" swimtime="00:00:29.31" resultid="47904" heatid="50833" lane="8" entrytime="00:00:29.34" entrycourse="LCM" />
                <RESULT eventid="46308" points="516" reactiontime="+72" swimtime="00:01:09.13" resultid="47905" heatid="50900" lane="3" entrytime="00:01:10.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="95" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="F">
              <RESULTS>
                <RESULT eventid="44401" points="465" reactiontime="+67" swimtime="00:04:57.25" resultid="50888" heatid="50887" lane="3" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="100" swimtime="00:01:18.06" />
                    <SPLIT distance="150" swimtime="00:01:56.41" />
                    <SPLIT distance="200" swimtime="00:02:40.60" />
                    <SPLIT distance="250" swimtime="00:03:13.66" />
                    <SPLIT distance="300" swimtime="00:03:53.69" />
                    <SPLIT distance="350" swimtime="00:04:23.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="47906" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="47901" number="2" reactiontime="+45" />
                    <RELAYPOSITION athleteid="47912" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="47917" number="4" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="01315" nation="POL" region="15" clubid="48623" name="UPKS Wodnik Rawicz">
          <ATHLETES>
            <ATHLETE firstname="Iga" lastname="Wendzonka" birthdate="2006-10-19" gender="F" nation="POL" license="101315600290" swrid="4953340" athleteid="48664">
              <RESULTS>
                <RESULT eventid="44384" points="347" swimtime="00:00:41.83" resultid="48665" heatid="50700" lane="4" entrytime="00:00:43.37" entrycourse="LCM" />
                <RESULT eventid="44409" points="333" swimtime="00:01:32.47" resultid="48666" heatid="50753" lane="5" entrytime="00:01:35.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="386" reactiontime="+78" swimtime="00:00:37.05" resultid="48667" heatid="50907" lane="9" entrytime="00:00:37.39" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Siama" birthdate="2006-06-13" gender="F" nation="POL" license="101315600285" swrid="4952635" athleteid="48656">
              <RESULTS>
                <RESULT eventid="44380" points="375" reactiontime="+74" swimtime="00:01:11.69" resultid="48657" heatid="50681" lane="4" entrytime="00:01:12.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="343" reactiontime="+79" swimtime="00:00:34.88" resultid="48658" heatid="50775" lane="6" entrytime="00:00:35.90" entrycourse="LCM" />
                <RESULT eventid="46300" points="379" reactiontime="+77" swimtime="00:00:32.68" resultid="48659" heatid="50829" lane="6" entrytime="00:00:33.20" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Nochelska" birthdate="2007-12-03" gender="F" nation="POL" license="101315600317" swrid="4951897" athleteid="48660">
              <RESULTS>
                <RESULT eventid="44384" points="302" reactiontime="+49" swimtime="00:00:43.80" resultid="48661" heatid="50701" lane="0" entrytime="00:00:42.87" entrycourse="LCM" />
                <RESULT eventid="44409" points="296" reactiontime="+67" swimtime="00:01:36.15" resultid="48662" heatid="50753" lane="3" entrytime="00:01:35.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="344" reactiontime="+50" swimtime="00:00:33.75" resultid="48663" heatid="50827" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Maruwka" birthdate="2003-10-29" gender="M" nation="POL" license="101315700208" swrid="4938119" athleteid="48668">
              <RESULTS>
                <RESULT eventid="44390" points="579" reactiontime="+73" swimtime="00:02:16.72" resultid="48669" heatid="50711" lane="5" entrytime="00:02:12.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.61" />
                    <SPLIT distance="100" swimtime="00:01:05.08" />
                    <SPLIT distance="150" swimtime="00:01:46.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="546" reactiontime="+76" swimtime="00:02:04.74" resultid="48670" heatid="50739" lane="7" entrytime="00:01:59.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.03" />
                    <SPLIT distance="100" swimtime="00:01:01.88" />
                    <SPLIT distance="150" swimtime="00:01:34.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="519" reactiontime="+77" swimtime="00:00:27.70" resultid="48671" heatid="50769" lane="1" entrytime="00:00:25.99" entrycourse="LCM" />
                <RESULT eventid="46306" points="624" reactiontime="+70" swimtime="00:00:57.91" resultid="48672" heatid="50849" lane="4" entrytime="00:00:57.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46310" points="573" reactiontime="+64" swimtime="00:00:28.88" resultid="48673" heatid="50862" lane="8" entrytime="00:00:29.93" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominik" lastname="Boryczka" birthdate="2004-09-10" gender="M" nation="POL" license="101315700226" swrid="4988285" athleteid="48624">
              <RESULTS>
                <RESULT eventid="44378" points="583" reactiontime="+71" swimtime="00:00:56.15" resultid="48625" heatid="50676" lane="0" entrytime="00:00:55.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="511" reactiontime="+67" swimtime="00:00:32.44" resultid="48626" heatid="50694" lane="5" entrytime="00:00:33.07" entrycourse="LCM" />
                <RESULT eventid="44411" points="584" reactiontime="+72" swimtime="00:00:26.64" resultid="48627" heatid="50769" lane="0" entrytime="00:00:26.46" entrycourse="LCM" />
                <RESULT eventid="46298" points="563" reactiontime="+70" swimtime="00:00:25.32" resultid="48628" heatid="50821" lane="5" entrytime="00:00:25.07" entrycourse="LCM" />
                <RESULT eventid="46306" points="484" reactiontime="+71" swimtime="00:01:03.04" resultid="48629" heatid="50849" lane="0" entrytime="00:01:01.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jeremiasz" lastname="Marakkala Manage" birthdate="2007-02-14" gender="M" nation="POL" license="101315700306" swrid="4952507" athleteid="48630">
              <RESULTS>
                <RESULT eventid="44378" points="402" reactiontime="+77" swimtime="00:01:03.52" resultid="48631" heatid="50671" lane="4" entrytime="00:01:02.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="324" reactiontime="+74" swimtime="00:00:32.40" resultid="48632" heatid="50764" lane="6" entrytime="00:00:32.37" entrycourse="LCM" />
                <RESULT eventid="46298" status="DNS" swimtime="00:00:00.00" resultid="48633" heatid="50817" lane="9" entrytime="00:00:28.51" entrycourse="LCM" />
                <RESULT eventid="46306" status="DNS" swimtime="00:00:00.00" resultid="48634" heatid="50846" lane="1" entrytime="00:01:20.31" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Bartkowiak" birthdate="2007-05-11" gender="F" nation="POL" license="101315600347" swrid="5214799" athleteid="48649">
              <RESULTS>
                <RESULT eventid="44380" points="455" reactiontime="+71" swimtime="00:01:07.20" resultid="48650" heatid="50684" lane="2" entrytime="00:01:07.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44396" points="431" reactiontime="+78" swimtime="00:01:16.19" resultid="48651" heatid="50727" lane="0" entrytime="00:01:17.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="447" reactiontime="+58" swimtime="00:00:31.93" resultid="48652" heatid="50777" lane="4" entrytime="00:00:32.39" entrycourse="LCM" />
                <RESULT eventid="46300" points="462" reactiontime="+63" swimtime="00:00:30.60" resultid="48653" heatid="50832" lane="2" entrytime="00:00:29.92" entrycourse="LCM" />
                <RESULT eventid="46308" points="347" reactiontime="+68" swimtime="00:01:18.92" resultid="48654" heatid="50897" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="447" reactiontime="+71" swimtime="00:00:35.28" resultid="48655" heatid="50907" lane="5" entrytime="00:00:35.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Twardy" birthdate="2006-02-04" gender="M" nation="POL" license="101315700302" swrid="4951976" athleteid="48635">
              <RESULTS>
                <RESULT eventid="44378" points="409" reactiontime="+74" swimtime="00:01:03.18" resultid="48636" heatid="50671" lane="2" entrytime="00:01:02.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="395" reactiontime="+74" swimtime="00:01:10.63" resultid="48637" heatid="50722" lane="2" entrytime="00:01:10.61" entrycourse="LCM" />
                <RESULT eventid="44411" points="326" reactiontime="+71" swimtime="00:00:32.35" resultid="48638" heatid="50764" lane="7" entrytime="00:00:32.51" entrycourse="LCM" />
                <RESULT eventid="44415" points="367" reactiontime="+76" swimtime="00:02:36.18" resultid="48639" heatid="50783" lane="5" entrytime="00:02:33.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.71" />
                    <SPLIT distance="100" swimtime="00:01:18.26" />
                    <SPLIT distance="150" swimtime="00:01:58.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="385" reactiontime="+71" swimtime="00:00:28.74" resultid="48640" heatid="50816" lane="8" entrytime="00:00:29.44" entrycourse="LCM" />
                <RESULT eventid="46310" points="407" reactiontime="+67" swimtime="00:00:32.36" resultid="48641" heatid="50860" lane="3" entrytime="00:00:32.68" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alan" lastname="Szymański" birthdate="2005-06-18" gender="M" nation="POL" license="101315700255" swrid="5147691" athleteid="48642">
              <RESULTS>
                <RESULT eventid="44378" points="533" reactiontime="+67" swimtime="00:00:57.83" resultid="48643" heatid="50663" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="438" reactiontime="+66" swimtime="00:00:34.16" resultid="48644" heatid="50694" lane="7" entrytime="00:00:33.56" entrycourse="LCM" />
                <RESULT eventid="44407" points="418" reactiontime="+66" swimtime="00:01:16.07" resultid="48645" heatid="50749" lane="5" entrytime="00:01:14.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="417" reactiontime="+67" swimtime="00:00:29.79" resultid="48646" heatid="50766" lane="2" entrytime="00:00:29.57" entrycourse="LCM" />
                <RESULT eventid="46298" points="502" reactiontime="+66" swimtime="00:00:26.30" resultid="48647" heatid="50819" lane="3" entrytime="00:00:26.35" entrycourse="LCM" />
                <RESULT eventid="46310" points="391" reactiontime="+68" swimtime="00:00:32.82" resultid="48648" heatid="50861" lane="8" entrytime="00:00:32.31" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="95" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="44399" points="507" reactiontime="+72" swimtime="00:04:19.81" resultid="48674" heatid="50730" lane="3" entrytime="00:04:11.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                    <SPLIT distance="100" swimtime="00:01:09.68" />
                    <SPLIT distance="150" swimtime="00:01:44.06" />
                    <SPLIT distance="200" swimtime="00:02:25.51" />
                    <SPLIT distance="250" swimtime="00:02:52.29" />
                    <SPLIT distance="300" swimtime="00:03:24.04" />
                    <SPLIT distance="350" swimtime="00:03:50.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="48635" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="48642" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="48668" number="3" reactiontime="+19" />
                    <RELAYPOSITION athleteid="48624" number="4" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00201" nation="POL" region="01" clubid="46550" name="KS AZS AWF Wrocław">
          <ATHLETES>
            <ATHLETE firstname="Wiktor" lastname="Kopacki" birthdate="1998-02-25" gender="M" nation="POL" license="100201700093" swrid="4373332" athleteid="46555">
              <RESULTS>
                <RESULT eventid="44378" points="770" reactiontime="+69" swimtime="00:00:51.16" resultid="46556" heatid="50677" lane="5" entrytime="00:00:50.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="710" reactiontime="+72" swimtime="00:00:23.43" resultid="46557" heatid="50822" lane="5" entrytime="00:00:23.31" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Sasin" birthdate="1994-05-29" gender="F" nation="POL" license="100201600097" swrid="4236079" athleteid="46573">
              <RESULTS>
                <RESULT eventid="44380" points="601" reactiontime="+68" swimtime="00:01:01.25" resultid="46574" heatid="50688" lane="7" entrytime="00:01:00.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44392" points="526" reactiontime="+73" swimtime="00:02:36.15" resultid="46575" heatid="50712" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.94" />
                    <SPLIT distance="100" swimtime="00:01:14.96" />
                    <SPLIT distance="150" swimtime="00:02:01.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="580" reactiontime="+63" swimtime="00:00:29.28" resultid="46576" heatid="50779" lane="3" entrytime="00:00:29.08" entrycourse="LCM" />
                <RESULT eventid="46300" points="602" reactiontime="+64" swimtime="00:00:28.03" resultid="46577" heatid="50835" lane="9" entrytime="00:00:28.01" entrycourse="LCM" />
                <RESULT eventid="46308" points="554" reactiontime="+67" swimtime="00:01:07.52" resultid="46578" heatid="50901" lane="5" entrytime="00:01:05.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anatolii" lastname="Chyvylenko" birthdate="2005-11-20" gender="M" nation="POL" license="100201700202" swrid="5250942" athleteid="46567">
              <RESULTS>
                <RESULT eventid="44378" points="469" reactiontime="+66" swimtime="00:01:00.35" resultid="46568" heatid="50670" lane="5" entrytime="00:01:03.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44390" points="370" reactiontime="+68" swimtime="00:02:38.76" resultid="46569" heatid="50708" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                    <SPLIT distance="100" swimtime="00:01:15.66" />
                    <SPLIT distance="150" swimtime="00:02:01.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="388" reactiontime="+65" swimtime="00:02:19.82" resultid="46570" heatid="50736" lane="9" entrytime="00:02:20.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.41" />
                    <SPLIT distance="100" swimtime="00:01:04.62" />
                    <SPLIT distance="150" swimtime="00:01:42.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="436" reactiontime="+70" swimtime="00:00:27.57" resultid="46571" heatid="50816" lane="7" entrytime="00:00:29.23" entrycourse="LCM" />
                <RESULT eventid="46310" points="356" reactiontime="+64" swimtime="00:00:33.85" resultid="46572" heatid="50857" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Pinkosz" birthdate="1998-04-26" gender="M" nation="POL" license="100201700138" swrid="4368915" athleteid="46551">
              <RESULTS>
                <RESULT eventid="44378" points="632" reactiontime="+63" swimtime="00:00:54.64" resultid="46552" heatid="50677" lane="0" entrytime="00:00:53.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="547" reactiontime="+62" swimtime="00:00:27.22" resultid="46553" heatid="50768" lane="6" entrytime="00:00:27.13" entrycourse="LCM" />
                <RESULT eventid="46298" points="601" reactiontime="+63" swimtime="00:00:24.77" resultid="46554" heatid="50822" lane="0" entrytime="00:00:24.82" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kinga" lastname="Kołecka" birthdate="2004-12-10" gender="F" nation="POL" license="100201600184" swrid="5360593" athleteid="46579">
              <RESULTS>
                <RESULT eventid="44380" status="DNS" swimtime="00:00:00.00" resultid="46580" heatid="50680" lane="5" entrytime="00:01:18.49" entrycourse="LCM" />
                <RESULT eventid="44384" points="361" reactiontime="+83" swimtime="00:00:41.27" resultid="46581" heatid="50700" lane="5" entrytime="00:00:43.51" entrycourse="LCM" />
                <RESULT eventid="46300" points="345" reactiontime="+75" swimtime="00:00:33.72" resultid="46582" heatid="50828" lane="5" entrytime="00:00:35.14" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maksymilian" lastname="Ujec" birthdate="2004-06-29" gender="M" nation="POL" license="100201700108" swrid="5043102" athleteid="46558">
              <RESULTS>
                <RESULT eventid="44378" points="517" reactiontime="+65" swimtime="00:00:58.42" resultid="46559" heatid="50674" lane="9" entrytime="00:00:59.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44386" status="DNS" swimtime="00:00:00.00" resultid="46560" heatid="50704" lane="3" />
                <RESULT eventid="46298" points="531" reactiontime="+64" swimtime="00:00:25.81" resultid="46561" heatid="50821" lane="9" entrytime="00:00:25.85" entrycourse="LCM" />
                <RESULT eventid="46306" points="467" reactiontime="+67" swimtime="00:01:03.78" resultid="46562" heatid="50848" lane="3" entrytime="00:01:04.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" status="DNS" swimtime="00:00:00.00" resultid="50893" heatid="50757" lane="8" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roman" lastname="Domagała" birthdate="2003-04-04" gender="M" nation="POL" license="100201700194" swrid="4840761" athleteid="46563">
              <RESULTS>
                <RESULT eventid="44378" points="520" reactiontime="+61" swimtime="00:00:58.30" resultid="46564" heatid="50665" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" status="DNS" swimtime="00:00:00.00" resultid="46565" heatid="50694" lane="2" entrytime="00:00:33.36" entrycourse="LCM" />
                <RESULT eventid="46298" points="526" reactiontime="+63" swimtime="00:00:25.89" resultid="46566" heatid="50820" lane="2" entrytime="00:00:26.14" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="95" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="46289" points="611" reactiontime="+65" swimtime="00:03:41.73" resultid="46583" heatid="50794" lane="4" entrytime="00:03:33.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.75" />
                    <SPLIT distance="100" swimtime="00:00:58.93" />
                    <SPLIT distance="150" swimtime="00:01:22.90" />
                    <SPLIT distance="200" swimtime="00:01:50.02" />
                    <SPLIT distance="250" swimtime="00:02:17.28" />
                    <SPLIT distance="300" swimtime="00:02:47.72" />
                    <SPLIT distance="350" swimtime="00:03:13.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="46558" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="46555" number="2" reactiontime="+20" />
                    <RELAYPOSITION athleteid="46563" number="3" reactiontime="+28" />
                    <RELAYPOSITION athleteid="46551" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="05201" nation="POL" region="01" clubid="46594" name="KS JUST SWIM Jelenia Góra">
          <ATHLETES>
            <ATHLETE firstname="Remigiusz" lastname="Ścigała" birthdate="2007-01-04" gender="M" nation="POL" license="105201700042" swrid="4576177" athleteid="46645">
              <RESULTS>
                <RESULT eventid="44378" points="437" reactiontime="+67" swimtime="00:01:01.78" resultid="46646" heatid="50673" lane="6" entrytime="00:00:59.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="286" reactiontime="+65" swimtime="00:00:39.35" resultid="46647" heatid="50691" lane="9" />
                <RESULT eventid="44390" points="388" reactiontime="+68" swimtime="00:02:36.25" resultid="46648" heatid="50710" lane="7" entrytime="00:02:33.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                    <SPLIT distance="100" swimtime="00:01:15.08" />
                    <SPLIT distance="150" swimtime="00:02:03.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="424" reactiontime="+66" swimtime="00:02:15.77" resultid="46649" heatid="50737" lane="0" entrytime="00:02:15.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.01" />
                    <SPLIT distance="100" swimtime="00:01:05.80" />
                    <SPLIT distance="150" swimtime="00:01:41.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="352" reactiontime="+65" swimtime="00:00:31.54" resultid="46650" heatid="50765" lane="9" entrytime="00:00:31.64" entrycourse="LCM" />
                <RESULT eventid="44415" points="297" reactiontime="+74" swimtime="00:02:47.72" resultid="46651" heatid="50783" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                    <SPLIT distance="100" swimtime="00:01:22.23" />
                    <SPLIT distance="150" swimtime="00:02:06.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="459" reactiontime="+66" swimtime="00:04:45.10" resultid="46652" heatid="50799" lane="8" entrytime="00:04:54.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                    <SPLIT distance="100" swimtime="00:01:06.58" />
                    <SPLIT distance="150" swimtime="00:01:44.15" />
                    <SPLIT distance="200" swimtime="00:02:21.38" />
                    <SPLIT distance="250" swimtime="00:02:59.31" />
                    <SPLIT distance="300" swimtime="00:03:35.82" />
                    <SPLIT distance="350" swimtime="00:04:12.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="415" reactiontime="+64" swimtime="00:00:28.02" resultid="46653" heatid="50816" lane="6" entrytime="00:00:29.00" entrycourse="LCM" />
                <RESULT eventid="46306" points="307" reactiontime="+65" swimtime="00:01:13.32" resultid="46654" heatid="50847" lane="8" entrytime="00:01:12.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Nowalińska" birthdate="2006-08-01" gender="F" nation="POL" license="105201600082" swrid="5194133" athleteid="46695">
              <RESULTS>
                <RESULT eventid="44380" points="441" reactiontime="+93" swimtime="00:01:07.91" resultid="46696" heatid="50683" lane="3" entrytime="00:01:08.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44384" points="313" reactiontime="+81" swimtime="00:00:43.27" resultid="46697" heatid="50697" lane="1" />
                <RESULT eventid="44392" points="411" reactiontime="+84" swimtime="00:02:49.54" resultid="46698" heatid="50714" lane="2" entrytime="00:02:51.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.88" />
                    <SPLIT distance="100" swimtime="00:01:21.60" />
                    <SPLIT distance="150" swimtime="00:02:13.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="448" reactiontime="+71" swimtime="00:02:27.61" resultid="46699" heatid="50742" lane="0" entrytime="00:02:29.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.60" />
                    <SPLIT distance="100" swimtime="00:01:11.90" />
                    <SPLIT distance="150" swimtime="00:01:50.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="311" reactiontime="+84" swimtime="00:00:36.05" resultid="46700" heatid="50773" lane="6" entrytime="00:00:49.97" entrycourse="LCM" />
                <RESULT eventid="44417" points="404" reactiontime="+75" swimtime="00:02:46.85" resultid="46701" heatid="50786" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.89" />
                    <SPLIT distance="100" swimtime="00:01:21.75" />
                    <SPLIT distance="150" swimtime="00:02:05.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="482" reactiontime="+82" swimtime="00:05:01.44" resultid="46702" heatid="50803" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.65" />
                    <SPLIT distance="100" swimtime="00:01:11.65" />
                    <SPLIT distance="150" swimtime="00:01:51.28" />
                    <SPLIT distance="200" swimtime="00:02:30.10" />
                    <SPLIT distance="250" swimtime="00:03:09.02" />
                    <SPLIT distance="300" swimtime="00:03:47.79" />
                    <SPLIT distance="350" swimtime="00:04:26.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="426" reactiontime="+78" swimtime="00:00:31.45" resultid="46703" heatid="50827" lane="7" />
                <RESULT eventid="46308" points="268" reactiontime="+61" swimtime="00:01:25.97" resultid="46704" heatid="50898" lane="4" entrytime="00:01:22.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Bancewicz" birthdate="2006-10-31" gender="M" nation="POL" license="105201700030" swrid="5190367" athleteid="46595">
              <RESULTS>
                <RESULT eventid="44378" points="363" reactiontime="+72" swimtime="00:01:05.72" resultid="46596" heatid="50667" lane="9" entrytime="00:01:13.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="223" reactiontime="+80" swimtime="00:00:42.77" resultid="46597" heatid="50690" lane="6" />
                <RESULT eventid="44390" points="298" swimtime="00:02:50.60" resultid="46598" heatid="50708" lane="4" entrytime="00:03:05.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                    <SPLIT distance="100" swimtime="00:01:22.19" />
                    <SPLIT distance="150" swimtime="00:02:13.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="328" reactiontime="+79" swimtime="00:02:27.90" resultid="46599" heatid="50734" lane="3" entrytime="00:02:30.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.01" />
                    <SPLIT distance="100" swimtime="00:01:12.13" />
                    <SPLIT distance="150" swimtime="00:01:50.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="272" reactiontime="+77" swimtime="00:00:34.33" resultid="46600" heatid="50761" lane="8" />
                <RESULT eventid="44415" points="273" reactiontime="+70" swimtime="00:02:52.37" resultid="46601" heatid="50782" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.69" />
                    <SPLIT distance="100" swimtime="00:01:24.46" />
                    <SPLIT distance="150" swimtime="00:02:09.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="319" reactiontime="+75" swimtime="00:05:21.90" resultid="46602" heatid="50797" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                    <SPLIT distance="100" swimtime="00:01:13.13" />
                    <SPLIT distance="150" swimtime="00:01:54.38" />
                    <SPLIT distance="200" swimtime="00:02:36.58" />
                    <SPLIT distance="250" swimtime="00:03:18.87" />
                    <SPLIT distance="300" swimtime="00:04:01.45" />
                    <SPLIT distance="350" swimtime="00:04:43.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="359" reactiontime="+76" swimtime="00:00:29.42" resultid="46603" heatid="50814" lane="0" entrytime="00:00:32.72" entrycourse="LCM" />
                <RESULT eventid="46306" points="208" reactiontime="+79" swimtime="00:01:23.53" resultid="46604" heatid="50844" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Niedzielska" birthdate="2006-04-12" gender="F" nation="POL" license="105201600056" swrid="5081136" athleteid="46675">
              <RESULTS>
                <RESULT eventid="44380" points="384" reactiontime="+68" swimtime="00:01:11.09" resultid="46676" heatid="50682" lane="8" entrytime="00:01:11.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44384" points="257" reactiontime="+69" swimtime="00:00:46.22" resultid="46677" heatid="50698" lane="1" />
                <RESULT eventid="44392" points="313" reactiontime="+68" swimtime="00:03:05.73" resultid="46678" heatid="50713" lane="3" entrytime="00:03:02.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.45" />
                    <SPLIT distance="100" swimtime="00:01:26.49" />
                    <SPLIT distance="150" swimtime="00:02:24.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="349" reactiontime="+65" swimtime="00:02:40.44" resultid="46679" heatid="50740" lane="2" entrytime="00:02:42.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.66" />
                    <SPLIT distance="100" swimtime="00:01:17.57" />
                    <SPLIT distance="150" swimtime="00:02:00.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="269" reactiontime="+54" swimtime="00:00:37.83" resultid="46680" heatid="50774" lane="0" entrytime="00:00:41.40" entrycourse="LCM" />
                <RESULT eventid="44417" points="308" reactiontime="+83" swimtime="00:03:02.62" resultid="46681" heatid="50786" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.19" />
                    <SPLIT distance="100" swimtime="00:01:28.63" />
                    <SPLIT distance="150" swimtime="00:02:17.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="351" reactiontime="+45" swimtime="00:05:34.94" resultid="46682" heatid="50801" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.91" />
                    <SPLIT distance="100" swimtime="00:01:17.19" />
                    <SPLIT distance="150" swimtime="00:02:00.14" />
                    <SPLIT distance="200" swimtime="00:02:43.53" />
                    <SPLIT distance="250" swimtime="00:03:27.51" />
                    <SPLIT distance="300" swimtime="00:04:11.37" />
                    <SPLIT distance="350" swimtime="00:04:54.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="376" reactiontime="+69" swimtime="00:00:32.78" resultid="46683" heatid="50825" lane="3" />
                <RESULT eventid="46308" points="249" reactiontime="+67" swimtime="00:01:28.09" resultid="46684" heatid="50898" lane="6" entrytime="00:01:26.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krystian" lastname="Kasprzak" birthdate="2007-05-05" gender="M" nation="POL" license="105201700035" swrid="5190366" athleteid="46625">
              <RESULTS>
                <RESULT eventid="44378" points="362" reactiontime="+65" swimtime="00:01:05.77" resultid="46626" heatid="50669" lane="2" entrytime="00:01:05.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="237" reactiontime="+65" swimtime="00:00:41.90" resultid="46627" heatid="50690" lane="7" />
                <RESULT eventid="44390" points="352" reactiontime="+54" swimtime="00:02:41.42" resultid="46628" heatid="50709" lane="5" entrytime="00:02:44.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                    <SPLIT distance="100" swimtime="00:01:16.83" />
                    <SPLIT distance="150" swimtime="00:02:04.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="354" reactiontime="+64" swimtime="00:02:24.08" resultid="46629" heatid="50735" lane="2" entrytime="00:02:25.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                    <SPLIT distance="100" swimtime="00:01:09.73" />
                    <SPLIT distance="150" swimtime="00:01:48.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="319" reactiontime="+54" swimtime="00:00:32.57" resultid="46630" heatid="50764" lane="0" entrytime="00:00:32.76" entrycourse="LCM" />
                <RESULT eventid="44415" points="301" reactiontime="+76" swimtime="00:02:46.86" resultid="46631" heatid="50782" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.83" />
                    <SPLIT distance="100" swimtime="00:01:22.31" />
                    <SPLIT distance="150" swimtime="00:02:05.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="374" reactiontime="+64" swimtime="00:05:05.19" resultid="46632" heatid="50798" lane="3" entrytime="00:05:14.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                    <SPLIT distance="100" swimtime="00:01:10.63" />
                    <SPLIT distance="150" swimtime="00:01:50.31" />
                    <SPLIT distance="200" swimtime="00:02:30.67" />
                    <SPLIT distance="250" swimtime="00:03:10.56" />
                    <SPLIT distance="300" swimtime="00:03:50.92" />
                    <SPLIT distance="350" swimtime="00:04:29.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="355" reactiontime="+47" swimtime="00:00:29.53" resultid="46633" heatid="50815" lane="2" entrytime="00:00:30.06" entrycourse="LCM" />
                <RESULT eventid="46306" points="265" reactiontime="+71" swimtime="00:01:16.98" resultid="46634" heatid="50846" lane="3" entrytime="00:01:17.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Niedzielska" birthdate="2007-12-12" gender="F" nation="POL" license="105201600057" swrid="5108628" athleteid="46685">
              <RESULTS>
                <RESULT eventid="44380" points="280" swimtime="00:01:19.00" resultid="46686" heatid="50681" lane="0" entrytime="00:01:17.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44384" status="DNS" swimtime="00:00:00.00" resultid="46687" heatid="50697" lane="4" />
                <RESULT eventid="44392" points="305" reactiontime="+76" swimtime="00:03:07.19" resultid="46688" heatid="50713" lane="7" entrytime="00:03:07.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.09" />
                    <SPLIT distance="100" swimtime="00:01:31.16" />
                    <SPLIT distance="150" swimtime="00:02:27.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="292" reactiontime="+57" swimtime="00:02:50.15" resultid="46689" heatid="50740" lane="1" entrytime="00:02:50.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                    <SPLIT distance="100" swimtime="00:01:23.39" />
                    <SPLIT distance="150" swimtime="00:02:07.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="187" reactiontime="+65" swimtime="00:00:42.69" resultid="46690" heatid="50773" lane="2" entrytime="00:00:53.76" entrycourse="LCM" />
                <RESULT eventid="44417" points="302" reactiontime="+85" swimtime="00:03:03.75" resultid="46691" heatid="50786" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.79" />
                    <SPLIT distance="100" swimtime="00:01:31.45" />
                    <SPLIT distance="150" swimtime="00:02:19.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="313" swimtime="00:05:48.10" resultid="46692" heatid="50804" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                    <SPLIT distance="100" swimtime="00:01:19.83" />
                    <SPLIT distance="150" swimtime="00:02:04.72" />
                    <SPLIT distance="200" swimtime="00:02:50.40" />
                    <SPLIT distance="250" swimtime="00:03:36.91" />
                    <SPLIT distance="300" swimtime="00:04:22.09" />
                    <SPLIT distance="350" swimtime="00:05:06.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="315" reactiontime="+68" swimtime="00:00:34.76" resultid="46693" heatid="50824" lane="8" />
                <RESULT eventid="46308" points="168" reactiontime="+55" swimtime="00:01:40.36" resultid="46694" heatid="50898" lane="9" entrytime="00:01:40.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amelia" lastname="Choroszy" birthdate="2008-04-18" gender="F" nation="POL" license="105201600058" swrid="4574174" athleteid="46705">
              <RESULTS>
                <RESULT eventid="44380" points="427" reactiontime="+87" swimtime="00:01:08.63" resultid="46706" heatid="50683" lane="2" entrytime="00:01:08.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44384" points="405" reactiontime="+66" swimtime="00:00:39.73" resultid="46707" heatid="50701" lane="9" entrytime="00:00:42.95" entrycourse="LCM" />
                <RESULT eventid="44392" points="377" reactiontime="+80" swimtime="00:02:54.58" resultid="46708" heatid="50714" lane="8" entrytime="00:02:52.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.35" />
                    <SPLIT distance="100" swimtime="00:01:25.79" />
                    <SPLIT distance="150" swimtime="00:02:15.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="383" reactiontime="+78" swimtime="00:02:35.54" resultid="46709" heatid="50741" lane="1" entrytime="00:02:35.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                    <SPLIT distance="100" swimtime="00:01:16.45" />
                    <SPLIT distance="150" swimtime="00:01:57.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="342" reactiontime="+83" swimtime="00:00:34.91" resultid="46710" heatid="50776" lane="8" entrytime="00:00:34.94" entrycourse="LCM" />
                <RESULT eventid="44417" points="361" reactiontime="+78" swimtime="00:02:53.11" resultid="46711" heatid="50785" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.41" />
                    <SPLIT distance="100" swimtime="00:01:26.17" />
                    <SPLIT distance="150" swimtime="00:02:11.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="383" reactiontime="+73" swimtime="00:05:25.54" resultid="46712" heatid="50803" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                    <SPLIT distance="100" swimtime="00:01:17.31" />
                    <SPLIT distance="150" swimtime="00:01:59.41" />
                    <SPLIT distance="200" swimtime="00:02:41.52" />
                    <SPLIT distance="250" swimtime="00:03:23.85" />
                    <SPLIT distance="300" swimtime="00:04:05.59" />
                    <SPLIT distance="350" swimtime="00:04:46.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="466" reactiontime="+77" swimtime="00:00:30.51" resultid="46713" heatid="50830" lane="2" entrytime="00:00:31.67" entrycourse="LCM" />
                <RESULT eventid="46308" points="248" reactiontime="+81" swimtime="00:01:28.27" resultid="46714" heatid="50898" lane="1" entrytime="00:01:28.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksander" lastname="Binasiewicz" birthdate="2006-05-03" gender="M" nation="POL" license="105201700061" swrid="4995364" athleteid="46615">
              <RESULTS>
                <RESULT eventid="44378" points="264" reactiontime="+72" swimtime="00:01:13.05" resultid="46616" heatid="50667" lane="7" entrytime="00:01:10.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="185" reactiontime="+60" swimtime="00:00:45.50" resultid="46617" heatid="50691" lane="4" />
                <RESULT eventid="44390" points="224" reactiontime="+81" swimtime="00:03:07.68" resultid="46618" heatid="50709" lane="0" entrytime="00:02:55.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.38" />
                    <SPLIT distance="100" swimtime="00:01:30.24" />
                    <SPLIT distance="150" swimtime="00:02:27.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="243" reactiontime="+71" swimtime="00:02:43.39" resultid="46619" heatid="50734" lane="8" entrytime="00:02:32.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.82" />
                    <SPLIT distance="100" swimtime="00:01:18.68" />
                    <SPLIT distance="150" swimtime="00:02:02.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="252" reactiontime="+75" swimtime="00:00:35.24" resultid="46620" heatid="50757" lane="6" />
                <RESULT eventid="44415" points="201" reactiontime="+96" swimtime="00:03:10.91" resultid="46621" heatid="50782" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.21" />
                    <SPLIT distance="100" swimtime="00:01:34.24" />
                    <SPLIT distance="150" swimtime="00:02:23.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="300" reactiontime="+69" swimtime="00:05:28.53" resultid="46622" heatid="50797" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                    <SPLIT distance="100" swimtime="00:01:17.28" />
                    <SPLIT distance="150" swimtime="00:01:59.01" />
                    <SPLIT distance="200" swimtime="00:02:42.03" />
                    <SPLIT distance="250" swimtime="00:03:24.51" />
                    <SPLIT distance="300" swimtime="00:04:07.50" />
                    <SPLIT distance="350" swimtime="00:04:49.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="275" reactiontime="+75" swimtime="00:00:32.15" resultid="46623" heatid="50810" lane="7" />
                <RESULT eventid="46306" points="205" reactiontime="+64" swimtime="00:01:23.92" resultid="46624" heatid="50845" lane="5" entrytime="00:01:24.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hubert" lastname="Skowron" birthdate="2006-05-25" gender="M" nation="POL" license="105201700039" swrid="5210843" athleteid="46635">
              <RESULTS>
                <RESULT eventid="44378" points="416" reactiontime="+83" swimtime="00:01:02.80" resultid="46636" heatid="50672" lane="1" entrytime="00:01:01.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="295" reactiontime="+85" swimtime="00:00:38.97" resultid="46637" heatid="50689" lane="6" />
                <RESULT eventid="44390" points="387" reactiontime="+82" swimtime="00:02:36.36" resultid="46638" heatid="50710" lane="1" entrytime="00:02:34.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                    <SPLIT distance="100" swimtime="00:01:15.78" />
                    <SPLIT distance="150" swimtime="00:02:01.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="419" reactiontime="+74" swimtime="00:02:16.26" resultid="46639" heatid="50736" lane="0" entrytime="00:02:20.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                    <SPLIT distance="100" swimtime="00:01:06.27" />
                    <SPLIT distance="150" swimtime="00:01:42.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="310" reactiontime="+76" swimtime="00:00:32.90" resultid="46640" heatid="50764" lane="1" entrytime="00:00:32.54" entrycourse="LCM" />
                <RESULT eventid="44415" points="324" reactiontime="+89" swimtime="00:02:42.88" resultid="46641" heatid="50782" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.85" />
                    <SPLIT distance="100" swimtime="00:01:20.49" />
                    <SPLIT distance="150" swimtime="00:02:02.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="451" reactiontime="+75" swimtime="00:04:46.92" resultid="46642" heatid="50799" lane="9" entrytime="00:05:01.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.55" />
                    <SPLIT distance="100" swimtime="00:01:07.19" />
                    <SPLIT distance="150" swimtime="00:01:44.77" />
                    <SPLIT distance="200" swimtime="00:02:22.33" />
                    <SPLIT distance="250" swimtime="00:02:59.83" />
                    <SPLIT distance="300" swimtime="00:03:36.33" />
                    <SPLIT distance="350" swimtime="00:04:12.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="381" reactiontime="+75" swimtime="00:00:28.83" resultid="46643" heatid="50816" lane="3" entrytime="00:00:28.87" entrycourse="LCM" />
                <RESULT eventid="46306" points="301" reactiontime="+80" swimtime="00:01:13.83" resultid="46644" heatid="50847" lane="1" entrytime="00:01:12.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwier" lastname="Barczyński" birthdate="2006-09-21" gender="M" nation="POL" license="105201700029" swrid="5194169" athleteid="46605">
              <RESULTS>
                <RESULT eventid="44378" points="381" reactiontime="+66" swimtime="00:01:04.68" resultid="46606" heatid="50669" lane="1" entrytime="00:01:05.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="203" reactiontime="+63" swimtime="00:00:44.13" resultid="46607" heatid="50691" lane="5" />
                <RESULT eventid="44390" points="318" reactiontime="+67" swimtime="00:02:46.86" resultid="46608" heatid="50709" lane="2" entrytime="00:02:47.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                    <SPLIT distance="100" swimtime="00:01:16.40" />
                    <SPLIT distance="150" swimtime="00:02:10.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="355" reactiontime="+66" swimtime="00:02:24.05" resultid="46609" heatid="50735" lane="1" entrytime="00:02:25.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.53" />
                    <SPLIT distance="100" swimtime="00:01:08.77" />
                    <SPLIT distance="150" swimtime="00:01:47.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="313" reactiontime="+51" swimtime="00:00:32.77" resultid="46610" heatid="50758" lane="9" />
                <RESULT eventid="44415" points="282" reactiontime="+53" swimtime="00:02:50.65" resultid="46611" heatid="50783" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.22" />
                    <SPLIT distance="100" swimtime="00:01:23.54" />
                    <SPLIT distance="150" swimtime="00:02:08.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="352" reactiontime="+69" swimtime="00:05:11.52" resultid="46612" heatid="50797" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                    <SPLIT distance="100" swimtime="00:01:10.91" />
                    <SPLIT distance="150" swimtime="00:01:51.12" />
                    <SPLIT distance="200" swimtime="00:02:31.58" />
                    <SPLIT distance="250" swimtime="00:03:12.15" />
                    <SPLIT distance="300" swimtime="00:03:53.16" />
                    <SPLIT distance="350" swimtime="00:04:33.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="342" reactiontime="+65" swimtime="00:00:29.90" resultid="46613" heatid="50813" lane="3" entrytime="00:00:33.10" entrycourse="LCM" />
                <RESULT eventid="46306" points="187" reactiontime="+65" swimtime="00:01:26.42" resultid="46614" heatid="50846" lane="9" entrytime="00:01:22.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Książek" birthdate="2005-02-23" gender="F" nation="POL" license="105201600022" swrid="4012868" athleteid="46665">
              <RESULTS>
                <RESULT eventid="44380" points="567" reactiontime="+73" swimtime="00:01:02.45" resultid="46666" heatid="50687" lane="1" entrytime="00:01:02.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44384" points="358" reactiontime="+67" swimtime="00:00:41.38" resultid="46667" heatid="50699" lane="2" />
                <RESULT eventid="44392" points="505" reactiontime="+80" swimtime="00:02:38.37" resultid="46668" heatid="50715" lane="6" entrytime="00:02:40.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                    <SPLIT distance="100" swimtime="00:01:14.36" />
                    <SPLIT distance="150" swimtime="00:02:03.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="529" reactiontime="+66" swimtime="00:02:19.64" resultid="46669" heatid="50743" lane="0" entrytime="00:02:20.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                    <SPLIT distance="100" swimtime="00:01:07.48" />
                    <SPLIT distance="150" swimtime="00:01:44.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="452" reactiontime="+76" swimtime="00:00:31.81" resultid="46670" heatid="50778" lane="8" entrytime="00:00:32.08" entrycourse="LCM" />
                <RESULT eventid="44417" points="410" reactiontime="+73" swimtime="00:02:45.95" resultid="46671" heatid="50785" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.52" />
                    <SPLIT distance="100" swimtime="00:01:21.21" />
                    <SPLIT distance="150" swimtime="00:02:04.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="500" swimtime="00:04:57.76" resultid="46672" heatid="50804" lane="4" entrytime="00:04:56.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.29" />
                    <SPLIT distance="100" swimtime="00:01:07.90" />
                    <SPLIT distance="150" swimtime="00:01:46.59" />
                    <SPLIT distance="200" swimtime="00:02:25.66" />
                    <SPLIT distance="250" swimtime="00:03:04.78" />
                    <SPLIT distance="300" swimtime="00:03:43.49" />
                    <SPLIT distance="350" swimtime="00:04:22.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="551" reactiontime="+75" swimtime="00:00:28.86" resultid="46673" heatid="50833" lane="1" entrytime="00:00:29.30" entrycourse="LCM" />
                <RESULT eventid="46308" points="404" reactiontime="+70" swimtime="00:01:15.02" resultid="46674" heatid="50899" lane="2" entrytime="00:01:18.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Gołębiewska" birthdate="2006-11-03" gender="F" nation="POL" license="105201600041" swrid="5081130" athleteid="46655">
              <RESULTS>
                <RESULT eventid="44380" points="305" reactiontime="+73" swimtime="00:01:16.76" resultid="46656" heatid="50681" lane="6" entrytime="00:01:15.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44384" status="DNS" swimtime="00:00:00.00" resultid="46657" heatid="50697" lane="8" />
                <RESULT eventid="44392" points="304" reactiontime="+75" swimtime="00:03:07.51" resultid="46658" heatid="50713" lane="6" entrytime="00:03:05.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.69" />
                    <SPLIT distance="100" swimtime="00:01:33.24" />
                    <SPLIT distance="150" swimtime="00:02:28.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="328" reactiontime="+76" swimtime="00:02:43.75" resultid="46659" heatid="50740" lane="6" entrytime="00:02:40.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.37" />
                    <SPLIT distance="100" swimtime="00:01:19.29" />
                    <SPLIT distance="150" swimtime="00:02:02.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="184" reactiontime="+77" swimtime="00:00:42.91" resultid="46660" heatid="50772" lane="6" />
                <RESULT eventid="44417" points="293" reactiontime="+75" swimtime="00:03:05.63" resultid="46661" heatid="50785" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.51" />
                    <SPLIT distance="100" swimtime="00:01:30.87" />
                    <SPLIT distance="150" swimtime="00:02:19.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="332" reactiontime="+74" swimtime="00:05:41.37" resultid="46662" heatid="50802" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.91" />
                    <SPLIT distance="100" swimtime="00:01:19.37" />
                    <SPLIT distance="150" swimtime="00:02:03.75" />
                    <SPLIT distance="200" swimtime="00:02:48.09" />
                    <SPLIT distance="250" swimtime="00:03:32.68" />
                    <SPLIT distance="300" swimtime="00:04:16.30" />
                    <SPLIT distance="350" swimtime="00:05:00.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="307" reactiontime="+69" swimtime="00:00:35.08" resultid="46663" heatid="50828" lane="1" entrytime="00:00:38.47" entrycourse="LCM" />
                <RESULT eventid="46308" points="177" reactiontime="+68" swimtime="00:01:38.65" resultid="46664" heatid="50898" lane="0" entrytime="00:01:37.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00801" nation="POL" region="01" clubid="47645" name="MKS Płetval Polkowice">
          <ATHLETES>
            <ATHLETE firstname="Bruno" lastname="Cios" birthdate="2007-11-28" gender="M" nation="POL" license="100801700017" swrid="5272062" athleteid="47646">
              <RESULTS>
                <RESULT eventid="46298" points="376" reactiontime="+78" swimtime="00:00:28.97" resultid="47647" heatid="50814" lane="6" entrytime="00:00:32.01" entrycourse="LCM" />
                <RESULT eventid="46306" points="196" reactiontime="+78" swimtime="00:01:25.14" resultid="47648" heatid="50846" lane="2" entrytime="00:01:18.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Zieliński" birthdate="2005-11-18" gender="M" nation="POL" license="100801700018" swrid="5043110" athleteid="47649">
              <RESULTS>
                <RESULT eventid="46298" points="463" reactiontime="+72" swimtime="00:00:27.02" resultid="47650" heatid="50816" lane="1" entrytime="00:00:29.32" entrycourse="LCM" />
                <RESULT eventid="46306" points="463" reactiontime="+74" swimtime="00:01:03.97" resultid="47651" heatid="50848" lane="6" entrytime="00:01:05.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06215" nation="POL" region="15" clubid="47823" name="UKS &quot;Dwójka&quot; w Obornikach">
          <ATHLETES>
            <ATHLETE firstname="Angelika" lastname="Bluge" birthdate="2000-03-20" gender="F" nation="POL" license="106215600042" swrid="4647713" athleteid="47824">
              <RESULTS>
                <RESULT eventid="44384" points="565" reactiontime="+74" swimtime="00:00:35.56" resultid="47825" heatid="50703" lane="8" entrytime="00:00:34.87" entrycourse="LCM" />
                <RESULT eventid="44409" points="479" reactiontime="+69" swimtime="00:01:21.95" resultid="47826" heatid="50756" lane="0" entrytime="00:01:18.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46304" points="497" reactiontime="+71" swimtime="00:02:55.60" resultid="47827" heatid="50843" lane="6" entrytime="00:02:47.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.94" />
                    <SPLIT distance="100" swimtime="00:01:23.25" />
                    <SPLIT distance="150" swimtime="00:02:09.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="05501" nation="POL" region="01" clubid="47922" name="UKS ,,HS&apos;&apos; Team Kryty Basen Kłodzko">
          <ATHLETES>
            <ATHLETE firstname="Cyprian" lastname="Liszka" birthdate="2007-02-18" gender="M" nation="POL" license="105501700036" swrid="5136362" athleteid="47923">
              <RESULTS>
                <RESULT eventid="44378" points="353" reactiontime="+70" swimtime="00:01:06.36" resultid="47924" heatid="50669" lane="5" entrytime="00:01:05.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="310" reactiontime="+69" swimtime="00:01:16.54" resultid="47925" heatid="50720" lane="5" entrytime="00:01:17.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" status="DNS" swimtime="00:00:00.00" resultid="47926" heatid="50760" lane="9" />
                <RESULT eventid="46298" points="391" reactiontime="+70" swimtime="00:00:28.59" resultid="47927" heatid="50811" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Poręba" birthdate="2007-09-12" gender="F" nation="POL" license="105501600006" swrid="5210814" athleteid="47937">
              <RESULTS>
                <RESULT eventid="44384" points="643" reactiontime="+66" swimtime="00:00:34.06" resultid="47938" heatid="50703" lane="1" entrytime="00:00:34.70" entrycourse="LCM" />
                <RESULT eventid="44392" points="535" reactiontime="+58" swimtime="00:02:35.35" resultid="47939" heatid="50715" lane="4" entrytime="00:02:34.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:15.89" />
                    <SPLIT distance="150" swimtime="00:01:58.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44409" points="596" reactiontime="+67" swimtime="00:01:16.19" resultid="47940" heatid="50755" lane="6" entrytime="00:01:19.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46304" points="582" reactiontime="+70" swimtime="00:02:46.61" resultid="47941" heatid="50842" lane="2" entrytime="00:03:09.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                    <SPLIT distance="100" swimtime="00:01:19.58" />
                    <SPLIT distance="150" swimtime="00:02:03.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Wierzbicka" birthdate="2007-08-04" gender="F" nation="POL" license="105501600020" swrid="5166030" athleteid="47932">
              <RESULTS>
                <RESULT eventid="44380" points="505" reactiontime="+74" swimtime="00:01:04.90" resultid="47933" heatid="50684" lane="6" entrytime="00:01:06.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="460" reactiontime="+74" swimtime="00:00:31.64" resultid="47934" heatid="50775" lane="8" entrytime="00:00:37.64" entrycourse="LCM" />
                <RESULT eventid="46308" points="467" reactiontime="+68" swimtime="00:01:11.50" resultid="47935" heatid="50900" lane="6" entrytime="00:01:11.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="482" reactiontime="+59" swimtime="00:00:34.40" resultid="47936" heatid="50905" lane="4" entrytime="00:00:42.12" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pascal" lastname="Blacheta" birthdate="2004-12-24" gender="M" nation="POL" license="105501700001" swrid="5118756" athleteid="47928">
              <RESULTS>
                <RESULT eventid="44378" points="521" reactiontime="+78" swimtime="00:00:58.27" resultid="47929" heatid="50668" lane="4" entrytime="00:01:06.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="431" reactiontime="+81" swimtime="00:01:08.60" resultid="47930" heatid="50721" lane="5" entrytime="00:01:14.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="433" reactiontime="+79" swimtime="00:02:27.93" resultid="47931" heatid="50783" lane="7" entrytime="00:02:43.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                    <SPLIT distance="100" swimtime="00:01:13.43" />
                    <SPLIT distance="150" swimtime="00:01:51.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hanna" lastname="Lewicka" birthdate="2007-07-26" gender="F" nation="POL" license="105501600009" swrid="5210829" athleteid="47952">
              <RESULTS>
                <RESULT eventid="44396" points="441" reactiontime="+63" swimtime="00:01:15.62" resultid="47953" heatid="50726" lane="6" entrytime="00:01:18.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44417" points="445" reactiontime="+73" swimtime="00:02:41.46" resultid="47954" heatid="50786" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.28" />
                    <SPLIT distance="100" swimtime="00:01:19.42" />
                    <SPLIT distance="150" swimtime="00:02:00.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="371" reactiontime="+72" swimtime="00:05:28.95" resultid="47955" heatid="50802" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.60" />
                    <SPLIT distance="100" swimtime="00:01:15.95" />
                    <SPLIT distance="150" swimtime="00:01:57.67" />
                    <SPLIT distance="200" swimtime="00:02:40.68" />
                    <SPLIT distance="250" swimtime="00:03:23.47" />
                    <SPLIT distance="300" swimtime="00:04:06.47" />
                    <SPLIT distance="350" swimtime="00:04:48.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="416" reactiontime="+81" swimtime="00:00:36.14" resultid="47956" heatid="50905" lane="3" entrytime="00:00:43.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zofia" lastname="Chilarska" birthdate="2008-07-09" gender="F" nation="POL" license="105501600035" swrid="5204354" athleteid="47942">
              <RESULTS>
                <RESULT eventid="44384" points="437" reactiontime="+61" swimtime="00:00:38.74" resultid="47943" heatid="50700" lane="2" entrytime="00:00:44.60" entrycourse="LCM" />
                <RESULT eventid="44409" points="419" reactiontime="+68" swimtime="00:01:25.64" resultid="47944" heatid="50754" lane="8" entrytime="00:01:29.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="372" reactiontime="+58" swimtime="00:00:33.95" resultid="47945" heatid="50777" lane="9" entrytime="00:00:33.55" entrycourse="LCM" />
                <RESULT eventid="46304" points="404" reactiontime="+65" swimtime="00:03:08.11" resultid="47946" heatid="50841" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.55" />
                    <SPLIT distance="100" swimtime="00:01:29.83" />
                    <SPLIT distance="150" swimtime="00:02:19.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zofia" lastname="Porębska" birthdate="2008-01-20" gender="F" nation="POL" license="105501600031" swrid="5001940" athleteid="47947">
              <RESULTS>
                <RESULT eventid="44384" points="325" reactiontime="+80" swimtime="00:00:42.75" resultid="47948" heatid="50700" lane="6" entrytime="00:00:43.87" entrycourse="LCM" />
                <RESULT eventid="44396" points="308" reactiontime="+87" swimtime="00:01:25.21" resultid="47949" heatid="50725" lane="5" entrytime="00:01:24.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44409" points="329" swimtime="00:01:32.88" resultid="47950" heatid="50753" lane="4" entrytime="00:01:34.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46304" points="362" reactiontime="+77" swimtime="00:03:15.11" resultid="47951" heatid="50841" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.39" />
                    <SPLIT distance="100" swimtime="00:01:32.52" />
                    <SPLIT distance="150" swimtime="00:02:23.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01006" nation="POL" region="06" clubid="47818" name="UKP Unia Oświęcim">
          <ATHLETES>
            <ATHLETE firstname="Karol" lastname="Cembala" birthdate="2005-07-31" gender="M" nation="POL" license="101006700460" swrid="5043014" athleteid="47819">
              <RESULTS>
                <RESULT eventid="44378" points="442" reactiontime="+75" swimtime="00:01:01.56" resultid="47820" heatid="50671" lane="0" entrytime="00:01:03.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="489" reactiontime="+77" swimtime="00:02:09.40" resultid="47821" heatid="50737" lane="1" entrytime="00:02:14.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.29" />
                    <SPLIT distance="100" swimtime="00:01:02.25" />
                    <SPLIT distance="150" swimtime="00:01:35.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="534" reactiontime="+76" swimtime="00:04:31.09" resultid="47822" heatid="50800" lane="0" entrytime="00:04:37.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.94" />
                    <SPLIT distance="100" swimtime="00:01:04.48" />
                    <SPLIT distance="150" swimtime="00:01:38.39" />
                    <SPLIT distance="200" swimtime="00:02:13.84" />
                    <SPLIT distance="250" swimtime="00:02:47.38" />
                    <SPLIT distance="300" swimtime="00:03:22.41" />
                    <SPLIT distance="350" swimtime="00:03:57.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00116" nation="POL" region="16" clubid="47078" name="MKP Szczecin">
          <ATHLETES>
            <ATHLETE firstname="Nikodem" lastname="Wieczorkowski" birthdate="2004-04-21" gender="M" nation="POL" license="100116701340" swrid="5011793" athleteid="47083">
              <RESULTS>
                <RESULT eventid="44378" points="513" reactiontime="+67" swimtime="00:00:58.58" resultid="47084" heatid="50675" lane="8" entrytime="00:00:57.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46285" points="603" reactiontime="+63" swimtime="00:17:10.98" resultid="47085" heatid="50790" lane="4" entrytime="00:16:54.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                    <SPLIT distance="100" swimtime="00:01:04.48" />
                    <SPLIT distance="150" swimtime="00:01:38.00" />
                    <SPLIT distance="200" swimtime="00:02:11.51" />
                    <SPLIT distance="250" swimtime="00:02:44.92" />
                    <SPLIT distance="300" swimtime="00:03:18.59" />
                    <SPLIT distance="350" swimtime="00:03:51.85" />
                    <SPLIT distance="400" swimtime="00:04:25.58" />
                    <SPLIT distance="450" swimtime="00:04:59.15" />
                    <SPLIT distance="500" swimtime="00:05:33.03" />
                    <SPLIT distance="550" swimtime="00:06:07.21" />
                    <SPLIT distance="600" swimtime="00:06:41.78" />
                    <SPLIT distance="650" swimtime="00:07:16.41" />
                    <SPLIT distance="700" swimtime="00:07:51.06" />
                    <SPLIT distance="750" swimtime="00:08:25.64" />
                    <SPLIT distance="800" swimtime="00:09:01.28" />
                    <SPLIT distance="850" swimtime="00:09:36.05" />
                    <SPLIT distance="900" swimtime="00:10:11.18" />
                    <SPLIT distance="950" swimtime="00:10:46.52" />
                    <SPLIT distance="1000" swimtime="00:11:21.55" />
                    <SPLIT distance="1050" swimtime="00:11:56.74" />
                    <SPLIT distance="1100" swimtime="00:12:31.88" />
                    <SPLIT distance="1150" swimtime="00:13:07.11" />
                    <SPLIT distance="1200" swimtime="00:13:42.83" />
                    <SPLIT distance="1250" swimtime="00:14:18.04" />
                    <SPLIT distance="1300" swimtime="00:14:53.42" />
                    <SPLIT distance="1350" swimtime="00:15:28.65" />
                    <SPLIT distance="1400" swimtime="00:16:03.87" />
                    <SPLIT distance="1450" swimtime="00:16:38.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="578" reactiontime="+70" swimtime="00:04:24.15" resultid="47086" heatid="50800" lane="3" entrytime="00:04:17.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.74" />
                    <SPLIT distance="100" swimtime="00:01:01.34" />
                    <SPLIT distance="150" swimtime="00:01:34.76" />
                    <SPLIT distance="200" swimtime="00:02:08.32" />
                    <SPLIT distance="250" swimtime="00:02:41.89" />
                    <SPLIT distance="300" swimtime="00:03:15.95" />
                    <SPLIT distance="350" swimtime="00:03:50.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Weronika" lastname="Mrożek" birthdate="2004-02-22" gender="F" nation="POL" license="100116601298" swrid="4939220" athleteid="47087">
              <RESULTS>
                <RESULT eventid="44380" points="574" reactiontime="+69" swimtime="00:01:02.21" resultid="47088" heatid="50688" lane="3" entrytime="00:01:00.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46287" points="655" reactiontime="+65" swimtime="00:09:18.06" resultid="47089" heatid="50792" lane="4" entrytime="00:09:25.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                    <SPLIT distance="100" swimtime="00:01:07.05" />
                    <SPLIT distance="150" swimtime="00:01:42.00" />
                    <SPLIT distance="200" swimtime="00:02:16.84" />
                    <SPLIT distance="250" swimtime="00:02:51.74" />
                    <SPLIT distance="300" swimtime="00:03:26.52" />
                    <SPLIT distance="350" swimtime="00:04:01.67" />
                    <SPLIT distance="400" swimtime="00:04:36.30" />
                    <SPLIT distance="450" swimtime="00:05:11.50" />
                    <SPLIT distance="500" swimtime="00:05:46.25" />
                    <SPLIT distance="550" swimtime="00:06:21.55" />
                    <SPLIT distance="600" swimtime="00:06:56.71" />
                    <SPLIT distance="650" swimtime="00:07:32.92" />
                    <SPLIT distance="700" swimtime="00:08:08.54" />
                    <SPLIT distance="750" swimtime="00:08:44.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="651" reactiontime="+54" swimtime="00:04:32.75" resultid="47090" heatid="50805" lane="4" entrytime="00:04:31.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.44" />
                    <SPLIT distance="100" swimtime="00:01:05.32" />
                    <SPLIT distance="150" swimtime="00:01:39.77" />
                    <SPLIT distance="200" swimtime="00:02:14.13" />
                    <SPLIT distance="250" swimtime="00:02:48.80" />
                    <SPLIT distance="300" swimtime="00:03:23.56" />
                    <SPLIT distance="350" swimtime="00:03:58.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Lisik" birthdate="2003-06-15" gender="M" nation="POL" license="100116701300" swrid="4793262" athleteid="47091">
              <RESULTS>
                <RESULT eventid="44382" points="481" reactiontime="+77" swimtime="00:00:33.10" resultid="47092" heatid="50695" lane="0" entrytime="00:00:32.48" entrycourse="LCM" />
                <RESULT eventid="44407" points="486" reactiontime="+68" swimtime="00:01:12.34" resultid="47093" heatid="50750" lane="9" entrytime="00:01:13.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Damian" lastname="Wojnowski" birthdate="2003-05-05" gender="M" nation="POL" license="100116701301" swrid="4902929" athleteid="47094">
              <RESULTS>
                <RESULT eventid="44394" points="687" reactiontime="+74" swimtime="00:00:58.75" resultid="47095" heatid="50723" lane="4" entrytime="00:00:59.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="588" reactiontime="+71" swimtime="00:02:13.57" resultid="47096" heatid="50784" lane="5" entrytime="00:02:09.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.62" />
                    <SPLIT distance="100" swimtime="00:01:05.12" />
                    <SPLIT distance="150" swimtime="00:01:39.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46310" points="661" reactiontime="+67" swimtime="00:00:27.54" resultid="47097" heatid="50862" lane="5" entrytime="00:00:26.76" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Szmit" birthdate="2004-03-17" gender="M" nation="POL" license="100116701303" swrid="4847864" athleteid="47079">
              <RESULTS>
                <RESULT eventid="44378" points="658" reactiontime="+65" swimtime="00:00:53.92" resultid="47080" heatid="50677" lane="8" entrytime="00:00:53.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="658" reactiontime="+66" swimtime="00:00:25.60" resultid="47081" heatid="50769" lane="6" entrytime="00:00:25.59" entrycourse="LCM" />
                <RESULT eventid="46298" points="620" reactiontime="+64" swimtime="00:00:24.51" resultid="47082" heatid="50822" lane="1" entrytime="00:00:24.59" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04401" nation="POL" region="01" clubid="49893" name="Bielawski KS Swim Team Bielawa">
          <ATHLETES>
            <ATHLETE firstname="Jakub" lastname="Grabowy" birthdate="2002-09-26" gender="M" nation="POL" license="104401700036" swrid="5202272" athleteid="49894">
              <RESULTS>
                <RESULT eventid="44403" points="387" reactiontime="+78" swimtime="00:02:19.87" resultid="49895" heatid="50732" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.88" />
                    <SPLIT distance="100" swimtime="00:01:04.39" />
                    <SPLIT distance="150" swimtime="00:01:41.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="439" reactiontime="+71" swimtime="00:01:14.80" resultid="49896" heatid="50746" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="503" reactiontime="+68" swimtime="00:00:26.29" resultid="49897" heatid="50814" lane="5" entrytime="00:00:31.16" entrycourse="LCM" />
                <RESULT eventid="46302" points="363" reactiontime="+67" swimtime="00:02:56.74" resultid="49898" heatid="50836" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.93" />
                    <SPLIT distance="100" swimtime="00:01:25.90" />
                    <SPLIT distance="150" swimtime="00:02:12.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03415" nation="POL" region="15" clubid="48054" name="Uks Cityzen">
          <ATHLETES>
            <ATHLETE firstname="Alex" lastname="Baranowski" birthdate="2007-02-27" gender="M" nation="POL" license="103415700115" swrid="5405709" athleteid="48055">
              <RESULTS>
                <RESULT eventid="44378" points="436" reactiontime="+71" swimtime="00:01:01.84" resultid="48056" heatid="50671" lane="3" entrytime="00:01:02.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="439" reactiontime="+71" swimtime="00:02:14.20" resultid="48057" heatid="50732" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.39" />
                    <SPLIT distance="100" swimtime="00:01:04.76" />
                    <SPLIT distance="150" swimtime="00:01:39.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="319" reactiontime="+71" swimtime="00:00:32.59" resultid="48058" heatid="50764" lane="8" entrytime="00:00:32.65" entrycourse="LCM" />
                <RESULT eventid="46294" points="439" reactiontime="+74" swimtime="00:04:49.56" resultid="48059" heatid="50799" lane="3" entrytime="00:04:48.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                    <SPLIT distance="100" swimtime="00:01:07.34" />
                    <SPLIT distance="150" swimtime="00:01:44.29" />
                    <SPLIT distance="200" swimtime="00:02:22.07" />
                    <SPLIT distance="250" swimtime="00:02:59.44" />
                    <SPLIT distance="300" swimtime="00:03:37.70" />
                    <SPLIT distance="350" swimtime="00:04:14.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46306" points="261" reactiontime="+68" swimtime="00:01:17.37" resultid="48060" heatid="50844" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kamil" lastname="Kaczmarek" birthdate="2007-12-22" gender="M" nation="POL" license="103415700092" swrid="5198919" athleteid="48090">
              <RESULTS>
                <RESULT eventid="44394" points="482" reactiontime="+63" swimtime="00:01:06.09" resultid="48091" heatid="50723" lane="9" entrytime="00:01:06.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="474" reactiontime="+60" swimtime="00:02:10.79" resultid="48092" heatid="50733" lane="5" entrytime="00:02:36.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.84" />
                    <SPLIT distance="100" swimtime="00:01:03.05" />
                    <SPLIT distance="150" swimtime="00:01:37.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="460" reactiontime="+61" swimtime="00:02:24.89" resultid="48093" heatid="50784" lane="0" entrytime="00:02:26.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                    <SPLIT distance="100" swimtime="00:01:12.67" />
                    <SPLIT distance="150" swimtime="00:01:49.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="491" reactiontime="+65" swimtime="00:04:38.78" resultid="48094" heatid="50798" lane="6" entrytime="00:05:16.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.06" />
                    <SPLIT distance="100" swimtime="00:01:03.60" />
                    <SPLIT distance="150" swimtime="00:01:39.03" />
                    <SPLIT distance="200" swimtime="00:02:15.10" />
                    <SPLIT distance="250" swimtime="00:02:51.93" />
                    <SPLIT distance="300" swimtime="00:03:28.55" />
                    <SPLIT distance="350" swimtime="00:04:04.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46310" points="440" reactiontime="+60" swimtime="00:00:31.54" resultid="48095" heatid="50860" lane="1" entrytime="00:00:35.09" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Norbert" lastname="Gorzeń" birthdate="2006-06-03" gender="M" nation="POL" license="103415700019" swrid="5138790" athleteid="48073">
              <RESULTS>
                <RESULT eventid="44378" points="434" reactiontime="+74" swimtime="00:01:01.95" resultid="48074" heatid="50666" lane="2" entrytime="00:01:16.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44390" points="397" reactiontime="+73" swimtime="00:02:35.03" resultid="48075" heatid="50708" lane="5" entrytime="00:03:08.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                    <SPLIT distance="100" swimtime="00:01:13.71" />
                    <SPLIT distance="150" swimtime="00:02:00.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46285" points="386" reactiontime="+77" swimtime="00:19:56.09" resultid="48076" heatid="50789" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.89" />
                    <SPLIT distance="100" swimtime="00:01:14.00" />
                    <SPLIT distance="150" swimtime="00:01:53.46" />
                    <SPLIT distance="200" swimtime="00:02:33.43" />
                    <SPLIT distance="250" swimtime="00:03:12.93" />
                    <SPLIT distance="300" swimtime="00:03:53.22" />
                    <SPLIT distance="350" swimtime="00:04:33.48" />
                    <SPLIT distance="400" swimtime="00:05:14.17" />
                    <SPLIT distance="450" swimtime="00:05:54.75" />
                    <SPLIT distance="500" swimtime="00:06:35.93" />
                    <SPLIT distance="550" swimtime="00:07:15.67" />
                    <SPLIT distance="600" swimtime="00:07:56.20" />
                    <SPLIT distance="650" swimtime="00:08:36.52" />
                    <SPLIT distance="700" swimtime="00:09:17.03" />
                    <SPLIT distance="750" swimtime="00:09:56.92" />
                    <SPLIT distance="800" swimtime="00:10:37.23" />
                    <SPLIT distance="850" swimtime="00:11:16.74" />
                    <SPLIT distance="900" swimtime="00:11:57.02" />
                    <SPLIT distance="950" swimtime="00:12:36.88" />
                    <SPLIT distance="1000" swimtime="00:13:17.23" />
                    <SPLIT distance="1050" swimtime="00:13:56.76" />
                    <SPLIT distance="1100" swimtime="00:14:36.92" />
                    <SPLIT distance="1150" swimtime="00:15:16.88" />
                    <SPLIT distance="1200" swimtime="00:15:57.61" />
                    <SPLIT distance="1250" swimtime="00:16:37.97" />
                    <SPLIT distance="1300" swimtime="00:17:18.48" />
                    <SPLIT distance="1350" swimtime="00:17:58.79" />
                    <SPLIT distance="1400" swimtime="00:18:38.90" />
                    <SPLIT distance="1450" swimtime="00:19:18.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="387" reactiontime="+74" swimtime="00:05:01.98" resultid="48077" heatid="50799" lane="0" entrytime="00:04:58.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                    <SPLIT distance="100" swimtime="00:01:09.05" />
                    <SPLIT distance="150" swimtime="00:01:46.26" />
                    <SPLIT distance="200" swimtime="00:02:25.34" />
                    <SPLIT distance="250" swimtime="00:03:04.12" />
                    <SPLIT distance="300" swimtime="00:03:44.12" />
                    <SPLIT distance="350" swimtime="00:04:23.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kostiantyn" lastname="Surkov" birthdate="2006-07-05" gender="M" nation="POL" license="103415700088" swrid="5058525" athleteid="48067">
              <RESULTS>
                <RESULT eventid="44378" points="293" reactiontime="+80" swimtime="00:01:10.57" resultid="48068" heatid="50666" lane="0" entrytime="00:01:26.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44390" points="257" reactiontime="+72" swimtime="00:02:59.13" resultid="48069" heatid="50708" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                    <SPLIT distance="100" swimtime="00:01:27.33" />
                    <SPLIT distance="150" swimtime="00:02:17.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="271" reactiontime="+76" swimtime="00:01:27.82" resultid="48070" heatid="50746" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="239" reactiontime="+74" swimtime="00:00:35.86" resultid="48071" heatid="50761" lane="3" />
                <RESULT eventid="46298" points="285" reactiontime="+66" swimtime="00:00:31.77" resultid="48072" heatid="50812" lane="7" entrytime="00:00:36.48" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Troszczyński" birthdate="2007-12-16" gender="M" nation="POL" license="103415700094" swrid="5198889" athleteid="48084">
              <RESULTS>
                <RESULT eventid="44386" points="368" reactiontime="+69" swimtime="00:02:34.46" resultid="48085" heatid="50705" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                    <SPLIT distance="100" swimtime="00:01:10.40" />
                    <SPLIT distance="150" swimtime="00:01:52.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="354" reactiontime="+75" swimtime="00:01:13.26" resultid="48086" heatid="50718" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="376" reactiontime="+69" swimtime="00:00:30.85" resultid="48087" heatid="50761" lane="6" />
                <RESULT eventid="46306" points="360" reactiontime="+66" swimtime="00:01:09.53" resultid="48088" heatid="50848" lane="9" entrytime="00:01:08.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46310" points="342" reactiontime="+67" swimtime="00:00:34.31" resultid="48089" heatid="50861" lane="0" entrytime="00:00:32.36" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Gulczyńska" birthdate="2007-08-25" gender="F" nation="POL" license="103415600093" swrid="5198895" athleteid="48078">
              <RESULTS>
                <RESULT eventid="44380" points="497" reactiontime="+65" swimtime="00:01:05.27" resultid="48079" heatid="50686" lane="0" entrytime="00:01:04.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44384" points="491" reactiontime="+63" swimtime="00:00:37.25" resultid="48080" heatid="50701" lane="5" entrytime="00:00:38.13" entrycourse="LCM" />
                <RESULT eventid="44409" points="444" reactiontime="+61" swimtime="00:01:24.01" resultid="48081" heatid="50751" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="407" reactiontime="+63" swimtime="00:00:32.95" resultid="48082" heatid="50777" lane="6" entrytime="00:00:32.86" entrycourse="LCM" />
                <RESULT eventid="46300" points="475" reactiontime="+60" swimtime="00:00:30.33" resultid="48083" heatid="50832" lane="8" entrytime="00:00:29.95" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kamil" lastname="Bosiacki" birthdate="2007-01-22" gender="M" nation="POL" license="103415700068" swrid="5278372" athleteid="48061">
              <RESULTS>
                <RESULT eventid="44378" points="298" reactiontime="+62" swimtime="00:01:10.21" resultid="48062" heatid="50666" lane="9" entrytime="00:01:29.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="332" reactiontime="+56" swimtime="00:00:37.47" resultid="48063" heatid="50694" lane="9" entrytime="00:00:36.18" entrycourse="LCM" />
                <RESULT eventid="44407" points="288" swimtime="00:01:26.11" resultid="48064" heatid="50748" lane="4" entrytime="00:01:23.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="267" reactiontime="+73" swimtime="00:00:32.47" resultid="48065" heatid="50812" lane="8" entrytime="00:00:37.85" entrycourse="LCM" />
                <RESULT eventid="46302" points="324" reactiontime="+74" swimtime="00:03:03.51" resultid="48066" heatid="50838" lane="2" entrytime="00:03:30.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.39" />
                    <SPLIT distance="100" swimtime="00:01:27.64" />
                    <SPLIT distance="150" swimtime="00:02:16.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="44399" points="390" reactiontime="+61" swimtime="00:04:43.70" resultid="48096" heatid="50730" lane="7" entrytime="00:04:37.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                    <SPLIT distance="100" swimtime="00:01:08.08" />
                    <SPLIT distance="150" swimtime="00:01:46.52" />
                    <SPLIT distance="200" swimtime="00:02:32.56" />
                    <SPLIT distance="250" swimtime="00:03:04.61" />
                    <SPLIT distance="300" swimtime="00:03:41.85" />
                    <SPLIT distance="350" swimtime="00:04:10.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="48090" number="1" reactiontime="+61" />
                    <RELAYPOSITION athleteid="48061" number="2" reactiontime="+28" />
                    <RELAYPOSITION athleteid="48084" number="3" reactiontime="+44" />
                    <RELAYPOSITION athleteid="48055" number="4" reactiontime="+52" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46289" points="398" reactiontime="+54" swimtime="00:04:15.71" resultid="48097" heatid="50794" lane="0" entrytime="00:04:10.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.37" />
                    <SPLIT distance="100" swimtime="00:00:59.85" />
                    <SPLIT distance="150" swimtime="00:01:29.00" />
                    <SPLIT distance="200" swimtime="00:02:02.20" />
                    <SPLIT distance="250" swimtime="00:02:36.07" />
                    <SPLIT distance="300" swimtime="00:03:12.78" />
                    <SPLIT distance="350" swimtime="00:03:42.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="48090" number="1" reactiontime="+54" />
                    <RELAYPOSITION athleteid="48084" number="2" reactiontime="+27" />
                    <RELAYPOSITION athleteid="48061" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="48055" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00114" nation="POL" region="14" clubid="46464" name="AZS AWF Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Marcelina" lastname="Dopart" birthdate="2003-04-14" gender="F" nation="POL" license="100114600105" swrid="4012857" athleteid="46465">
              <RESULTS>
                <RESULT eventid="44384" points="572" reactiontime="+72" swimtime="00:00:35.41" resultid="46466" heatid="50703" lane="6" entrytime="00:00:34.33" entrycourse="LCM" />
                <RESULT eventid="44392" points="545" reactiontime="+73" swimtime="00:02:34.36" resultid="46467" heatid="50716" lane="9" entrytime="00:02:34.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                    <SPLIT distance="100" swimtime="00:01:14.45" />
                    <SPLIT distance="150" swimtime="00:01:58.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44409" points="491" reactiontime="+72" swimtime="00:01:21.25" resultid="46468" heatid="50756" lane="2" entrytime="00:01:16.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="562" reactiontime="+71" swimtime="00:00:28.67" resultid="46469" heatid="50834" lane="4" entrytime="00:00:28.05" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Obajtek" birthdate="2003-01-19" gender="F" nation="POL" license="100114600108" swrid="4695906" athleteid="46470">
              <RESULTS>
                <RESULT eventid="44384" points="612" reactiontime="+63" swimtime="00:00:34.61" resultid="46471" heatid="50703" lane="3" entrytime="00:00:34.25" entrycourse="LCM" />
                <RESULT eventid="44392" points="622" reactiontime="+66" swimtime="00:02:27.71" resultid="46472" heatid="50716" lane="3" entrytime="00:02:27.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                    <SPLIT distance="100" swimtime="00:01:12.41" />
                    <SPLIT distance="150" swimtime="00:01:53.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44409" points="620" reactiontime="+64" swimtime="00:01:15.19" resultid="46473" heatid="50756" lane="5" entrytime="00:01:15.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46304" points="618" reactiontime="+57" swimtime="00:02:43.28" resultid="46474" heatid="50843" lane="4" entrytime="00:02:41.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.38" />
                    <SPLIT distance="100" swimtime="00:01:18.96" />
                    <SPLIT distance="150" swimtime="00:02:00.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00501" nation="POL" region="01" clubid="48160" name="UKS Energetyk Zgorzelec">
          <ATHLETES>
            <ATHLETE firstname="Natalia" lastname="Skoczylas" birthdate="2008-10-07" gender="F" nation="POL" license="100501600035" swrid="5334425" athleteid="48191">
              <RESULTS>
                <RESULT eventid="44380" points="353" reactiontime="+57" swimtime="00:01:13.12" resultid="48192" heatid="50679" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="331" swimtime="00:00:35.31" resultid="48193" heatid="50772" lane="5" />
                <RESULT eventid="46300" points="395" reactiontime="+56" swimtime="00:00:32.26" resultid="48194" heatid="50823" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Borowiecki" birthdate="2004-09-07" gender="M" nation="POL" license="100501700034" athleteid="48173">
              <RESULTS>
                <RESULT eventid="44378" points="582" reactiontime="+64" swimtime="00:00:56.16" resultid="48174" heatid="50663" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="510" reactiontime="+66" swimtime="00:00:32.47" resultid="48175" heatid="50690" lane="4" />
                <RESULT eventid="44411" points="599" reactiontime="+66" swimtime="00:00:26.41" resultid="48176" heatid="50760" lane="7" />
                <RESULT eventid="46298" points="592" reactiontime="+68" swimtime="00:00:24.89" resultid="48177" heatid="50806" lane="3" />
                <RESULT eventid="46310" points="512" reactiontime="+60" swimtime="00:00:29.99" resultid="48178" heatid="50857" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sebastian" lastname="Bałdyga" birthdate="2006-06-05" gender="M" nation="POL" license="100501700022" swrid="5024299" athleteid="48161">
              <RESULTS>
                <RESULT eventid="44378" points="481" reactiontime="+79" swimtime="00:00:59.84" resultid="48162" heatid="50663" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="431" reactiontime="+54" swimtime="00:01:08.59" resultid="48163" heatid="50719" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="403" reactiontime="+59" swimtime="00:02:31.45" resultid="48164" heatid="50781" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                    <SPLIT distance="100" swimtime="00:01:12.70" />
                    <SPLIT distance="150" swimtime="00:01:52.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="474" reactiontime="+74" swimtime="00:00:26.80" resultid="48165" heatid="50807" lane="8" />
                <RESULT eventid="46310" points="419" reactiontime="+54" swimtime="00:00:32.07" resultid="48166" heatid="50858" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Leśniewska" birthdate="2006-06-01" gender="F" nation="POL" license="100501600026" swrid="5072876" athleteid="48179">
              <RESULTS>
                <RESULT eventid="44380" points="372" reactiontime="+79" swimtime="00:01:11.88" resultid="48180" heatid="50679" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="349" reactiontime="+77" swimtime="00:00:34.68" resultid="48181" heatid="50772" lane="3" />
                <RESULT eventid="46300" points="408" reactiontime="+78" swimtime="00:00:31.89" resultid="48182" heatid="50825" lane="1" />
                <RESULT eventid="46308" points="278" reactiontime="+79" swimtime="00:01:24.92" resultid="48183" heatid="50897" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Daszyński" birthdate="1948-11-29" gender="M" nation="POL" athleteid="50884">
              <RESULTS>
                <RESULT eventid="44394" points="84" reactiontime="+89" swimtime="00:01:58.39" resultid="50885" heatid="50717" lane="6" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44386" points="33" swimtime="00:05:41.91" resultid="50886" heatid="50704" lane="6" late="yes">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:04:14.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="69" reactiontime="+87" swimtime="00:02:18.48" resultid="50889" heatid="50745" lane="6" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="87" reactiontime="+90" swimtime="00:04:11.88" resultid="50890" heatid="50780" lane="6" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.76" />
                    <SPLIT distance="100" swimtime="00:02:05.80" />
                    <SPLIT distance="150" swimtime="00:03:10.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" status="DNS" swimtime="00:00:00.00" resultid="50891" heatid="50796" lane="2" late="yes" />
                <RESULT eventid="46306" points="36" reactiontime="+98" swimtime="00:02:29.24" resultid="50892" heatid="50844" lane="8" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="107" reactiontime="+92" swimtime="00:00:43.92" resultid="50910" heatid="50806" lane="7" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Kurasiewicz" birthdate="2007-03-15" gender="F" nation="POL" license="100501600033" swrid="4901148" athleteid="48184">
              <RESULTS>
                <RESULT eventid="44380" points="362" reactiontime="+91" swimtime="00:01:12.51" resultid="48185" heatid="50678" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44392" points="288" reactiontime="+76" swimtime="00:03:10.91" resultid="48186" heatid="50712" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.65" />
                    <SPLIT distance="100" swimtime="00:01:29.75" />
                    <SPLIT distance="150" swimtime="00:02:27.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44396" points="275" reactiontime="+66" swimtime="00:01:28.45" resultid="48187" heatid="50724" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="278" reactiontime="+82" swimtime="00:00:37.40" resultid="48188" heatid="50770" lane="1" />
                <RESULT eventid="46300" points="383" reactiontime="+74" swimtime="00:00:32.57" resultid="48189" heatid="50825" lane="5" />
                <RESULT eventid="46312" points="284" reactiontime="+63" swimtime="00:00:41.03" resultid="48190" heatid="50903" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominik" lastname="Leśniewski" birthdate="2004-08-02" gender="M" nation="POL" license="100501700025" swrid="4931181" athleteid="48167">
              <RESULTS>
                <RESULT eventid="44378" points="483" reactiontime="+71" swimtime="00:00:59.76" resultid="48168" heatid="50671" lane="1" entrytime="00:01:03.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="378" reactiontime="+68" swimtime="00:01:11.69" resultid="48169" heatid="50718" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="516" reactiontime="+70" swimtime="00:00:27.76" resultid="48170" heatid="50765" lane="8" entrytime="00:00:30.93" entrycourse="LCM" />
                <RESULT eventid="46298" points="465" reactiontime="+70" swimtime="00:00:26.99" resultid="48171" heatid="50816" lane="4" entrytime="00:00:28.53" entrycourse="LCM" />
                <RESULT eventid="46306" points="366" reactiontime="+69" swimtime="00:01:09.20" resultid="48172" heatid="50845" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Koprowicz" birthdate="2005-01-26" gender="F" nation="POL" license="100501600046" swrid="5458593" athleteid="48195">
              <RESULTS>
                <RESULT eventid="44384" points="350" reactiontime="+53" swimtime="00:00:41.70" resultid="48196" heatid="50698" lane="9" />
                <RESULT eventid="46300" points="433" reactiontime="+62" swimtime="00:00:31.27" resultid="48197" heatid="50827" lane="0" />
                <RESULT eventid="46312" points="378" reactiontime="+56" swimtime="00:00:37.29" resultid="48198" heatid="50905" lane="1" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01015" nation="POL" region="15" clubid="48585" name="UKS Trójka Środa Wlkp.">
          <ATHLETES>
            <ATHLETE firstname="Krystyna" lastname="Kwiecińska" birthdate="2004-12-12" gender="F" nation="POL" license="101015600048" swrid="5163617" athleteid="48600">
              <RESULTS>
                <RESULT eventid="44384" points="476" reactiontime="+53" swimtime="00:00:37.63" resultid="48601" heatid="50701" lane="4" entrytime="00:00:37.98" entrycourse="LCM" />
                <RESULT eventid="44409" points="483" reactiontime="+77" swimtime="00:01:21.73" resultid="48602" heatid="50755" lane="2" entrytime="00:01:21.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46304" points="504" reactiontime="+76" swimtime="00:02:54.76" resultid="48603" heatid="50843" lane="0" entrytime="00:02:56.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.28" />
                    <SPLIT distance="100" swimtime="00:01:23.60" />
                    <SPLIT distance="150" swimtime="00:02:09.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcelina" lastname="Mieloch" birthdate="2005-07-24" gender="F" nation="POL" license="101015600044" swrid="5117134" athleteid="48604">
              <RESULTS>
                <RESULT eventid="44396" points="418" reactiontime="+61" swimtime="00:01:16.95" resultid="48605" heatid="50726" lane="5" entrytime="00:01:17.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44417" points="378" reactiontime="+70" swimtime="00:02:50.46" resultid="48606" heatid="50788" lane="9" entrytime="00:02:48.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.26" />
                    <SPLIT distance="100" swimtime="00:01:21.94" />
                    <SPLIT distance="150" swimtime="00:02:07.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="452" reactiontime="+63" swimtime="00:00:35.14" resultid="48607" heatid="50907" lane="6" entrytime="00:00:35.87" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kamil" lastname="Nowak" birthdate="2005-08-04" gender="M" nation="POL" license="101015700036" swrid="5117131" athleteid="48586">
              <RESULTS>
                <RESULT eventid="44378" points="488" reactiontime="+69" swimtime="00:00:59.58" resultid="48587" heatid="50673" lane="9" entrytime="00:01:01.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="429" reactiontime="+76" swimtime="00:00:29.51" resultid="48588" heatid="50765" lane="7" entrytime="00:00:30.74" entrycourse="LCM" />
                <RESULT eventid="46298" points="452" reactiontime="+79" swimtime="00:00:27.23" resultid="48589" heatid="50817" lane="7" entrytime="00:00:28.16" entrycourse="LCM" />
                <RESULT eventid="46306" points="395" reactiontime="+69" swimtime="00:01:07.41" resultid="48590" heatid="50847" lane="4" entrytime="00:01:08.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Perlik" birthdate="2006-09-24" gender="F" nation="POL" license="101015600057" swrid="5153534" athleteid="48591">
              <RESULTS>
                <RESULT eventid="44380" points="479" reactiontime="+79" swimtime="00:01:06.07" resultid="48592" heatid="50683" lane="7" entrytime="00:01:09.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="377" swimtime="00:00:33.80" resultid="48593" heatid="50776" lane="4" entrytime="00:00:33.64" entrycourse="LCM" />
                <RESULT eventid="46300" points="488" reactiontime="+79" swimtime="00:00:30.05" resultid="48594" heatid="50831" lane="0" entrytime="00:00:31.02" entrycourse="LCM" />
                <RESULT eventid="46308" points="362" reactiontime="+74" swimtime="00:01:17.81" resultid="48595" heatid="50899" lane="7" entrytime="00:01:19.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Kucharska" birthdate="2005-01-04" gender="F" nation="POL" license="101015600037" swrid="5096958" athleteid="48596">
              <RESULTS>
                <RESULT eventid="44384" points="606" reactiontime="+68" swimtime="00:00:34.73" resultid="48597" heatid="50703" lane="0" entrytime="00:00:34.93" entrycourse="LCM" />
                <RESULT eventid="44409" points="515" reactiontime="+69" swimtime="00:01:19.98" resultid="48598" heatid="50756" lane="1" entrytime="00:01:17.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46304" points="447" reactiontime="+65" swimtime="00:03:01.89" resultid="48599" heatid="50843" lane="8" entrytime="00:02:53.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                    <SPLIT distance="100" swimtime="00:01:27.37" />
                    <SPLIT distance="150" swimtime="00:02:15.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00101" nation="POL" region="01" clubid="50312" name="MKS Juvenia Wrocław">
          <ATHLETES>
            <ATHLETE firstname="Igor" lastname="Wierzbicki" birthdate="2005-06-25" gender="M" nation="POL" license="100101701334" swrid="5147678" athleteid="50560">
              <RESULTS>
                <RESULT eventid="44390" points="523" reactiontime="+68" swimtime="00:02:21.49" resultid="50561" heatid="50711" lane="3" entrytime="00:02:20.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.35" />
                    <SPLIT distance="100" swimtime="00:01:05.69" />
                    <SPLIT distance="150" swimtime="00:01:49.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="564" reactiontime="+63" swimtime="00:02:03.43" resultid="50562" heatid="50738" lane="4" entrytime="00:02:04.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.68" />
                    <SPLIT distance="100" swimtime="00:00:58.96" />
                    <SPLIT distance="150" swimtime="00:01:32.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="497" reactiontime="+65" swimtime="00:00:28.11" resultid="50563" heatid="50768" lane="9" entrytime="00:00:27.88" entrycourse="LCM" />
                <RESULT eventid="46298" points="501" reactiontime="+66" swimtime="00:00:26.32" resultid="50564" heatid="50819" lane="1" entrytime="00:00:26.56" entrycourse="LCM" />
                <RESULT eventid="46310" points="474" reactiontime="+64" swimtime="00:00:30.76" resultid="50565" heatid="50861" lane="3" entrytime="00:00:30.87" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hanna" lastname="Gryncewicz" birthdate="2008-05-22" gender="F" nation="POL" license="100101601340" swrid="5165967" athleteid="50532">
              <RESULTS>
                <RESULT eventid="44384" points="278" reactiontime="+77" swimtime="00:00:45.04" resultid="50533" heatid="50699" lane="4" entrytime="00:00:47.74" entrycourse="LCM" />
                <RESULT eventid="44396" points="284" reactiontime="+87" swimtime="00:01:27.58" resultid="50534" heatid="50725" lane="8" entrytime="00:01:27.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44409" points="247" reactiontime="+90" swimtime="00:01:42.15" resultid="50535" heatid="50753" lane="9" entrytime="00:01:43.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="365" reactiontime="+89" swimtime="00:00:33.12" resultid="50536" heatid="50823" lane="3" />
                <RESULT eventid="46312" points="279" reactiontime="+86" swimtime="00:00:41.26" resultid="50537" heatid="50906" lane="5" entrytime="00:00:39.05" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Malik" birthdate="2007-02-01" gender="M" nation="POL" license="100101701290" swrid="5244057" athleteid="50369">
              <RESULTS>
                <RESULT eventid="44378" points="366" reactiontime="+71" swimtime="00:01:05.55" resultid="50370" heatid="50669" lane="0" entrytime="00:01:06.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="331" reactiontime="+78" swimtime="00:00:37.49" resultid="50371" heatid="50692" lane="1" />
                <RESULT eventid="44407" points="332" reactiontime="+77" swimtime="00:01:22.12" resultid="50372" heatid="50748" lane="6" entrytime="00:01:25.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="346" reactiontime="+58" swimtime="00:02:39.42" resultid="50373" heatid="50781" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.07" />
                    <SPLIT distance="100" swimtime="00:01:19.59" />
                    <SPLIT distance="150" swimtime="00:02:00.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="344" reactiontime="+73" swimtime="00:00:29.84" resultid="50374" heatid="50808" lane="2" />
                <RESULT eventid="46310" points="349" reactiontime="+59" swimtime="00:00:34.07" resultid="50375" heatid="50858" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Kołtuniewicz" birthdate="2007-09-02" gender="F" nation="POL" license="100101601189" swrid="5088589" athleteid="50508">
              <RESULTS>
                <RESULT eventid="44384" points="418" reactiontime="+71" swimtime="00:00:39.29" resultid="50509" heatid="50697" lane="0" />
                <RESULT eventid="44392" points="422" reactiontime="+76" swimtime="00:02:48.02" resultid="50510" heatid="50714" lane="1" entrytime="00:02:52.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.96" />
                    <SPLIT distance="100" swimtime="00:01:20.76" />
                    <SPLIT distance="150" swimtime="00:02:07.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44409" points="416" reactiontime="+78" swimtime="00:01:25.87" resultid="50511" heatid="50754" lane="1" entrytime="00:01:28.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="373" reactiontime="+65" swimtime="00:00:33.91" resultid="50512" heatid="50772" lane="4" />
                <RESULT eventid="46304" points="462" reactiontime="+75" swimtime="00:02:59.92" resultid="50513" heatid="50841" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.49" />
                    <SPLIT distance="100" swimtime="00:01:26.89" />
                    <SPLIT distance="150" swimtime="00:02:13.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46308" points="331" reactiontime="+74" swimtime="00:01:20.17" resultid="50514" heatid="50899" lane="1" entrytime="00:01:20.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Olszowiec" birthdate="2007-01-04" gender="M" nation="POL" license="100101701258" swrid="5001973" athleteid="50313">
              <RESULTS>
                <RESULT eventid="44378" points="482" reactiontime="+74" swimtime="00:00:59.79" resultid="50314" heatid="50673" lane="5" entrytime="00:00:59.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="327" reactiontime="+76" swimtime="00:00:37.66" resultid="50315" heatid="50689" lane="7" />
                <RESULT eventid="44403" points="423" reactiontime="+74" swimtime="00:02:15.84" resultid="50316" heatid="50736" lane="8" entrytime="00:02:19.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                    <SPLIT distance="100" swimtime="00:01:05.61" />
                    <SPLIT distance="150" swimtime="00:01:41.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="411" reactiontime="+77" swimtime="00:00:29.93" resultid="50317" heatid="50764" lane="3" entrytime="00:00:32.06" entrycourse="LCM" />
                <RESULT eventid="46298" points="455" reactiontime="+76" swimtime="00:00:27.17" resultid="50318" heatid="50809" lane="6" />
                <RESULT eventid="46310" points="378" reactiontime="+75" swimtime="00:00:33.18" resultid="50319" heatid="50856" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mikołaj" lastname="Koczerga" birthdate="2007-08-28" gender="M" nation="POL" license="100101701366" swrid="5416712" athleteid="50335">
              <RESULTS>
                <RESULT eventid="44378" points="333" reactiontime="+66" swimtime="00:01:07.66" resultid="50336" heatid="50667" lane="5" entrytime="00:01:07.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44390" points="336" reactiontime="+62" swimtime="00:02:43.90" resultid="50337" heatid="50709" lane="4" entrytime="00:02:43.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.81" />
                    <SPLIT distance="100" swimtime="00:01:19.97" />
                    <SPLIT distance="150" swimtime="00:02:07.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="320" reactiontime="+66" swimtime="00:02:29.05" resultid="50338" heatid="50735" lane="9" entrytime="00:02:28.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.30" />
                    <SPLIT distance="100" swimtime="00:01:13.31" />
                    <SPLIT distance="150" swimtime="00:01:53.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="271" reactiontime="+63" swimtime="00:00:34.40" resultid="50339" heatid="50758" lane="0" />
                <RESULT eventid="46294" points="360" reactiontime="+66" swimtime="00:05:09.21" resultid="50340" heatid="50798" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.49" />
                    <SPLIT distance="100" swimtime="00:01:13.14" />
                    <SPLIT distance="150" swimtime="00:01:52.83" />
                    <SPLIT distance="200" swimtime="00:02:32.64" />
                    <SPLIT distance="250" swimtime="00:03:12.89" />
                    <SPLIT distance="300" swimtime="00:03:52.53" />
                    <SPLIT distance="350" swimtime="00:04:32.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46306" points="279" reactiontime="+64" swimtime="00:01:15.70" resultid="50341" heatid="50846" lane="5" entrytime="00:01:16.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mikołaj" lastname="Rosiński" birthdate="2007-12-06" gender="M" nation="POL" license="100101701295" swrid="5244108" athleteid="50376">
              <RESULTS>
                <RESULT eventid="44378" points="362" reactiontime="+80" swimtime="00:01:05.78" resultid="50377" heatid="50668" lane="7" entrytime="00:01:06.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="329" reactiontime="+91" swimtime="00:01:15.05" resultid="50378" heatid="50721" lane="6" entrytime="00:01:15.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="279" reactiontime="+78" swimtime="00:00:34.06" resultid="50379" heatid="50760" lane="6" />
                <RESULT eventid="44415" points="323" reactiontime="+91" swimtime="00:02:43.01" resultid="50380" heatid="50781" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.80" />
                    <SPLIT distance="100" swimtime="00:01:19.36" />
                    <SPLIT distance="150" swimtime="00:02:01.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="336" reactiontime="+82" swimtime="00:00:30.05" resultid="50381" heatid="50807" lane="1" />
                <RESULT eventid="46306" points="284" reactiontime="+80" swimtime="00:01:15.23" resultid="50382" heatid="50846" lane="6" entrytime="00:01:17.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Mazurkiewicz" birthdate="2006-03-21" gender="F" nation="POL" license="100101601195" swrid="5088591" athleteid="50416">
              <RESULTS>
                <RESULT eventid="44380" points="428" reactiontime="+74" swimtime="00:01:08.57" resultid="50417" heatid="50683" lane="4" entrytime="00:01:08.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44392" points="456" reactiontime="+73" swimtime="00:02:43.79" resultid="50418" heatid="50715" lane="1" entrytime="00:02:42.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.83" />
                    <SPLIT distance="100" swimtime="00:01:17.92" />
                    <SPLIT distance="150" swimtime="00:02:06.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="423" reactiontime="+76" swimtime="00:02:30.47" resultid="50419" heatid="50742" lane="8" entrytime="00:02:28.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                    <SPLIT distance="100" swimtime="00:01:12.21" />
                    <SPLIT distance="150" swimtime="00:01:51.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46287" points="372" reactiontime="+76" swimtime="00:11:14.07" resultid="50420" heatid="50791" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                    <SPLIT distance="100" swimtime="00:01:14.95" />
                    <SPLIT distance="150" swimtime="00:01:56.45" />
                    <SPLIT distance="200" swimtime="00:02:39.09" />
                    <SPLIT distance="250" swimtime="00:03:21.45" />
                    <SPLIT distance="300" swimtime="00:04:04.69" />
                    <SPLIT distance="350" swimtime="00:04:47.85" />
                    <SPLIT distance="400" swimtime="00:05:31.00" />
                    <SPLIT distance="450" swimtime="00:06:14.07" />
                    <SPLIT distance="500" swimtime="00:06:57.28" />
                    <SPLIT distance="550" swimtime="00:07:40.74" />
                    <SPLIT distance="600" swimtime="00:08:24.75" />
                    <SPLIT distance="650" swimtime="00:09:07.91" />
                    <SPLIT distance="700" swimtime="00:09:51.18" />
                    <SPLIT distance="750" swimtime="00:10:33.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="400" reactiontime="+77" swimtime="00:05:20.70" resultid="50421" heatid="50803" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                    <SPLIT distance="100" swimtime="00:01:14.20" />
                    <SPLIT distance="150" swimtime="00:01:55.22" />
                    <SPLIT distance="200" swimtime="00:02:36.79" />
                    <SPLIT distance="250" swimtime="00:03:18.08" />
                    <SPLIT distance="300" swimtime="00:04:00.07" />
                    <SPLIT distance="350" swimtime="00:04:41.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46308" points="318" reactiontime="+77" swimtime="00:01:21.26" resultid="50422" heatid="50899" lane="6" entrytime="00:01:18.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Szymczak" birthdate="2003-05-27" gender="M" nation="POL" license="100101701175" swrid="4995388" athleteid="50404">
              <RESULTS>
                <RESULT eventid="44378" points="600" reactiontime="+65" swimtime="00:00:55.59" resultid="50405" heatid="50676" lane="8" entrytime="00:00:55.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="582" reactiontime="+66" swimtime="00:02:02.15" resultid="50406" heatid="50739" lane="1" entrytime="00:02:01.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.38" />
                    <SPLIT distance="100" swimtime="00:00:59.45" />
                    <SPLIT distance="150" swimtime="00:01:31.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="627" reactiontime="+69" swimtime="00:04:17.12" resultid="50407" heatid="50800" lane="5" entrytime="00:04:16.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.21" />
                    <SPLIT distance="100" swimtime="00:01:01.42" />
                    <SPLIT distance="150" swimtime="00:01:34.37" />
                    <SPLIT distance="200" swimtime="00:02:07.61" />
                    <SPLIT distance="250" swimtime="00:02:40.67" />
                    <SPLIT distance="300" swimtime="00:03:14.04" />
                    <SPLIT distance="350" swimtime="00:03:46.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46306" points="561" reactiontime="+67" swimtime="00:01:00.01" resultid="50408" heatid="50849" lane="2" entrytime="00:00:59.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daria" lastname="Shevhenko" birthdate="2006-06-24" gender="F" nation="POL" license="100101601370" swrid="4979441" athleteid="50409">
              <RESULTS>
                <RESULT eventid="44380" points="504" reactiontime="+75" swimtime="00:01:04.95" resultid="50410" heatid="50686" lane="2" entrytime="00:01:04.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44388" points="357" reactiontime="+69" swimtime="00:02:51.58" resultid="50411" heatid="50706" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                    <SPLIT distance="100" swimtime="00:01:18.70" />
                    <SPLIT distance="150" swimtime="00:02:04.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="430" reactiontime="+72" swimtime="00:02:29.68" resultid="50412" heatid="50742" lane="3" entrytime="00:02:23.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                    <SPLIT distance="100" swimtime="00:01:11.87" />
                    <SPLIT distance="150" swimtime="00:01:51.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="446" reactiontime="+71" swimtime="00:00:31.97" resultid="50413" heatid="50771" lane="8" />
                <RESULT eventid="46300" points="510" reactiontime="+77" swimtime="00:00:29.61" resultid="50414" heatid="50826" lane="6" />
                <RESULT eventid="46308" points="453" reactiontime="+73" swimtime="00:01:12.22" resultid="50415" heatid="50900" lane="2" entrytime="00:01:12.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nadia" lastname="Kertyńska" birthdate="2003-12-18" gender="F" nation="POL" license="100101601331" swrid="5023597" athleteid="50588">
              <RESULTS>
                <RESULT eventid="44392" points="647" reactiontime="+64" swimtime="00:02:25.77" resultid="50589" heatid="50716" lane="4" entrytime="00:02:25.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.22" />
                    <SPLIT distance="100" swimtime="00:01:10.36" />
                    <SPLIT distance="150" swimtime="00:01:52.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="669" reactiontime="+66" swimtime="00:02:09.14" resultid="50590" heatid="50744" lane="5" entrytime="00:02:10.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.73" />
                    <SPLIT distance="100" swimtime="00:01:02.92" />
                    <SPLIT distance="150" swimtime="00:01:36.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="528" reactiontime="+71" swimtime="00:00:30.21" resultid="50591" heatid="50771" lane="5" />
                <RESULT eventid="46300" points="697" reactiontime="+64" swimtime="00:00:26.69" resultid="50592" heatid="50835" lane="3" entrytime="00:00:26.97" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwia" lastname="Zagdańska" birthdate="2005-07-08" gender="F" nation="POL" license="100101601397" swrid="5024239" athleteid="50484">
              <RESULTS>
                <RESULT eventid="44380" points="615" reactiontime="+74" swimtime="00:01:00.80" resultid="50485" heatid="50688" lane="2" entrytime="00:01:00.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44392" points="608" reactiontime="+71" swimtime="00:02:28.86" resultid="50486" heatid="50716" lane="6" entrytime="00:02:29.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                    <SPLIT distance="100" swimtime="00:01:10.87" />
                    <SPLIT distance="150" swimtime="00:01:54.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="621" reactiontime="+73" swimtime="00:02:12.42" resultid="50487" heatid="50744" lane="7" entrytime="00:02:12.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.07" />
                    <SPLIT distance="100" swimtime="00:01:05.17" />
                    <SPLIT distance="150" swimtime="00:01:39.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="617" reactiontime="+72" swimtime="00:04:37.71" resultid="50488" heatid="50805" lane="5" entrytime="00:04:39.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="100" swimtime="00:01:05.71" />
                    <SPLIT distance="150" swimtime="00:01:40.80" />
                    <SPLIT distance="200" swimtime="00:02:16.15" />
                    <SPLIT distance="250" swimtime="00:02:52.00" />
                    <SPLIT distance="300" swimtime="00:03:27.85" />
                    <SPLIT distance="350" swimtime="00:04:03.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="584" reactiontime="+71" swimtime="00:00:28.31" resultid="50489" heatid="50834" lane="3" entrytime="00:00:28.14" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Polina" lastname="Żurawel" birthdate="2008-09-06" gender="F" nation="POL" license="100101601286" swrid="5266496" athleteid="50459">
              <RESULTS>
                <RESULT eventid="44380" points="448" reactiontime="+66" swimtime="00:01:07.53" resultid="50460" heatid="50684" lane="4" entrytime="00:01:06.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44396" points="425" reactiontime="+69" swimtime="00:01:16.52" resultid="50461" heatid="50727" lane="5" entrytime="00:01:13.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="409" reactiontime="+74" swimtime="00:00:32.91" resultid="50462" heatid="50776" lane="3" entrytime="00:00:33.88" entrycourse="LCM" />
                <RESULT eventid="44417" points="424" reactiontime="+74" swimtime="00:02:44.18" resultid="50463" heatid="50786" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.51" />
                    <SPLIT distance="100" swimtime="00:01:21.54" />
                    <SPLIT distance="150" swimtime="00:02:04.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="521" reactiontime="+72" swimtime="00:00:29.41" resultid="50464" heatid="50831" lane="2" entrytime="00:00:30.67" entrycourse="LCM" />
                <RESULT eventid="46312" points="508" reactiontime="+64" swimtime="00:00:33.81" resultid="50465" heatid="50908" lane="9" entrytime="00:00:35.43" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcel" lastname="Jaworski" birthdate="2004-01-17" gender="M" nation="POL" license="100101701332" swrid="5088670" athleteid="50593">
              <RESULTS>
                <RESULT eventid="44411" points="598" reactiontime="+64" swimtime="00:00:26.42" resultid="50594" heatid="50768" lane="4" entrytime="00:00:26.69" entrycourse="LCM" />
                <RESULT eventid="46298" points="559" reactiontime="+63" swimtime="00:00:25.37" resultid="50595" heatid="50821" lane="3" entrytime="00:00:25.18" entrycourse="LCM" />
                <RESULT eventid="46306" points="586" reactiontime="+66" swimtime="00:00:59.13" resultid="50596" heatid="50849" lane="1" entrytime="00:01:00.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Malwina" lastname="Malaczewska" birthdate="2005-07-05" gender="F" nation="POL" license="100101601337" swrid="5088658" athleteid="50521">
              <RESULTS>
                <RESULT eventid="44384" points="635" reactiontime="+70" swimtime="00:00:34.19" resultid="50522" heatid="50703" lane="2" entrytime="00:00:34.39" entrycourse="LCM" />
                <RESULT eventid="44409" points="621" reactiontime="+66" swimtime="00:01:15.16" resultid="50523" heatid="50756" lane="3" entrytime="00:01:16.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="537" reactiontime="+66" swimtime="00:00:30.05" resultid="50524" heatid="50779" lane="8" entrytime="00:00:30.06" entrycourse="LCM" />
                <RESULT eventid="46300" points="657" reactiontime="+70" swimtime="00:00:27.22" resultid="50525" heatid="50835" lane="2" entrytime="00:00:27.63" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michalina" lastname="Głowiak" birthdate="2007-03-18" gender="F" nation="POL" license="100101601444" swrid="5166102" athleteid="50478">
              <RESULTS>
                <RESULT eventid="44380" points="521" reactiontime="+72" swimtime="00:01:04.23" resultid="50479" heatid="50686" lane="5" entrytime="00:01:04.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44392" points="496" reactiontime="+72" swimtime="00:02:39.31" resultid="50480" heatid="50715" lane="5" entrytime="00:02:38.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                    <SPLIT distance="100" swimtime="00:01:17.09" />
                    <SPLIT distance="150" swimtime="00:02:02.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="512" reactiontime="+70" swimtime="00:02:21.14" resultid="50481" heatid="50743" lane="8" entrytime="00:02:20.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                    <SPLIT distance="100" swimtime="00:01:09.16" />
                    <SPLIT distance="150" swimtime="00:01:45.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="438" reactiontime="+67" swimtime="00:00:32.16" resultid="50482" heatid="50772" lane="0" />
                <RESULT eventid="46300" points="521" reactiontime="+70" swimtime="00:00:29.40" resultid="50483" heatid="50832" lane="3" entrytime="00:00:29.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Michalczuk" birthdate="2007-07-06" gender="M" nation="POL" license="100101701255" swrid="5266466" athleteid="50320">
              <RESULTS>
                <RESULT eventid="44378" points="411" reactiontime="+80" swimtime="00:01:03.05" resultid="50321" heatid="50670" lane="1" entrytime="00:01:04.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="342" reactiontime="+80" swimtime="00:02:25.78" resultid="50322" heatid="50735" lane="0" entrytime="00:02:27.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.75" />
                    <SPLIT distance="100" swimtime="00:01:09.11" />
                    <SPLIT distance="150" swimtime="00:01:48.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="341" reactiontime="+80" swimtime="00:00:31.85" resultid="50323" heatid="50763" lane="3" entrytime="00:00:33.23" entrycourse="LCM" />
                <RESULT eventid="46298" points="396" reactiontime="+71" swimtime="00:00:28.46" resultid="50324" heatid="50816" lane="0" entrytime="00:00:29.61" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Wołkowska" birthdate="2008-02-19" gender="F" nation="POL" license="100101601324" swrid="5244031" athleteid="50441">
              <RESULTS>
                <RESULT eventid="44380" points="366" reactiontime="+74" swimtime="00:01:12.27" resultid="50442" heatid="50682" lane="2" entrytime="00:01:10.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44396" points="365" reactiontime="+60" swimtime="00:01:20.50" resultid="50443" heatid="50726" lane="3" entrytime="00:01:18.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44417" points="358" reactiontime="+62" swimtime="00:02:53.71" resultid="50444" heatid="50785" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.03" />
                    <SPLIT distance="100" swimtime="00:01:25.05" />
                    <SPLIT distance="150" swimtime="00:02:10.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="400" reactiontime="+68" swimtime="00:00:32.11" resultid="50445" heatid="50827" lane="5" />
                <RESULT eventid="46312" points="403" reactiontime="+60" swimtime="00:00:36.52" resultid="50446" heatid="50907" lane="8" entrytime="00:00:36.71" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Borowiecki" birthdate="2007-07-29" gender="M" nation="POL" license="100101701284" swrid="5244090" athleteid="50389">
              <RESULTS>
                <RESULT eventid="44378" points="321" reactiontime="+88" swimtime="00:01:08.49" resultid="50390" heatid="50664" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="240" reactiontime="+75" swimtime="00:01:23.34" resultid="50391" heatid="50719" lane="2" entrytime="00:01:24.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="307" reactiontime="+91" swimtime="00:02:31.19" resultid="50392" heatid="50734" lane="7" entrytime="00:02:31.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                    <SPLIT distance="100" swimtime="00:01:12.36" />
                    <SPLIT distance="150" swimtime="00:01:53.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="308" reactiontime="+87" swimtime="00:00:30.93" resultid="50393" heatid="50810" lane="8" />
                <RESULT eventid="46310" points="253" reactiontime="+70" swimtime="00:00:37.90" resultid="50394" heatid="50855" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miłosz" lastname="Frankowski" birthdate="2005-09-03" gender="M" nation="POL" license="100101701055" swrid="4911027" athleteid="50566">
              <RESULTS>
                <RESULT eventid="44390" points="579" reactiontime="+61" swimtime="00:02:16.76" resultid="50567" heatid="50711" lane="1" entrytime="00:02:24.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.76" />
                    <SPLIT distance="100" swimtime="00:01:04.40" />
                    <SPLIT distance="150" swimtime="00:01:44.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="565" reactiontime="+48" swimtime="00:01:08.80" resultid="50568" heatid="50750" lane="4" entrytime="00:01:10.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="594" reactiontime="+58" swimtime="00:00:26.48" resultid="50569" heatid="50768" lane="3" entrytime="00:00:27.07" entrycourse="LCM" />
                <RESULT eventid="46302" points="566" reactiontime="+63" swimtime="00:02:32.44" resultid="50570" heatid="50839" lane="1" entrytime="00:02:37.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                    <SPLIT distance="100" swimtime="00:01:12.01" />
                    <SPLIT distance="150" swimtime="00:01:52.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwia" lastname="Kaniak" birthdate="2002-09-18" gender="F" nation="POL" license="100101601082" swrid="4949111" athleteid="50538">
              <RESULTS>
                <RESULT eventid="44384" points="634" reactiontime="+64" swimtime="00:00:34.22" resultid="50539" heatid="50703" lane="4" entrytime="00:00:33.43" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zofia" lastname="Urbaniak" birthdate="2008-02-02" gender="F" nation="POL" license="100101601283" swrid="5244050" athleteid="50447">
              <RESULTS>
                <RESULT eventid="44380" points="361" swimtime="00:01:12.59" resultid="50448" heatid="50682" lane="0" entrytime="00:01:11.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44384" points="255" reactiontime="+86" swimtime="00:00:46.35" resultid="50449" heatid="50700" lane="7" entrytime="00:00:44.73" entrycourse="LCM" />
                <RESULT eventid="44409" points="264" reactiontime="+82" swimtime="00:01:39.87" resultid="50450" heatid="50753" lane="7" entrytime="00:01:38.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="371" reactiontime="+81" swimtime="00:00:32.92" resultid="50451" heatid="50829" lane="2" entrytime="00:00:33.28" entrycourse="LCM" />
                <RESULT eventid="46304" points="276" swimtime="00:03:33.53" resultid="50452" heatid="50842" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.89" />
                    <SPLIT distance="100" swimtime="00:01:42.47" />
                    <SPLIT distance="150" swimtime="00:02:38.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Liwia" lastname="Bawolska" birthdate="2006-03-06" gender="F" nation="POL" license="100101601410" swrid="5166061" athleteid="50423">
              <RESULTS>
                <RESULT eventid="44380" points="511" reactiontime="+79" swimtime="00:01:04.64" resultid="50424" heatid="50686" lane="7" entrytime="00:01:04.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44392" points="458" reactiontime="+75" swimtime="00:02:43.58" resultid="50425" heatid="50715" lane="2" entrytime="00:02:41.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                    <SPLIT distance="100" swimtime="00:01:16.34" />
                    <SPLIT distance="150" swimtime="00:02:05.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="447" reactiontime="+79" swimtime="00:02:27.70" resultid="50426" heatid="50742" lane="1" entrytime="00:02:27.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                    <SPLIT distance="100" swimtime="00:01:11.30" />
                    <SPLIT distance="150" swimtime="00:01:50.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="470" reactiontime="+76" swimtime="00:00:31.40" resultid="50427" heatid="50775" lane="9" entrytime="00:00:37.77" entrycourse="LCM" />
                <RESULT eventid="46300" points="527" reactiontime="+61" swimtime="00:00:29.30" resultid="50428" heatid="50829" lane="4" entrytime="00:00:32.80" entrycourse="LCM" />
                <RESULT eventid="46312" points="444" reactiontime="+92" swimtime="00:00:35.36" resultid="50429" heatid="50906" lane="1" entrytime="00:00:40.35" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Makuszewska" birthdate="2005-12-12" gender="F" nation="POL" license="100101601133" swrid="5117240" athleteid="50471">
              <RESULTS>
                <RESULT eventid="44380" points="615" reactiontime="+67" swimtime="00:01:00.79" resultid="50472" heatid="50685" lane="3" entrytime="00:01:05.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44392" points="578" reactiontime="+67" swimtime="00:02:31.38" resultid="50473" heatid="50716" lane="7" entrytime="00:02:30.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                    <SPLIT distance="100" swimtime="00:01:11.93" />
                    <SPLIT distance="150" swimtime="00:01:55.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="577" reactiontime="+66" swimtime="00:02:15.67" resultid="50474" heatid="50744" lane="2" entrytime="00:02:12.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.69" />
                    <SPLIT distance="100" swimtime="00:01:04.99" />
                    <SPLIT distance="150" swimtime="00:01:40.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="549" reactiontime="+70" swimtime="00:00:29.82" resultid="50475" heatid="50775" lane="7" entrytime="00:00:36.48" entrycourse="LCM" />
                <RESULT eventid="46300" points="619" reactiontime="+67" swimtime="00:00:27.77" resultid="50476" heatid="50835" lane="7" entrytime="00:00:27.71" entrycourse="LCM" />
                <RESULT eventid="46308" points="514" reactiontime="+66" swimtime="00:01:09.24" resultid="50477" heatid="50901" lane="7" entrytime="00:01:08.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amelia" lastname="Władyczka" birthdate="2007-07-27" gender="F" nation="POL" license="100101601339" swrid="5272080" athleteid="50434">
              <RESULTS>
                <RESULT eventid="44380" points="580" reactiontime="+83" swimtime="00:01:02.00" resultid="50435" heatid="50687" lane="3" entrytime="00:01:02.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44396" points="520" reactiontime="+84" swimtime="00:01:11.55" resultid="50436" heatid="50728" lane="0" entrytime="00:01:11.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="561" reactiontime="+78" swimtime="00:02:16.95" resultid="50437" heatid="50743" lane="5" entrytime="00:02:16.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                    <SPLIT distance="100" swimtime="00:01:07.00" />
                    <SPLIT distance="150" swimtime="00:01:43.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44417" points="461" reactiontime="+90" swimtime="00:02:39.62" resultid="50438" heatid="50787" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                    <SPLIT distance="100" swimtime="00:01:19.20" />
                    <SPLIT distance="150" swimtime="00:02:00.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="499" reactiontime="+80" swimtime="00:04:57.93" resultid="50439" heatid="50802" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                    <SPLIT distance="100" swimtime="00:01:09.09" />
                    <SPLIT distance="150" swimtime="00:01:47.49" />
                    <SPLIT distance="200" swimtime="00:02:26.05" />
                    <SPLIT distance="250" swimtime="00:03:05.22" />
                    <SPLIT distance="300" swimtime="00:03:44.48" />
                    <SPLIT distance="350" swimtime="00:04:21.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="582" reactiontime="+78" swimtime="00:00:28.35" resultid="50440" heatid="50827" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maksym" lastname="Woźny" birthdate="2005-02-17" gender="M" nation="POL" license="100101701371" swrid="4929885" athleteid="50395">
              <RESULTS>
                <RESULT eventid="44378" points="569" reactiontime="+66" swimtime="00:00:56.59" resultid="50396" heatid="50675" lane="2" entrytime="00:00:57.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="556" reactiontime="+64" swimtime="00:02:03.98" resultid="50397" heatid="50739" lane="9" entrytime="00:02:03.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.75" />
                    <SPLIT distance="100" swimtime="00:01:00.42" />
                    <SPLIT distance="150" swimtime="00:01:32.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46285" points="553" reactiontime="+65" swimtime="00:17:40.79" resultid="50398" heatid="50790" lane="5" entrytime="00:18:02.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.17" />
                    <SPLIT distance="100" swimtime="00:01:04.37" />
                    <SPLIT distance="150" swimtime="00:01:38.80" />
                    <SPLIT distance="200" swimtime="00:02:13.47" />
                    <SPLIT distance="250" swimtime="00:02:48.00" />
                    <SPLIT distance="300" swimtime="00:03:23.43" />
                    <SPLIT distance="350" swimtime="00:03:58.62" />
                    <SPLIT distance="400" swimtime="00:04:34.11" />
                    <SPLIT distance="450" swimtime="00:05:09.44" />
                    <SPLIT distance="500" swimtime="00:05:45.23" />
                    <SPLIT distance="550" swimtime="00:06:20.95" />
                    <SPLIT distance="600" swimtime="00:06:56.90" />
                    <SPLIT distance="650" swimtime="00:07:32.77" />
                    <SPLIT distance="700" swimtime="00:08:08.47" />
                    <SPLIT distance="750" swimtime="00:08:44.28" />
                    <SPLIT distance="800" swimtime="00:09:19.98" />
                    <SPLIT distance="850" swimtime="00:09:55.73" />
                    <SPLIT distance="900" swimtime="00:10:31.84" />
                    <SPLIT distance="950" swimtime="00:11:07.73" />
                    <SPLIT distance="1000" swimtime="00:11:43.91" />
                    <SPLIT distance="1050" swimtime="00:12:19.90" />
                    <SPLIT distance="1100" swimtime="00:12:56.07" />
                    <SPLIT distance="1150" swimtime="00:13:32.14" />
                    <SPLIT distance="1200" swimtime="00:14:08.33" />
                    <SPLIT distance="1250" swimtime="00:14:44.19" />
                    <SPLIT distance="1300" swimtime="00:15:20.36" />
                    <SPLIT distance="1350" swimtime="00:15:56.38" />
                    <SPLIT distance="1400" swimtime="00:16:32.30" />
                    <SPLIT distance="1450" swimtime="00:17:07.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="567" reactiontime="+64" swimtime="00:04:25.87" resultid="50399" heatid="50800" lane="2" entrytime="00:04:20.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.08" />
                    <SPLIT distance="100" swimtime="00:01:01.66" />
                    <SPLIT distance="150" swimtime="00:01:35.56" />
                    <SPLIT distance="200" swimtime="00:02:09.88" />
                    <SPLIT distance="250" swimtime="00:02:44.43" />
                    <SPLIT distance="300" swimtime="00:03:19.20" />
                    <SPLIT distance="350" swimtime="00:03:53.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Ziemiaszewski" birthdate="2007-07-17" gender="M" nation="POL" license="100101701265" swrid="5001959" athleteid="50325">
              <RESULTS>
                <RESULT eventid="44378" points="302" reactiontime="+63" swimtime="00:01:09.85" resultid="50326" heatid="50666" lane="4" entrytime="00:01:13.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="286" reactiontime="+77" swimtime="00:01:26.24" resultid="50327" heatid="50748" lane="9" entrytime="00:01:28.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="289" reactiontime="+89" swimtime="00:00:33.65" resultid="50328" heatid="50760" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alex" lastname="Rytkowski" birthdate="2005-03-21" gender="M" nation="POL" license="100101701227" swrid="5113513" athleteid="50502">
              <RESULTS>
                <RESULT eventid="44382" points="542" reactiontime="+61" swimtime="00:00:31.81" resultid="50503" heatid="50695" lane="5" entrytime="00:00:31.40" entrycourse="LCM" />
                <RESULT eventid="44407" points="517" reactiontime="+63" swimtime="00:01:10.85" resultid="50504" heatid="50750" lane="7" entrytime="00:01:11.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="474" reactiontime="+62" swimtime="00:00:28.55" resultid="50505" heatid="50894" lane="0" entrytime="00:00:28.85" entrycourse="LCM" />
                <RESULT eventid="46298" points="484" reactiontime="+61" swimtime="00:00:26.62" resultid="50506" heatid="50820" lane="0" entrytime="00:00:26.23" entrycourse="LCM" />
                <RESULT eventid="46302" points="512" reactiontime="+65" swimtime="00:02:37.63" resultid="50507" heatid="50839" lane="3" entrytime="00:02:35.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                    <SPLIT distance="100" swimtime="00:01:14.70" />
                    <SPLIT distance="150" swimtime="00:01:56.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karol" lastname="Grudziński" birthdate="2006-03-12" gender="M" nation="POL" license="100101701403" swrid="5219616" athleteid="50349">
              <RESULTS>
                <RESULT eventid="44378" points="495" reactiontime="+65" swimtime="00:00:59.30" resultid="50350" heatid="50675" lane="3" entrytime="00:00:56.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44386" points="485" reactiontime="+71" swimtime="00:02:20.87" resultid="50351" heatid="50705" lane="1" entrytime="00:02:40.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                    <SPLIT distance="100" swimtime="00:01:09.28" />
                    <SPLIT distance="150" swimtime="00:01:46.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="406" reactiontime="+67" swimtime="00:02:17.72" resultid="50352" heatid="50738" lane="8" entrytime="00:02:10.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.46" />
                    <SPLIT distance="100" swimtime="00:01:05.60" />
                    <SPLIT distance="150" swimtime="00:01:42.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="541" reactiontime="+64" swimtime="00:00:27.33" resultid="50353" heatid="50766" lane="3" entrytime="00:00:29.23" entrycourse="LCM" />
                <RESULT eventid="46294" points="453" reactiontime="+72" swimtime="00:04:46.41" resultid="50354" heatid="50797" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                    <SPLIT distance="100" swimtime="00:01:08.73" />
                    <SPLIT distance="150" swimtime="00:01:46.36" />
                    <SPLIT distance="200" swimtime="00:02:24.66" />
                    <SPLIT distance="250" swimtime="00:03:02.62" />
                    <SPLIT distance="300" swimtime="00:03:38.68" />
                    <SPLIT distance="350" swimtime="00:04:14.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46306" points="526" reactiontime="+59" swimtime="00:01:01.29" resultid="50355" heatid="50849" lane="8" entrytime="00:01:01.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartłomiej" lastname="Maciołek" birthdate="2005-01-22" gender="M" nation="POL" license="100101701428" swrid="5024108" athleteid="50540">
              <RESULTS>
                <RESULT eventid="44386" points="486" reactiontime="+65" swimtime="00:02:20.79" resultid="50541" heatid="50705" lane="7" entrytime="00:02:30.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.88" />
                    <SPLIT distance="100" swimtime="00:01:04.03" />
                    <SPLIT distance="150" swimtime="00:01:41.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="479" reactiontime="+63" swimtime="00:00:28.46" resultid="50542" heatid="50766" lane="9" entrytime="00:00:29.78" entrycourse="LCM" />
                <RESULT eventid="44415" points="493" reactiontime="+67" swimtime="00:02:21.67" resultid="50543" heatid="50784" lane="7" entrytime="00:02:18.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.38" />
                    <SPLIT distance="100" swimtime="00:01:09.61" />
                    <SPLIT distance="150" swimtime="00:01:46.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46306" points="487" reactiontime="+65" swimtime="00:01:02.89" resultid="50544" heatid="50848" lane="4" entrytime="00:01:02.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Lech" birthdate="2005-03-22" gender="M" nation="POL" license="100101701441" swrid="5166050" athleteid="50400">
              <RESULTS>
                <RESULT eventid="44378" points="522" reactiontime="+69" swimtime="00:00:58.26" resultid="50401" heatid="50664" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="451" reactiontime="+72" swimtime="00:01:14.16" resultid="50402" heatid="50750" lane="8" entrytime="00:01:12.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46302" points="474" reactiontime="+71" swimtime="00:02:41.71" resultid="50403" heatid="50839" lane="2" entrytime="00:02:36.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.17" />
                    <SPLIT distance="100" swimtime="00:01:16.90" />
                    <SPLIT distance="150" swimtime="00:01:59.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Traczyk" birthdate="2006-06-14" gender="F" nation="POL" license="100101601203" swrid="5191060" athleteid="50571">
              <RESULTS>
                <RESULT eventid="44392" points="583" reactiontime="+77" swimtime="00:02:30.96" resultid="50572" heatid="50716" lane="1" entrytime="00:02:31.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                    <SPLIT distance="100" swimtime="00:01:09.53" />
                    <SPLIT distance="150" swimtime="00:01:55.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44396" points="550" reactiontime="+78" swimtime="00:01:10.26" resultid="50573" heatid="50728" lane="7" entrytime="00:01:09.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44417" points="605" reactiontime="+79" swimtime="00:02:25.84" resultid="50574" heatid="50786" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.36" />
                    <SPLIT distance="100" swimtime="00:01:11.57" />
                    <SPLIT distance="150" swimtime="00:01:49.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46287" points="510" reactiontime="+75" swimtime="00:10:06.58" resultid="50575" heatid="50792" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                    <SPLIT distance="100" swimtime="00:01:11.39" />
                    <SPLIT distance="150" swimtime="00:01:49.65" />
                    <SPLIT distance="200" swimtime="00:02:28.38" />
                    <SPLIT distance="250" swimtime="00:03:06.78" />
                    <SPLIT distance="300" swimtime="00:03:45.19" />
                    <SPLIT distance="350" swimtime="00:04:23.65" />
                    <SPLIT distance="400" swimtime="00:05:02.79" />
                    <SPLIT distance="450" swimtime="00:05:41.91" />
                    <SPLIT distance="500" swimtime="00:06:20.29" />
                    <SPLIT distance="550" swimtime="00:06:58.90" />
                    <SPLIT distance="600" swimtime="00:07:37.22" />
                    <SPLIT distance="650" swimtime="00:08:15.38" />
                    <SPLIT distance="700" swimtime="00:08:53.51" />
                    <SPLIT distance="750" swimtime="00:09:30.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="563" reactiontime="+73" swimtime="00:04:46.23" resultid="50576" heatid="50802" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.90" />
                    <SPLIT distance="100" swimtime="00:01:07.42" />
                    <SPLIT distance="150" swimtime="00:01:44.38" />
                    <SPLIT distance="200" swimtime="00:02:21.25" />
                    <SPLIT distance="250" swimtime="00:02:58.28" />
                    <SPLIT distance="300" swimtime="00:03:35.56" />
                    <SPLIT distance="350" swimtime="00:04:11.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46308" points="465" reactiontime="+76" swimtime="00:01:11.57" resultid="50577" heatid="50901" lane="8" entrytime="00:01:08.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrianna" lastname="Michałowska" birthdate="2008-03-01" gender="F" nation="POL" license="100101601256" swrid="5266485" athleteid="50545">
              <RESULTS>
                <RESULT eventid="44388" points="335" reactiontime="+67" swimtime="00:02:55.30" resultid="50546" heatid="50706" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.87" />
                    <SPLIT distance="100" swimtime="00:01:19.00" />
                    <SPLIT distance="150" swimtime="00:02:06.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46308" points="412" reactiontime="+74" swimtime="00:01:14.55" resultid="50547" heatid="50900" lane="1" entrytime="00:01:13.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Kramkowska" birthdate="2004-09-29" gender="F" nation="POL" license="100101601287" swrid="4990815" athleteid="50430">
              <RESULTS>
                <RESULT eventid="44380" points="587" reactiontime="+70" swimtime="00:01:01.73" resultid="50431" heatid="50687" lane="2" entrytime="00:01:02.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="596" reactiontime="+70" swimtime="00:02:14.22" resultid="50432" heatid="50744" lane="8" entrytime="00:02:14.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.39" />
                    <SPLIT distance="100" swimtime="00:01:05.38" />
                    <SPLIT distance="150" swimtime="00:01:40.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="583" reactiontime="+70" swimtime="00:00:28.33" resultid="50433" heatid="50834" lane="6" entrytime="00:00:28.25" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Malaczewska" birthdate="2005-07-05" gender="F" nation="POL" license="100101601336" swrid="5088657" athleteid="50583">
              <RESULTS>
                <RESULT eventid="44392" points="509" reactiontime="+68" swimtime="00:02:37.95" resultid="50584" heatid="50715" lane="3" entrytime="00:02:39.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                    <SPLIT distance="100" swimtime="00:01:12.98" />
                    <SPLIT distance="150" swimtime="00:02:00.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44417" points="500" reactiontime="+69" swimtime="00:02:35.39" resultid="50585" heatid="50788" lane="2" entrytime="00:02:32.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.08" />
                    <SPLIT distance="100" swimtime="00:01:15.97" />
                    <SPLIT distance="150" swimtime="00:01:55.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="585" reactiontime="+67" swimtime="00:00:28.30" resultid="50586" heatid="50833" lane="5" entrytime="00:00:29.07" entrycourse="LCM" />
                <RESULT eventid="46312" points="593" reactiontime="+62" swimtime="00:00:32.10" resultid="50587" heatid="50909" lane="8" entrytime="00:00:32.03" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Durlik" birthdate="2005-04-30" gender="M" nation="POL" license="100101701335" swrid="5118820" athleteid="50554">
              <RESULTS>
                <RESULT eventid="44390" points="486" reactiontime="+67" swimtime="00:02:24.90" resultid="50555" heatid="50711" lane="0" entrytime="00:02:26.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.37" />
                    <SPLIT distance="100" swimtime="00:01:07.77" />
                    <SPLIT distance="150" swimtime="00:01:51.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="493" reactiontime="+66" swimtime="00:02:09.06" resultid="50556" heatid="50737" lane="2" entrytime="00:02:12.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.62" />
                    <SPLIT distance="100" swimtime="00:01:01.05" />
                    <SPLIT distance="150" swimtime="00:01:35.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="533" reactiontime="+63" swimtime="00:00:27.45" resultid="50557" heatid="50768" lane="1" entrytime="00:00:27.49" entrycourse="LCM" />
                <RESULT eventid="46298" points="524" reactiontime="+62" swimtime="00:00:25.93" resultid="50558" heatid="50819" lane="6" entrytime="00:00:26.41" entrycourse="LCM" />
                <RESULT eventid="46306" points="533" reactiontime="+62" swimtime="00:01:01.03" resultid="50559" heatid="50849" lane="9" entrytime="00:01:01.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maksymilian" lastname="Czarny" birthdate="2006-09-11" gender="M" nation="POL" license="100101701401" swrid="5222193" athleteid="50490">
              <RESULTS>
                <RESULT eventid="44382" points="479" reactiontime="+59" swimtime="00:00:33.16" resultid="50491" heatid="50691" lane="6" />
                <RESULT eventid="44394" points="375" reactiontime="+70" swimtime="00:01:11.87" resultid="50492" heatid="50722" lane="4" entrytime="00:01:07.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="455" reactiontime="+66" swimtime="00:01:13.92" resultid="50493" heatid="50750" lane="0" entrytime="00:01:13.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="177" reactiontime="+95" swimtime="00:00:39.66" resultid="50494" heatid="50759" lane="9" />
                <RESULT eventid="46302" points="449" reactiontime="+65" swimtime="00:02:44.70" resultid="50495" heatid="50837" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                    <SPLIT distance="100" swimtime="00:01:20.61" />
                    <SPLIT distance="150" swimtime="00:02:03.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46310" points="375" reactiontime="+72" swimtime="00:00:33.28" resultid="50496" heatid="50858" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Strużyk" birthdate="2004-06-27" gender="F" nation="POL" license="100101601049" swrid="5072852" athleteid="50578">
              <RESULTS>
                <RESULT eventid="44392" points="557" reactiontime="+76" swimtime="00:02:33.24" resultid="50579" heatid="50716" lane="0" entrytime="00:02:34.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                    <SPLIT distance="100" swimtime="00:01:11.56" />
                    <SPLIT distance="150" swimtime="00:01:56.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44417" points="575" reactiontime="+62" swimtime="00:02:28.32" resultid="50580" heatid="50788" lane="3" entrytime="00:02:29.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                    <SPLIT distance="100" swimtime="00:01:12.23" />
                    <SPLIT distance="150" swimtime="00:01:51.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="553" reactiontime="+73" swimtime="00:04:48.08" resultid="50581" heatid="50805" lane="7" entrytime="00:04:45.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                    <SPLIT distance="100" swimtime="00:01:06.95" />
                    <SPLIT distance="150" swimtime="00:01:43.56" />
                    <SPLIT distance="200" swimtime="00:02:20.63" />
                    <SPLIT distance="250" swimtime="00:02:57.58" />
                    <SPLIT distance="300" swimtime="00:03:34.80" />
                    <SPLIT distance="350" swimtime="00:04:12.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="598" reactiontime="+59" swimtime="00:00:32.02" resultid="50582" heatid="50909" lane="7" entrytime="00:00:31.80" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Iga" lastname="Maślej" birthdate="2003-05-15" gender="F" nation="POL" license="100101601020" swrid="5043142" athleteid="50548">
              <RESULTS>
                <RESULT eventid="44388" points="447" reactiontime="+54" swimtime="00:02:39.28" resultid="50549" heatid="50706" lane="5" entrytime="00:02:36.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                    <SPLIT distance="100" swimtime="00:01:11.33" />
                    <SPLIT distance="150" swimtime="00:01:54.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="557" reactiontime="+56" swimtime="00:02:17.29" resultid="50550" heatid="50743" lane="4" entrytime="00:02:16.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                    <SPLIT distance="100" swimtime="00:01:06.71" />
                    <SPLIT distance="150" swimtime="00:01:42.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46287" points="504" reactiontime="+73" swimtime="00:10:08.92" resultid="50551" heatid="50792" lane="3" entrytime="00:10:04.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.46" />
                    <SPLIT distance="100" swimtime="00:01:12.56" />
                    <SPLIT distance="150" swimtime="00:01:51.19" />
                    <SPLIT distance="200" swimtime="00:02:30.16" />
                    <SPLIT distance="250" swimtime="00:03:08.91" />
                    <SPLIT distance="300" swimtime="00:03:47.63" />
                    <SPLIT distance="350" swimtime="00:04:26.23" />
                    <SPLIT distance="400" swimtime="00:05:04.79" />
                    <SPLIT distance="450" swimtime="00:05:43.30" />
                    <SPLIT distance="500" swimtime="00:06:21.44" />
                    <SPLIT distance="550" swimtime="00:06:59.73" />
                    <SPLIT distance="600" swimtime="00:07:37.85" />
                    <SPLIT distance="650" swimtime="00:08:15.95" />
                    <SPLIT distance="700" swimtime="00:08:54.26" />
                    <SPLIT distance="750" swimtime="00:09:32.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="537" reactiontime="+69" swimtime="00:04:50.88" resultid="50552" heatid="50805" lane="8" entrytime="00:04:49.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                    <SPLIT distance="100" swimtime="00:01:08.35" />
                    <SPLIT distance="150" swimtime="00:01:45.28" />
                    <SPLIT distance="200" swimtime="00:02:22.18" />
                    <SPLIT distance="250" swimtime="00:02:59.44" />
                    <SPLIT distance="300" swimtime="00:03:37.23" />
                    <SPLIT distance="350" swimtime="00:04:14.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46308" points="516" reactiontime="+61" swimtime="00:01:09.16" resultid="50553" heatid="50901" lane="0" entrytime="00:01:09.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Maciuszek" birthdate="2004-05-11" gender="F" nation="POL" license="100101601407" swrid="4858842" athleteid="50466">
              <RESULTS>
                <RESULT eventid="44380" points="683" reactiontime="+64" swimtime="00:00:58.69" resultid="50467" heatid="50688" lane="5" entrytime="00:00:58.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44396" points="607" reactiontime="+59" swimtime="00:01:07.99" resultid="50468" heatid="50728" lane="3" entrytime="00:01:04.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="659" reactiontime="+65" swimtime="00:00:27.19" resultid="50469" heatid="50835" lane="6" entrytime="00:00:27.19" entrycourse="LCM" />
                <RESULT eventid="46312" points="676" reactiontime="+57" swimtime="00:00:30.74" resultid="50470" heatid="50909" lane="2" entrytime="00:00:30.56" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leon" lastname="Bednorz" birthdate="2008-08-13" gender="M" nation="POL" license="100101701291" swrid="5318117" athleteid="50383">
              <RESULTS>
                <RESULT eventid="44378" points="265" reactiontime="+53" swimtime="00:01:12.97" resultid="50384" heatid="50666" lane="5" entrytime="00:01:14.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="191" reactiontime="+54" swimtime="00:00:45.04" resultid="50385" heatid="50692" lane="5" entrytime="00:00:46.98" entrycourse="LCM" />
                <RESULT eventid="44407" points="205" reactiontime="+73" swimtime="00:01:36.39" resultid="50386" heatid="50747" lane="1" entrytime="00:01:38.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="157" reactiontime="+67" swimtime="00:00:41.20" resultid="50387" heatid="50762" lane="8" entrytime="00:00:45.53" entrycourse="LCM" />
                <RESULT eventid="46298" points="234" reactiontime="+53" swimtime="00:00:33.89" resultid="50388" heatid="50813" lane="0" entrytime="00:00:34.82" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Kędzia" birthdate="2007-06-06" gender="M" nation="POL" license="100101701249" swrid="5266462" athleteid="50329">
              <RESULTS>
                <RESULT eventid="44378" points="327" reactiontime="+76" swimtime="00:01:08.05" resultid="50330" heatid="50668" lane="1" entrytime="00:01:07.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="319" reactiontime="+83" swimtime="00:02:29.23" resultid="50331" heatid="50734" lane="1" entrytime="00:02:31.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                    <SPLIT distance="100" swimtime="00:01:14.02" />
                    <SPLIT distance="150" swimtime="00:01:53.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46285" points="346" reactiontime="+83" swimtime="00:20:40.30" resultid="50332" heatid="50790" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                    <SPLIT distance="100" swimtime="00:01:15.25" />
                    <SPLIT distance="150" swimtime="00:01:56.17" />
                    <SPLIT distance="200" swimtime="00:02:36.77" />
                    <SPLIT distance="250" swimtime="00:03:18.05" />
                    <SPLIT distance="300" swimtime="00:03:59.81" />
                    <SPLIT distance="350" swimtime="00:04:41.96" />
                    <SPLIT distance="400" swimtime="00:05:23.94" />
                    <SPLIT distance="450" swimtime="00:06:06.07" />
                    <SPLIT distance="500" swimtime="00:06:48.55" />
                    <SPLIT distance="550" swimtime="00:07:32.31" />
                    <SPLIT distance="600" swimtime="00:08:13.83" />
                    <SPLIT distance="650" swimtime="00:08:56.36" />
                    <SPLIT distance="700" swimtime="00:09:39.74" />
                    <SPLIT distance="750" swimtime="00:10:20.43" />
                    <SPLIT distance="800" swimtime="00:11:03.51" />
                    <SPLIT distance="850" swimtime="00:11:45.70" />
                    <SPLIT distance="900" swimtime="00:12:27.88" />
                    <SPLIT distance="950" swimtime="00:13:09.90" />
                    <SPLIT distance="1000" swimtime="00:13:52.26" />
                    <SPLIT distance="1050" swimtime="00:14:34.21" />
                    <SPLIT distance="1100" swimtime="00:15:15.60" />
                    <SPLIT distance="1150" swimtime="00:15:57.39" />
                    <SPLIT distance="1200" swimtime="00:16:40.51" />
                    <SPLIT distance="1250" swimtime="00:17:22.34" />
                    <SPLIT distance="1300" swimtime="00:18:02.88" />
                    <SPLIT distance="1350" swimtime="00:18:43.38" />
                    <SPLIT distance="1400" swimtime="00:19:23.64" />
                    <SPLIT distance="1450" swimtime="00:20:02.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="324" reactiontime="+83" swimtime="00:05:20.34" resultid="50333" heatid="50797" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                    <SPLIT distance="100" swimtime="00:01:14.10" />
                    <SPLIT distance="150" swimtime="00:01:54.89" />
                    <SPLIT distance="200" swimtime="00:02:36.33" />
                    <SPLIT distance="250" swimtime="00:03:18.30" />
                    <SPLIT distance="300" swimtime="00:04:00.80" />
                    <SPLIT distance="350" swimtime="00:04:41.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46306" points="185" reactiontime="+83" swimtime="00:01:26.79" resultid="50334" heatid="50844" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leon" lastname="Fischer" birthdate="2007-04-14" gender="M" nation="POL" license="100101701277" swrid="5136358" athleteid="50362">
              <RESULTS>
                <RESULT eventid="44378" points="478" reactiontime="+86" swimtime="00:00:59.96" resultid="50363" heatid="50665" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="359" reactiontime="+78" swimtime="00:00:36.49" resultid="50364" heatid="50692" lane="2" entrytime="00:00:48.40" entrycourse="LCM" />
                <RESULT eventid="44407" points="317" reactiontime="+85" swimtime="00:01:23.35" resultid="50365" heatid="50748" lane="2" entrytime="00:01:25.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="349" reactiontime="+86" swimtime="00:00:31.61" resultid="50366" heatid="50760" lane="0" />
                <RESULT eventid="46298" points="420" reactiontime="+75" swimtime="00:00:27.92" resultid="50367" heatid="50811" lane="4" entrytime="00:00:44.12" entrycourse="LCM" />
                <RESULT eventid="46302" points="340" reactiontime="+82" swimtime="00:03:00.65" resultid="50368" heatid="50836" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.60" />
                    <SPLIT distance="100" swimtime="00:01:26.31" />
                    <SPLIT distance="150" swimtime="00:02:13.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Dyrda" birthdate="2006-04-26" gender="M" nation="POL" license="100101701402" swrid="5219618" athleteid="50342">
              <RESULTS>
                <RESULT eventid="44378" points="502" reactiontime="+71" swimtime="00:00:59.00" resultid="50343" heatid="50673" lane="4" entrytime="00:00:59.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="492" reactiontime="+70" swimtime="00:01:05.67" resultid="50344" heatid="50723" lane="1" entrytime="00:01:05.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="385" reactiontime="+79" swimtime="00:00:30.60" resultid="50345" heatid="50757" lane="3" />
                <RESULT eventid="44415" points="382" reactiontime="+82" swimtime="00:02:34.13" resultid="50346" heatid="50781" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                    <SPLIT distance="100" swimtime="00:01:15.46" />
                    <SPLIT distance="150" swimtime="00:01:56.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="467" reactiontime="+71" swimtime="00:00:26.95" resultid="50347" heatid="50811" lane="9" />
                <RESULT eventid="46310" points="516" reactiontime="+71" swimtime="00:00:29.92" resultid="50348" heatid="50856" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Klaudia" lastname="Naziębło" birthdate="1993-12-03" gender="F" nation="POL" license="100101600997" swrid="4087213" athleteid="50881">
              <RESULTS>
                <RESULT eventid="46308" points="828" reactiontime="+69" swimtime="00:00:59.06" resultid="50882" heatid="50901" lane="4" late="yes" entrytime="00:00:59.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="856" reactiontime="+55" swimtime="00:00:28.41" resultid="50883" heatid="50909" lane="4" entrytime="00:00:28.60" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Leśniak" birthdate="2008-03-20" gender="F" nation="POL" license="100101601296" swrid="5244041" athleteid="50453">
              <RESULTS>
                <RESULT eventid="44380" points="283" reactiontime="+88" swimtime="00:01:18.71" resultid="50454" heatid="50681" lane="2" entrytime="00:01:15.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44396" points="286" reactiontime="+95" swimtime="00:01:27.30" resultid="50455" heatid="50726" lane="9" entrytime="00:01:24.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44417" points="302" reactiontime="+86" swimtime="00:03:03.75" resultid="50456" heatid="50786" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.56" />
                    <SPLIT distance="100" swimtime="00:01:31.21" />
                    <SPLIT distance="150" swimtime="00:02:17.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="291" reactiontime="+89" swimtime="00:00:35.68" resultid="50457" heatid="50829" lane="0" entrytime="00:00:34.45" entrycourse="LCM" />
                <RESULT eventid="46312" points="302" reactiontime="+71" swimtime="00:00:40.19" resultid="50458" heatid="50906" lane="9" entrytime="00:00:42.06" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Zakrzewska" birthdate="2003-01-29" gender="F" nation="POL" license="100101601297" swrid="4911016" athleteid="50515">
              <RESULTS>
                <RESULT eventid="44384" points="546" reactiontime="+66" swimtime="00:00:35.97" resultid="50516" heatid="50702" lane="5" entrytime="00:00:35.70" entrycourse="LCM" />
                <RESULT eventid="44396" points="567" reactiontime="+61" swimtime="00:01:09.52" resultid="50517" heatid="50728" lane="1" entrytime="00:01:09.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44417" points="564" reactiontime="+61" swimtime="00:02:29.27" resultid="50518" heatid="50788" lane="7" entrytime="00:02:33.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                    <SPLIT distance="100" swimtime="00:01:12.21" />
                    <SPLIT distance="150" swimtime="00:01:50.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="587" reactiontime="+66" swimtime="00:00:28.26" resultid="50519" heatid="50834" lane="5" entrytime="00:00:28.08" entrycourse="LCM" />
                <RESULT eventid="46312" points="601" reactiontime="+60" swimtime="00:00:31.97" resultid="50520" heatid="50909" lane="1" entrytime="00:00:31.92" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Kochańska" birthdate="2008-04-11" gender="F" nation="POL" license="100101601299" swrid="4838369" athleteid="50526">
              <RESULTS>
                <RESULT eventid="44384" points="421" reactiontime="+67" swimtime="00:00:39.21" resultid="50527" heatid="50701" lane="7" entrytime="00:00:41.27" entrycourse="LCM" />
                <RESULT eventid="44392" points="362" reactiontime="+53" swimtime="00:02:56.92" resultid="50528" heatid="50714" lane="0" entrytime="00:02:53.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                    <SPLIT distance="100" swimtime="00:01:28.01" />
                    <SPLIT distance="150" swimtime="00:02:17.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44409" points="382" reactiontime="+65" swimtime="00:01:28.34" resultid="50529" heatid="50754" lane="6" entrytime="00:01:25.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="402" reactiontime="+62" swimtime="00:05:20.31" resultid="50530" heatid="50803" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.53" />
                    <SPLIT distance="100" swimtime="00:01:16.46" />
                    <SPLIT distance="150" swimtime="00:01:57.88" />
                    <SPLIT distance="200" swimtime="00:02:39.12" />
                    <SPLIT distance="250" swimtime="00:03:20.78" />
                    <SPLIT distance="300" swimtime="00:04:01.91" />
                    <SPLIT distance="350" swimtime="00:04:43.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="374" reactiontime="+64" swimtime="00:00:32.85" resultid="50531" heatid="50830" lane="7" entrytime="00:00:31.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Sarnowicz" birthdate="2004-03-01" gender="M" nation="POL" license="100101701073" swrid="5118745" athleteid="50497">
              <RESULTS>
                <RESULT eventid="44382" points="555" reactiontime="+63" swimtime="00:00:31.57" resultid="50498" heatid="50695" lane="4" entrytime="00:00:31.22" entrycourse="LCM" />
                <RESULT eventid="44407" points="512" reactiontime="+63" swimtime="00:01:11.10" resultid="50499" heatid="50750" lane="3" entrytime="00:01:10.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="494" reactiontime="+63" swimtime="00:00:26.45" resultid="50500" heatid="50819" lane="9" entrytime="00:00:26.67" entrycourse="LCM" />
                <RESULT eventid="46302" points="486" reactiontime="+67" swimtime="00:02:40.33" resultid="50501" heatid="50839" lane="6" entrytime="00:02:36.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                    <SPLIT distance="100" swimtime="00:01:15.10" />
                    <SPLIT distance="150" swimtime="00:01:56.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oskar" lastname="Nowak" birthdate="2006-03-22" gender="M" nation="POL" license="100101701178" swrid="4834359" athleteid="50356">
              <RESULTS>
                <RESULT eventid="44378" points="460" reactiontime="+82" swimtime="00:01:00.74" resultid="50357" heatid="50673" lane="8" entrytime="00:01:00.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="365" reactiontime="+76" swimtime="00:01:12.49" resultid="50358" heatid="50721" lane="1" entrytime="00:01:15.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="434" reactiontime="+80" swimtime="00:02:14.67" resultid="50359" heatid="50736" lane="1" entrytime="00:02:17.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.20" />
                    <SPLIT distance="100" swimtime="00:01:05.19" />
                    <SPLIT distance="150" swimtime="00:01:41.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="447" reactiontime="+75" swimtime="00:04:47.81" resultid="50360" heatid="50797" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                    <SPLIT distance="100" swimtime="00:01:08.05" />
                    <SPLIT distance="150" swimtime="00:01:45.92" />
                    <SPLIT distance="200" swimtime="00:02:23.46" />
                    <SPLIT distance="250" swimtime="00:03:00.93" />
                    <SPLIT distance="300" swimtime="00:03:38.36" />
                    <SPLIT distance="350" swimtime="00:04:15.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="431" reactiontime="+77" swimtime="00:00:27.67" resultid="50361" heatid="50812" lane="5" entrytime="00:00:35.66" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="95" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="44399" points="565" reactiontime="+65" swimtime="00:04:10.61" resultid="47530" heatid="50730" lane="6" entrytime="00:04:12.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.06" />
                    <SPLIT distance="100" swimtime="00:01:03.52" />
                    <SPLIT distance="150" swimtime="00:01:35.56" />
                    <SPLIT distance="200" swimtime="00:02:12.16" />
                    <SPLIT distance="250" swimtime="00:02:40.29" />
                    <SPLIT distance="300" swimtime="00:03:13.69" />
                    <SPLIT distance="350" swimtime="00:03:41.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="50540" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="50566" number="2" reactiontime="+11" />
                    <RELAYPOSITION athleteid="50554" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="50395" number="4" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46314" points="594" reactiontime="+47" swimtime="00:08:17.65" resultid="50608" heatid="50870" lane="4" entrytime="00:08:13.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.33" />
                    <SPLIT distance="100" swimtime="00:00:57.92" />
                    <SPLIT distance="150" swimtime="00:01:30.71" />
                    <SPLIT distance="200" swimtime="00:02:03.53" />
                    <SPLIT distance="250" swimtime="00:02:31.62" />
                    <SPLIT distance="300" swimtime="00:03:03.28" />
                    <SPLIT distance="350" swimtime="00:03:37.43" />
                    <SPLIT distance="400" swimtime="00:04:09.62" />
                    <SPLIT distance="450" swimtime="00:04:38.73" />
                    <SPLIT distance="500" swimtime="00:05:11.44" />
                    <SPLIT distance="550" swimtime="00:05:46.20" />
                    <SPLIT distance="600" swimtime="00:06:17.22" />
                    <SPLIT distance="650" swimtime="00:06:44.38" />
                    <SPLIT distance="700" swimtime="00:07:14.89" />
                    <SPLIT distance="750" swimtime="00:07:47.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="50566" number="1" reactiontime="+47" />
                    <RELAYPOSITION athleteid="50560" number="2" reactiontime="+13" />
                    <RELAYPOSITION athleteid="50540" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="50593" number="4" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="44399" points="480" reactiontime="+73" swimtime="00:04:24.69" resultid="50598" heatid="50730" lane="5" entrytime="00:04:10.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                    <SPLIT distance="100" swimtime="00:01:08.04" />
                    <SPLIT distance="150" swimtime="00:01:42.38" />
                    <SPLIT distance="200" swimtime="00:02:22.59" />
                    <SPLIT distance="250" swimtime="00:02:50.44" />
                    <SPLIT distance="300" swimtime="00:03:24.17" />
                    <SPLIT distance="350" swimtime="00:03:52.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="50342" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="50490" number="2" reactiontime="+45" />
                    <RELAYPOSITION athleteid="50349" number="3" reactiontime="+21" />
                    <RELAYPOSITION athleteid="50356" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="95" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="46289" points="594" reactiontime="+64" swimtime="00:03:43.83" resultid="50603" heatid="50794" lane="5" entrytime="00:03:39.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.99" />
                    <SPLIT distance="100" swimtime="00:00:54.21" />
                    <SPLIT distance="150" swimtime="00:01:19.94" />
                    <SPLIT distance="200" swimtime="00:01:48.57" />
                    <SPLIT distance="250" swimtime="00:02:15.58" />
                    <SPLIT distance="300" swimtime="00:02:45.46" />
                    <SPLIT distance="350" swimtime="00:03:12.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="50593" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="50404" number="2" reactiontime="+6" />
                    <RELAYPOSITION athleteid="50554" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="50497" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="95" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="46289" points="557" reactiontime="+70" swimtime="00:03:48.75" resultid="50604" heatid="50794" lane="3" entrytime="00:03:45.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.31" />
                    <SPLIT distance="100" swimtime="00:00:57.20" />
                    <SPLIT distance="150" swimtime="00:01:24.75" />
                    <SPLIT distance="200" swimtime="00:01:56.05" />
                    <SPLIT distance="250" swimtime="00:02:23.55" />
                    <SPLIT distance="300" swimtime="00:02:54.20" />
                    <SPLIT distance="350" swimtime="00:03:19.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="50560" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="50395" number="2" reactiontime="+9" />
                    <RELAYPOSITION athleteid="50540" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="50566" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="46289" points="493" reactiontime="+72" swimtime="00:03:58.20" resultid="50662" heatid="50794" lane="2" entrytime="00:03:52.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.97" />
                    <SPLIT distance="100" swimtime="00:00:59.48" />
                    <SPLIT distance="150" swimtime="00:01:27.92" />
                    <SPLIT distance="200" swimtime="00:02:00.15" />
                    <SPLIT distance="250" swimtime="00:02:28.91" />
                    <SPLIT distance="300" swimtime="00:03:00.85" />
                    <SPLIT distance="350" swimtime="00:03:28.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="50342" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="50490" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="50356" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="50349" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="95" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="44401" points="543" reactiontime="+63" swimtime="00:04:42.36" resultid="50599" heatid="50731" lane="5" entrytime="00:04:26.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                    <SPLIT distance="100" swimtime="00:01:09.05" />
                    <SPLIT distance="150" swimtime="00:01:45.99" />
                    <SPLIT distance="200" swimtime="00:02:28.87" />
                    <SPLIT distance="250" swimtime="00:02:59.99" />
                    <SPLIT distance="300" swimtime="00:03:38.83" />
                    <SPLIT distance="350" swimtime="00:04:08.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="50578" number="1" reactiontime="+63" />
                    <RELAYPOSITION athleteid="50588" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="50430" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="50548" number="4" reactiontime="+16" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46291" points="622" reactiontime="+65" swimtime="00:04:05.94" resultid="50605" heatid="50795" lane="5" entrytime="00:04:00.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.76" />
                    <SPLIT distance="100" swimtime="00:00:59.08" />
                    <SPLIT distance="150" swimtime="00:01:28.57" />
                    <SPLIT distance="200" swimtime="00:02:00.91" />
                    <SPLIT distance="250" swimtime="00:02:30.46" />
                    <SPLIT distance="300" swimtime="00:03:03.91" />
                    <SPLIT distance="350" swimtime="00:03:32.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="50588" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="50430" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="50578" number="3" reactiontime="+25" />
                    <RELAYPOSITION athleteid="50515" number="4" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46316" points="616" reactiontime="+52" swimtime="00:09:02.23" resultid="50609" heatid="50871" lane="4" entrytime="00:08:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                    <SPLIT distance="100" swimtime="00:01:06.12" />
                    <SPLIT distance="150" swimtime="00:01:40.94" />
                    <SPLIT distance="200" swimtime="00:02:14.35" />
                    <SPLIT distance="250" swimtime="00:02:44.01" />
                    <SPLIT distance="300" swimtime="00:03:18.26" />
                    <SPLIT distance="350" swimtime="00:03:53.62" />
                    <SPLIT distance="400" swimtime="00:04:28.61" />
                    <SPLIT distance="450" swimtime="00:05:01.32" />
                    <SPLIT distance="500" swimtime="00:05:37.40" />
                    <SPLIT distance="550" swimtime="00:06:14.13" />
                    <SPLIT distance="600" swimtime="00:06:49.60" />
                    <SPLIT distance="650" swimtime="00:07:20.33" />
                    <SPLIT distance="700" swimtime="00:07:54.70" />
                    <SPLIT distance="750" swimtime="00:08:29.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="50521" number="1" reactiontime="+52" />
                    <RELAYPOSITION athleteid="50471" number="2" reactiontime="+8" />
                    <RELAYPOSITION athleteid="50583" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="50484" number="4" reactiontime="+13" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="95" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="44401" points="598" reactiontime="+63" swimtime="00:04:33.41" resultid="50600" heatid="50731" lane="4" entrytime="00:04:22.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                    <SPLIT distance="100" swimtime="00:01:10.01" />
                    <SPLIT distance="150" swimtime="00:01:44.51" />
                    <SPLIT distance="200" swimtime="00:02:23.95" />
                    <SPLIT distance="250" swimtime="00:02:54.79" />
                    <SPLIT distance="300" swimtime="00:03:32.90" />
                    <SPLIT distance="350" swimtime="00:04:02.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="50583" number="1" reactiontime="+63" />
                    <RELAYPOSITION athleteid="50521" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="50471" number="3" reactiontime="+23" />
                    <RELAYPOSITION athleteid="50484" number="4" reactiontime="-10" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46291" points="649" reactiontime="+54" swimtime="00:04:02.54" resultid="50606" heatid="50795" lane="4" entrytime="00:03:55.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.06" />
                    <SPLIT distance="100" swimtime="00:01:03.16" />
                    <SPLIT distance="150" swimtime="00:01:32.37" />
                    <SPLIT distance="200" swimtime="00:02:03.60" />
                    <SPLIT distance="250" swimtime="00:02:31.58" />
                    <SPLIT distance="300" swimtime="00:03:02.89" />
                    <SPLIT distance="350" swimtime="00:03:31.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="50583" number="1" reactiontime="+54" />
                    <RELAYPOSITION athleteid="50484" number="2" reactiontime="+20" />
                    <RELAYPOSITION athleteid="50521" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="50471" number="4" reactiontime="+16" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="F" number="3">
              <RESULTS>
                <RESULT eventid="44401" points="481" reactiontime="+78" swimtime="00:04:53.92" resultid="50601" heatid="50731" lane="3" entrytime="00:04:42.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                    <SPLIT distance="100" swimtime="00:01:11.25" />
                    <SPLIT distance="150" swimtime="00:01:51.49" />
                    <SPLIT distance="200" swimtime="00:02:36.70" />
                    <SPLIT distance="250" swimtime="00:03:09.32" />
                    <SPLIT distance="300" swimtime="00:03:48.43" />
                    <SPLIT distance="350" swimtime="00:04:18.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="50571" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="50508" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="50409" number="3" reactiontime="+26" />
                    <RELAYPOSITION athleteid="50423" number="4" reactiontime="+18" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46291" points="526" reactiontime="+82" swimtime="00:04:20.19" resultid="50607" heatid="50795" lane="3" entrytime="00:04:16.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                    <SPLIT distance="100" swimtime="00:01:02.77" />
                    <SPLIT distance="150" swimtime="00:01:34.03" />
                    <SPLIT distance="200" swimtime="00:02:07.73" />
                    <SPLIT distance="250" swimtime="00:02:40.51" />
                    <SPLIT distance="300" swimtime="00:03:17.00" />
                    <SPLIT distance="350" swimtime="00:03:46.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="50434" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="50409" number="2" reactiontime="+27" />
                    <RELAYPOSITION athleteid="50416" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="50423" number="4" reactiontime="+18" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="03401" nation="POL" region="01" clubid="48489" name="UKS PATOMSWIM Bogatynia">
          <ATHLETES>
            <ATHLETE firstname="Julia" lastname="Kameduła" birthdate="2007-02-10" gender="F" nation="POL" license="103401600030" swrid="5190421" athleteid="48543">
              <RESULTS>
                <RESULT eventid="44384" points="290" reactiontime="+81" swimtime="00:00:44.38" resultid="48544" heatid="50697" lane="7" />
                <RESULT eventid="44409" points="257" reactiontime="+79" swimtime="00:01:40.74" resultid="48545" heatid="50752" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="185" reactiontime="+77" swimtime="00:00:42.81" resultid="48546" heatid="50773" lane="7" />
                <RESULT eventid="46300" points="270" reactiontime="+86" swimtime="00:00:36.60" resultid="48547" heatid="50828" lane="0" />
                <RESULT eventid="46304" points="262" reactiontime="+64" swimtime="00:03:37.22" resultid="48548" heatid="50840" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.44" />
                    <SPLIT distance="100" swimtime="00:01:44.21" />
                    <SPLIT distance="150" swimtime="00:02:42.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" status="DNS" swimtime="00:00:00.00" resultid="48549" heatid="50904" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Listkiewicz" birthdate="2006-08-04" gender="F" nation="POL" license="103401600027" swrid="5173443" athleteid="48535">
              <RESULTS>
                <RESULT eventid="44380" points="381" reactiontime="+72" swimtime="00:01:11.31" resultid="48536" heatid="50679" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44396" points="392" reactiontime="+53" swimtime="00:01:18.65" resultid="48537" heatid="50724" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" status="DNS" swimtime="00:00:00.00" resultid="48538" heatid="50773" lane="1" />
                <RESULT eventid="44417" points="350" reactiontime="+63" swimtime="00:02:54.97" resultid="48539" heatid="50786" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.63" />
                    <SPLIT distance="100" swimtime="00:01:25.68" />
                    <SPLIT distance="150" swimtime="00:02:11.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="400" reactiontime="+68" swimtime="00:00:32.10" resultid="48540" heatid="50825" lane="2" />
                <RESULT eventid="46308" points="326" reactiontime="+54" swimtime="00:01:20.53" resultid="48541" heatid="50897" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="416" reactiontime="+63" swimtime="00:00:36.12" resultid="48542" heatid="50903" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martyna" lastname="Fuławka" birthdate="2008-04-21" gender="F" nation="POL" license="103401600022" swrid="5173436" athleteid="48517">
              <RESULTS>
                <RESULT eventid="44380" points="317" reactiontime="+69" swimtime="00:01:15.76" resultid="48518" heatid="50678" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44384" points="328" reactiontime="+69" swimtime="00:00:42.61" resultid="48519" heatid="50698" lane="7" />
                <RESULT eventid="44392" points="274" reactiontime="+71" swimtime="00:03:14.07" resultid="48520" heatid="50713" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.09" />
                    <SPLIT distance="100" swimtime="00:01:33.86" />
                    <SPLIT distance="150" swimtime="00:02:31.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44396" points="262" reactiontime="+65" swimtime="00:01:29.86" resultid="48521" heatid="50724" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44409" points="275" reactiontime="+68" swimtime="00:01:38.54" resultid="48522" heatid="50751" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="290" reactiontime="+71" swimtime="00:00:36.89" resultid="48523" heatid="50771" lane="0" />
                <RESULT eventid="44417" status="DNS" swimtime="00:00:00.00" resultid="48524" heatid="50785" lane="7" />
                <RESULT eventid="46300" points="353" reactiontime="+57" swimtime="00:00:33.47" resultid="48525" heatid="50825" lane="4" />
                <RESULT eventid="46308" points="171" reactiontime="+69" swimtime="00:01:39.83" resultid="48526" heatid="50897" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="288" reactiontime="+62" swimtime="00:00:40.81" resultid="48527" heatid="50903" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Polak" birthdate="2006-01-21" gender="F" nation="POL" license="103401600026" swrid="4941793" athleteid="48528">
              <RESULTS>
                <RESULT eventid="44380" points="440" reactiontime="+58" swimtime="00:01:07.96" resultid="48529" heatid="50678" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44392" points="320" reactiontime="+76" swimtime="00:03:04.21" resultid="48530" heatid="50713" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                    <SPLIT distance="100" swimtime="00:01:24.57" />
                    <SPLIT distance="150" swimtime="00:02:20.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="398" reactiontime="+71" swimtime="00:00:33.19" resultid="48531" heatid="50770" lane="3" />
                <RESULT eventid="46300" points="508" reactiontime="+72" swimtime="00:00:29.65" resultid="48532" heatid="50825" lane="8" />
                <RESULT eventid="46308" points="314" reactiontime="+74" swimtime="00:01:21.60" resultid="48533" heatid="50897" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" status="DNS" swimtime="00:00:00.00" resultid="48534" heatid="50902" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksander" lastname="Peremicki" birthdate="2007-12-18" gender="M" nation="POL" license="103401700031" swrid="5081222" athleteid="48501">
              <RESULTS>
                <RESULT eventid="44378" points="423" reactiontime="+68" swimtime="00:01:02.45" resultid="48502" heatid="50663" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="507" reactiontime="+67" swimtime="00:00:32.54" resultid="48503" heatid="50691" lane="8" />
                <RESULT eventid="44390" status="DNS" swimtime="00:00:00.00" resultid="48504" heatid="50708" lane="1" />
                <RESULT eventid="44407" points="462" reactiontime="+65" swimtime="00:01:13.54" resultid="48505" heatid="50746" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="323" reactiontime="+64" swimtime="00:00:32.45" resultid="48506" heatid="50761" lane="9" />
                <RESULT eventid="46298" points="412" reactiontime="+63" swimtime="00:00:28.08" resultid="48507" heatid="50808" lane="9" />
                <RESULT eventid="46302" points="398" reactiontime="+69" swimtime="00:02:51.43" resultid="48508" heatid="50838" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.48" />
                    <SPLIT distance="100" swimtime="00:01:21.85" />
                    <SPLIT distance="150" swimtime="00:02:07.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46310" points="303" reactiontime="+73" swimtime="00:00:35.73" resultid="48509" heatid="50856" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Kołodziej" birthdate="2007-05-05" gender="M" nation="POL" license="103401700025" swrid="5081224" athleteid="48490">
              <RESULTS>
                <RESULT eventid="44378" points="375" reactiontime="+67" swimtime="00:01:05.04" resultid="48491" heatid="50664" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44390" points="367" reactiontime="+64" swimtime="00:02:39.13" resultid="48492" heatid="50708" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                    <SPLIT distance="100" swimtime="00:01:15.13" />
                    <SPLIT distance="150" swimtime="00:02:02.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="333" reactiontime="+62" swimtime="00:01:14.80" resultid="48493" heatid="50719" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" status="DNS" swimtime="00:00:00.00" resultid="48494" heatid="50732" lane="3" />
                <RESULT eventid="44411" points="341" reactiontime="+59" swimtime="00:00:31.85" resultid="48495" heatid="50760" lane="8" />
                <RESULT eventid="44415" points="321" reactiontime="+61" swimtime="00:02:43.42" resultid="48496" heatid="50781" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.76" />
                    <SPLIT distance="100" swimtime="00:01:19.74" />
                    <SPLIT distance="150" swimtime="00:02:02.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="352" reactiontime="+66" swimtime="00:05:11.48" resultid="48497" heatid="50797" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                    <SPLIT distance="100" swimtime="00:01:10.71" />
                    <SPLIT distance="150" swimtime="00:01:50.41" />
                    <SPLIT distance="200" swimtime="00:02:31.43" />
                    <SPLIT distance="250" swimtime="00:03:12.67" />
                    <SPLIT distance="300" swimtime="00:03:53.84" />
                    <SPLIT distance="350" swimtime="00:04:34.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="351" reactiontime="+52" swimtime="00:00:29.63" resultid="48498" heatid="50809" lane="9" />
                <RESULT eventid="46306" points="278" reactiontime="+63" swimtime="00:01:15.83" resultid="48499" heatid="50845" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46310" points="340" reactiontime="+68" swimtime="00:00:34.38" resultid="48500" heatid="50858" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Poźniak" birthdate="2008-02-29" gender="M" nation="POL" license="103401700024" swrid="5287582" athleteid="48510">
              <RESULTS>
                <RESULT eventid="44378" points="198" reactiontime="+65" swimtime="00:01:20.43" resultid="48511" heatid="50665" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="174" reactiontime="+72" swimtime="00:01:32.75" resultid="48512" heatid="50717" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="144" reactiontime="+55" swimtime="00:00:42.41" resultid="48513" heatid="50761" lane="0" />
                <RESULT eventid="46298" points="210" reactiontime="+47" swimtime="00:00:35.13" resultid="48514" heatid="50811" lane="0" />
                <RESULT eventid="46306" status="DNS" swimtime="00:00:00.00" resultid="48515" heatid="50845" lane="7" />
                <RESULT eventid="46310" points="181" reactiontime="+86" swimtime="00:00:42.38" resultid="48516" heatid="50856" lane="7" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="05114" nation="POL" region="14" clubid="48199" name="UKS G-8 Bielany Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Jakub" lastname="Kotarski" birthdate="2001-05-07" gender="M" nation="POL" license="105114700823" swrid="5019900" athleteid="48200">
              <RESULTS>
                <RESULT eventid="44378" points="654" reactiontime="+70" swimtime="00:00:54.04" resultid="48201" heatid="50676" lane="7" entrytime="00:00:55.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="565" reactiontime="+72" swimtime="00:00:25.29" resultid="48202" heatid="50820" lane="3" entrytime="00:00:26.02" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02001" nation="POL" region="01" clubid="46855" name="KS Rekin Świebodzice">
          <ATHLETES>
            <ATHLETE firstname="Jakub" lastname="Gadacz" birthdate="2006-09-04" gender="M" nation="POL" license="102001700177" swrid="5165957" athleteid="46863">
              <RESULTS>
                <RESULT eventid="44378" points="384" reactiontime="+46" swimtime="00:01:04.51" resultid="46864" heatid="50670" lane="4" entrytime="00:01:03.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="306" reactiontime="+65" swimtime="00:00:33.04" resultid="46865" heatid="50762" lane="0" entrytime="00:00:47.84" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Gajdowska" birthdate="1995-07-17" gender="F" nation="POL" license="102001600173" swrid="4258728" athleteid="46881">
              <RESULTS>
                <RESULT eventid="44380" points="588" reactiontime="+69" swimtime="00:01:01.69" resultid="46882" heatid="50688" lane="1" entrytime="00:01:01.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="574" reactiontime="+68" swimtime="00:00:28.47" resultid="46883" heatid="50835" lane="1" entrytime="00:00:27.93" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Jachym" birthdate="2003-10-30" gender="M" nation="POL" license="102001700089" swrid="4792710" athleteid="46870">
              <RESULTS>
                <RESULT eventid="44378" points="553" reactiontime="+70" swimtime="00:00:57.12" resultid="46871" heatid="50674" lane="6" entrytime="00:00:58.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44390" points="524" reactiontime="+68" swimtime="00:02:21.36" resultid="46872" heatid="50711" lane="6" entrytime="00:02:23.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.13" />
                    <SPLIT distance="100" swimtime="00:01:06.62" />
                    <SPLIT distance="150" swimtime="00:01:48.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="496" reactiontime="+65" swimtime="00:00:28.13" resultid="46873" heatid="50894" lane="1" entrytime="00:00:28.82" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Skowron" birthdate="2006-12-29" gender="M" nation="POL" license="102001700182" swrid="5281325" athleteid="46878">
              <RESULTS>
                <RESULT eventid="44378" points="452" reactiontime="+62" swimtime="00:01:01.10" resultid="46879" heatid="50672" lane="3" entrytime="00:01:01.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="392" reactiontime="+63" swimtime="00:00:30.42" resultid="46880" heatid="50761" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Glejzer" birthdate="2006-02-26" gender="M" nation="POL" license="102001700112" swrid="4995330" athleteid="46866">
              <RESULTS>
                <RESULT eventid="44378" points="509" reactiontime="+47" swimtime="00:00:58.72" resultid="46867" heatid="50674" lane="8" entrytime="00:00:58.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="447" reactiontime="+56" swimtime="00:00:29.11" resultid="46868" heatid="50763" lane="9" entrytime="00:00:35.21" entrycourse="LCM" />
                <RESULT comment="O-1" eventid="46298" status="DSQ" swimtime="00:00:00.00" resultid="46869" heatid="50815" lane="1" entrytime="00:00:30.38" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Franciszek" lastname="Horbacz" birthdate="2007-07-16" gender="M" nation="POL" license="102001700170" swrid="5260099" athleteid="46856">
              <RESULTS>
                <RESULT eventid="44378" points="337" reactiontime="+80" swimtime="00:01:07.37" resultid="46857" heatid="50668" lane="6" entrytime="00:01:06.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="284" reactiontime="+80" swimtime="00:01:18.87" resultid="46858" heatid="50720" lane="2" entrytime="00:01:19.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="307" reactiontime="+78" swimtime="00:02:31.11" resultid="46859" heatid="50734" lane="6" entrytime="00:02:30.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                    <SPLIT distance="100" swimtime="00:01:12.91" />
                    <SPLIT distance="150" swimtime="00:01:53.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="307" reactiontime="+76" swimtime="00:00:33.00" resultid="46860" heatid="50760" lane="2" />
                <RESULT eventid="46298" points="332" reactiontime="+73" swimtime="00:00:30.19" resultid="46861" heatid="50810" lane="5" />
                <RESULT eventid="46310" points="334" reactiontime="+66" swimtime="00:00:34.56" resultid="46862" heatid="50858" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonina" lastname="Horbacz" birthdate="2007-07-16" gender="F" nation="POL" license="102001600171" swrid="5323392" athleteid="46884">
              <RESULTS>
                <RESULT eventid="44380" points="322" reactiontime="+84" swimtime="00:01:15.44" resultid="46885" heatid="50681" lane="7" entrytime="00:01:15.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44396" points="237" reactiontime="+67" swimtime="00:01:33.00" resultid="46886" heatid="50725" lane="9" entrytime="00:01:27.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="253" reactiontime="+81" swimtime="00:00:38.59" resultid="46887" heatid="50770" lane="6" />
                <RESULT eventid="46300" points="381" swimtime="00:00:32.64" resultid="46888" heatid="50824" lane="4" />
                <RESULT eventid="46312" points="258" reactiontime="+69" swimtime="00:00:42.35" resultid="46889" heatid="50904" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Angelika" lastname="Kurowska" birthdate="2007-04-11" gender="F" nation="POL" license="102001600134" swrid="4135401" athleteid="46890">
              <RESULTS>
                <RESULT eventid="44380" points="457" reactiontime="+65" swimtime="00:01:07.13" resultid="46891" heatid="50684" lane="7" entrytime="00:01:07.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44384" status="DNS" swimtime="00:00:00.00" resultid="46892" heatid="50701" lane="8" entrytime="00:00:42.66" entrycourse="LCM" />
                <RESULT eventid="44413" points="334" reactiontime="+68" swimtime="00:00:35.20" resultid="46893" heatid="50774" lane="6" entrytime="00:00:38.51" entrycourse="LCM" />
                <RESULT eventid="46300" status="DNS" swimtime="00:00:00.00" resultid="46894" heatid="50830" lane="8" entrytime="00:00:32.09" entrycourse="LCM" />
                <RESULT eventid="46312" status="DNS" swimtime="00:00:00.00" resultid="46895" heatid="50905" lane="5" entrytime="00:00:42.12" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kornel" lastname="Skowron" birthdate="2005-04-12" gender="M" nation="POL" license="102001700156" swrid="5285295" athleteid="46874">
              <RESULTS>
                <RESULT eventid="44378" points="296" reactiontime="+79" swimtime="00:01:10.36" resultid="46875" heatid="50665" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="270" reactiontime="+59" swimtime="00:01:20.21" resultid="46876" heatid="50718" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="269" swimtime="00:02:53.37" resultid="46877" heatid="50780" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.11" />
                    <SPLIT distance="100" swimtime="00:01:22.53" />
                    <SPLIT distance="150" swimtime="00:02:08.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06601" nation="POL" region="01" clubid="48036" name="UKS ALFA Wałbrzych">
          <ATHLETES>
            <ATHLETE firstname="Michał" lastname="Stelmach" birthdate="2003-02-17" gender="M" nation="POL" license="106601700012" swrid="5088632" athleteid="48050">
              <RESULTS>
                <RESULT eventid="44411" status="DNS" swimtime="00:00:00.00" resultid="48051" heatid="50766" lane="5" entrytime="00:00:29.21" entrycourse="LCM" />
                <RESULT eventid="46298" points="453" reactiontime="+63" swimtime="00:00:27.21" resultid="48052" heatid="50818" lane="7" entrytime="00:00:27.14" entrycourse="LCM" />
                <RESULT eventid="46310" points="441" reactiontime="+85" swimtime="00:00:31.53" resultid="48053" heatid="50860" lane="5" entrytime="00:00:32.46" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alicja" lastname="Maziar" birthdate="2002-07-14" gender="F" nation="POL" license="106601600051" swrid="4792709" athleteid="48041">
              <RESULTS>
                <RESULT eventid="44380" points="470" reactiontime="+65" swimtime="00:01:06.49" resultid="48042" heatid="50686" lane="4" entrytime="00:01:03.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44396" points="429" reactiontime="+73" swimtime="00:01:16.31" resultid="48043" heatid="50728" lane="9" entrytime="00:01:12.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="504" reactiontime="+77" swimtime="00:00:29.73" resultid="48044" heatid="50833" lane="3" entrytime="00:00:29.08" entrycourse="LCM" />
                <RESULT eventid="46312" points="478" reactiontime="+76" swimtime="00:00:34.50" resultid="48045" heatid="50908" lane="3" entrytime="00:00:33.43" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Franczyk" birthdate="2002-09-13" gender="M" nation="POL" license="106601700008" swrid="5166072" athleteid="48037">
              <RESULTS>
                <RESULT eventid="44378" points="433" reactiontime="+63" swimtime="00:01:02.00" resultid="48038" heatid="50672" lane="6" entrytime="00:01:01.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="347" reactiontime="+74" swimtime="00:01:13.74" resultid="48039" heatid="50722" lane="6" entrytime="00:01:10.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="386" reactiontime="+61" swimtime="00:02:20.07" resultid="48040" heatid="50737" lane="9" entrytime="00:02:15.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                    <SPLIT distance="100" swimtime="00:01:07.13" />
                    <SPLIT distance="150" swimtime="00:01:44.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Turków" birthdate="2003-12-03" gender="M" nation="POL" license="106601700002" swrid="5108819" athleteid="48046">
              <RESULTS>
                <RESULT eventid="44382" points="533" reactiontime="+70" swimtime="00:00:32.00" resultid="48047" heatid="50694" lane="4" entrytime="00:00:33.06" entrycourse="LCM" />
                <RESULT eventid="44411" points="476" reactiontime="+69" swimtime="00:00:28.51" resultid="48048" heatid="50759" lane="3" />
                <RESULT eventid="46298" points="468" reactiontime="+70" swimtime="00:00:26.92" resultid="48049" heatid="50819" lane="8" entrytime="00:00:26.59" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00401" nation="POL" region="01" clubid="47098" name="MKS ,,ROKITA&quot; Brzeg Dolny">
          <ATHLETES>
            <ATHLETE firstname="Bartosz" lastname="Geisler" birthdate="2007-03-12" gender="M" nation="POL" license="100401700073" swrid="5219596" athleteid="47099">
              <RESULTS>
                <RESULT eventid="44378" points="233" reactiontime="+45" swimtime="00:01:16.20" resultid="47100" heatid="50665" lane="5" entrytime="00:01:48.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="224" reactiontime="+84" swimtime="00:02:47.75" resultid="47101" heatid="50733" lane="8" entrytime="00:02:48.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.83" />
                    <SPLIT distance="100" swimtime="00:01:18.83" />
                    <SPLIT distance="150" swimtime="00:02:03.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="220" reactiontime="+88" swimtime="00:06:04.49" resultid="47102" heatid="50798" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                    <SPLIT distance="100" swimtime="00:01:19.64" />
                    <SPLIT distance="150" swimtime="00:02:05.36" />
                    <SPLIT distance="200" swimtime="00:02:53.40" />
                    <SPLIT distance="250" swimtime="00:03:41.11" />
                    <SPLIT distance="300" swimtime="00:04:29.58" />
                    <SPLIT distance="350" swimtime="00:05:19.25" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O-1" eventid="46298" reactiontime="+59" status="DSQ" swimtime="00:00:00.00" resultid="47103" heatid="50811" lane="5" entrytime="00:00:49.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Szerszeń" birthdate="2005-11-11" gender="F" nation="POL" license="100401600065" swrid="5213716" athleteid="47130">
              <RESULTS>
                <RESULT eventid="44380" points="306" reactiontime="+91" swimtime="00:01:16.73" resultid="47131" heatid="50682" lane="5" entrytime="00:01:09.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44392" points="284" reactiontime="+90" swimtime="00:03:11.85" resultid="47132" heatid="50713" lane="2" entrytime="00:03:07.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.44" />
                    <SPLIT distance="100" swimtime="00:01:32.40" />
                    <SPLIT distance="150" swimtime="00:02:26.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="282" reactiontime="+89" swimtime="00:02:52.15" resultid="47133" heatid="50740" lane="5" entrytime="00:02:39.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                    <SPLIT distance="100" swimtime="00:01:21.99" />
                    <SPLIT distance="150" swimtime="00:02:09.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="369" reactiontime="+88" swimtime="00:00:33.00" resultid="47134" heatid="50829" lane="3" entrytime="00:00:33.15" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Jurkowski" birthdate="2007-02-15" gender="M" nation="POL" license="100401700077" swrid="5193004" athleteid="47111">
              <RESULTS>
                <RESULT eventid="44378" points="213" reactiontime="+77" swimtime="00:01:18.49" resultid="47112" heatid="50666" lane="8" entrytime="00:01:25.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="376" reactiontime="+80" swimtime="00:00:35.95" resultid="47113" heatid="50690" lane="0" />
                <RESULT eventid="44407" points="371" reactiontime="+75" swimtime="00:01:19.10" resultid="47114" heatid="50748" lane="1" entrytime="00:01:26.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="256" reactiontime="+76" swimtime="00:00:32.92" resultid="47115" heatid="50810" lane="0" />
                <RESULT eventid="46302" points="329" reactiontime="+86" swimtime="00:03:02.57" resultid="47116" heatid="50837" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                    <SPLIT distance="100" swimtime="00:01:26.01" />
                    <SPLIT distance="150" swimtime="00:02:14.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46310" points="201" reactiontime="+85" swimtime="00:00:40.94" resultid="47117" heatid="50857" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Rak" birthdate="2005-07-10" gender="F" nation="POL" license="100401600061" swrid="5088606" athleteid="47124">
              <RESULTS>
                <RESULT eventid="44380" points="472" reactiontime="+75" swimtime="00:01:06.38" resultid="47125" heatid="50685" lane="6" entrytime="00:01:05.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44392" points="436" reactiontime="+76" swimtime="00:02:46.26" resultid="47126" heatid="50714" lane="5" entrytime="00:02:48.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                    <SPLIT distance="100" swimtime="00:01:16.63" />
                    <SPLIT distance="150" swimtime="00:02:08.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="447" reactiontime="+76" swimtime="00:00:31.95" resultid="47127" heatid="50778" lane="1" entrytime="00:00:31.82" entrycourse="LCM" />
                <RESULT eventid="46300" points="489" reactiontime="+71" swimtime="00:00:30.04" resultid="47128" heatid="50833" lane="9" entrytime="00:00:29.60" entrycourse="LCM" />
                <RESULT eventid="46308" points="348" reactiontime="+79" swimtime="00:01:18.86" resultid="47129" heatid="50900" lane="8" entrytime="00:01:16.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Kuźma" birthdate="2005-09-10" gender="F" nation="POL" license="100401600066" swrid="5112213" athleteid="47118">
              <RESULTS>
                <RESULT eventid="44380" status="DNS" swimtime="00:00:00.00" resultid="47119" heatid="50680" lane="4" entrytime="00:01:18.27" entrycourse="LCM" />
                <RESULT eventid="44384" status="DNS" swimtime="00:00:00.00" resultid="47120" heatid="50700" lane="8" entrytime="00:00:45.50" entrycourse="LCM" />
                <RESULT eventid="44409" status="DNS" swimtime="00:00:00.00" resultid="47121" heatid="50753" lane="8" entrytime="00:01:40.87" entrycourse="LCM" />
                <RESULT eventid="46300" status="DNS" swimtime="00:00:00.00" resultid="47122" heatid="50829" lane="9" entrytime="00:00:35.04" entrycourse="LCM" />
                <RESULT eventid="46304" status="DNS" swimtime="00:00:00.00" resultid="47123" heatid="50841" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Jacukiewicz" birthdate="2004-03-21" gender="M" nation="POL" license="100401700074" swrid="4840789" athleteid="47104">
              <RESULTS>
                <RESULT eventid="44378" points="441" reactiontime="+76" swimtime="00:01:01.61" resultid="47105" heatid="50664" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="384" reactiontime="+77" swimtime="00:00:35.68" resultid="47106" heatid="50691" lane="7" />
                <RESULT eventid="44390" points="338" reactiontime="+74" swimtime="00:02:43.64" resultid="47107" heatid="50707" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.78" />
                    <SPLIT distance="100" swimtime="00:01:14.77" />
                    <SPLIT distance="150" swimtime="00:02:01.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="328" reactiontime="+77" swimtime="00:01:22.41" resultid="47108" heatid="50746" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="408" reactiontime="+71" swimtime="00:00:28.19" resultid="47109" heatid="50811" lane="2" />
                <RESULT eventid="46302" points="352" reactiontime="+72" swimtime="00:02:58.57" resultid="47110" heatid="50838" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.04" />
                    <SPLIT distance="100" swimtime="00:01:23.01" />
                    <SPLIT distance="150" swimtime="00:02:10.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00115" nation="POL" region="15" clubid="46954" name="KS Warta Poznań">
          <ATHLETES>
            <ATHLETE firstname="Maja" lastname="Rybak" birthdate="2007-04-23" gender="F" nation="POL" license="100115600454" swrid="5162165" athleteid="46982">
              <RESULTS>
                <RESULT eventid="44384" points="552" reactiontime="+60" swimtime="00:00:35.82" resultid="46983" heatid="50703" lane="9" entrytime="00:00:35.43" entrycourse="LCM" />
                <RESULT eventid="44392" points="539" reactiontime="+61" swimtime="00:02:34.92" resultid="46984" heatid="50714" lane="7" entrytime="00:02:51.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                    <SPLIT distance="100" swimtime="00:01:13.20" />
                    <SPLIT distance="150" swimtime="00:01:58.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44409" points="540" reactiontime="+51" swimtime="00:01:18.72" resultid="46985" heatid="50755" lane="4" entrytime="00:01:18.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46304" points="502" reactiontime="+60" swimtime="00:02:54.93" resultid="46986" heatid="50843" lane="1" entrytime="00:02:50.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.33" />
                    <SPLIT distance="100" swimtime="00:01:22.02" />
                    <SPLIT distance="150" swimtime="00:02:08.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Kolańczyk" birthdate="2006-09-05" gender="F" nation="POL" license="100115600428" swrid="5162144" athleteid="46960">
              <RESULTS>
                <RESULT eventid="44380" points="598" reactiontime="+55" swimtime="00:01:01.36" resultid="46961" heatid="50687" lane="4" entrytime="00:01:01.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="537" reactiontime="+64" swimtime="00:02:18.96" resultid="46962" heatid="50743" lane="3" entrytime="00:02:17.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                    <SPLIT distance="100" swimtime="00:01:08.47" />
                    <SPLIT distance="150" swimtime="00:01:44.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="556" reactiontime="+64" swimtime="00:00:29.70" resultid="46963" heatid="50779" lane="6" entrytime="00:00:29.71" entrycourse="LCM" />
                <RESULT eventid="46300" points="623" reactiontime="+50" swimtime="00:00:27.71" resultid="46964" heatid="50832" lane="4" entrytime="00:00:29.66" entrycourse="LCM" />
                <RESULT eventid="46308" points="520" reactiontime="+69" swimtime="00:01:08.96" resultid="46965" heatid="50901" lane="2" entrytime="00:01:08.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Krasowski" birthdate="2006-10-12" gender="M" nation="POL" license="100115700430" swrid="5162163" athleteid="46977">
              <RESULTS>
                <RESULT eventid="44382" points="483" reactiontime="+67" swimtime="00:00:33.06" resultid="46978" heatid="50694" lane="3" entrytime="00:00:33.19" entrycourse="LCM" />
                <RESULT eventid="44390" points="474" reactiontime="+67" swimtime="00:02:26.20" resultid="46979" heatid="50707" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.05" />
                    <SPLIT distance="100" swimtime="00:01:09.92" />
                    <SPLIT distance="150" swimtime="00:01:50.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="515" reactiontime="+71" swimtime="00:01:10.94" resultid="46980" heatid="50750" lane="2" entrytime="00:01:11.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46306" points="430" reactiontime="+70" swimtime="00:01:05.56" resultid="46981" heatid="50847" lane="7" entrytime="00:01:11.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Celmer" birthdate="2007-03-26" gender="F" nation="POL" license="100115600449" swrid="5162156" athleteid="46996">
              <RESULTS>
                <RESULT eventid="44413" points="569" reactiontime="+66" swimtime="00:00:29.47" resultid="46997" heatid="50779" lane="2" entrytime="00:00:29.72" entrycourse="LCM" />
                <RESULT eventid="46300" points="654" reactiontime="+59" swimtime="00:00:27.26" resultid="46998" heatid="50835" lane="5" entrytime="00:00:26.74" entrycourse="LCM" />
                <RESULT eventid="46312" points="620" reactiontime="+76" swimtime="00:00:31.63" resultid="46999" heatid="50908" lane="4" entrytime="00:00:32.69" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kajetan" lastname="Krucki" birthdate="2006-09-16" gender="M" nation="POL" license="100115700431" swrid="5162145" athleteid="46966">
              <RESULTS>
                <RESULT eventid="44382" points="538" reactiontime="+60" swimtime="00:00:31.90" resultid="46967" heatid="50693" lane="4" entrytime="00:00:36.87" entrycourse="LCM" />
                <RESULT eventid="44411" points="591" reactiontime="+60" swimtime="00:00:26.53" resultid="46968" heatid="50769" lane="9" entrytime="00:00:26.49" entrycourse="LCM" />
                <RESULT eventid="46298" points="590" reactiontime="+62" swimtime="00:00:24.92" resultid="46969" heatid="50821" lane="4" entrytime="00:00:25.03" entrycourse="LCM" />
                <RESULT eventid="46310" points="553" reactiontime="+59" swimtime="00:00:29.23" resultid="46970" heatid="50860" lane="6" entrytime="00:00:33.02" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Chruściel" birthdate="2007-04-23" gender="M" nation="POL" license="100115700450" swrid="5162166" athleteid="46987">
              <RESULTS>
                <RESULT eventid="44394" points="361" reactiontime="+69" swimtime="00:01:12.78" resultid="46988" heatid="50721" lane="3" entrytime="00:01:14.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="352" reactiontime="+70" swimtime="00:00:31.53" resultid="46989" heatid="50764" lane="5" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="46298" points="343" reactiontime="+70" swimtime="00:00:29.85" resultid="46990" heatid="50813" lane="2" entrytime="00:00:33.36" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maksymilian" lastname="Budny" birthdate="2006-05-04" gender="M" nation="POL" license="100115700424" swrid="5162174" athleteid="46971">
              <RESULTS>
                <RESULT eventid="44382" points="495" reactiontime="+65" swimtime="00:00:32.80" resultid="46972" heatid="50692" lane="3" entrytime="00:00:47.32" entrycourse="LCM" />
                <RESULT eventid="44390" points="517" reactiontime="+67" swimtime="00:02:22.02" resultid="46973" heatid="50711" lane="8" entrytime="00:02:25.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.36" />
                    <SPLIT distance="100" swimtime="00:01:08.01" />
                    <SPLIT distance="150" swimtime="00:01:47.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="453" reactiontime="+63" swimtime="00:01:14.03" resultid="46974" heatid="50749" lane="9" entrytime="00:01:21.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="524" reactiontime="+66" swimtime="00:00:25.93" resultid="46975" heatid="50820" lane="1" entrytime="00:00:26.17" entrycourse="LCM" />
                <RESULT eventid="46310" points="517" reactiontime="+69" swimtime="00:00:29.90" resultid="46976" heatid="50861" lane="1" entrytime="00:00:31.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Wrzeszczyńska" birthdate="2007-07-03" gender="F" nation="POL" license="100115600456" swrid="5162152" athleteid="46955">
              <RESULTS>
                <RESULT eventid="44380" points="626" reactiontime="+74" swimtime="00:01:00.42" resultid="46956" heatid="50688" lane="6" entrytime="00:01:00.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="504" reactiontime="+76" swimtime="00:02:21.89" resultid="46957" heatid="50743" lane="6" entrytime="00:02:17.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.38" />
                    <SPLIT distance="100" swimtime="00:01:08.54" />
                    <SPLIT distance="150" swimtime="00:01:45.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="526" reactiontime="+73" swimtime="00:00:30.25" resultid="46958" heatid="50779" lane="0" entrytime="00:00:30.10" entrycourse="LCM" />
                <RESULT eventid="46308" points="576" reactiontime="+74" swimtime="00:01:06.67" resultid="46959" heatid="50901" lane="6" entrytime="00:01:07.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Jarecki" birthdate="2006-10-18" gender="M" nation="POL" license="100115700427" swrid="5162157" athleteid="46991">
              <RESULTS>
                <RESULT eventid="44394" points="396" reactiontime="+74" swimtime="00:01:10.55" resultid="46992" heatid="50722" lane="1" entrytime="00:01:10.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="411" reactiontime="+72" swimtime="00:00:29.95" resultid="46993" heatid="50766" lane="1" entrytime="00:00:29.69" entrycourse="LCM" />
                <RESULT eventid="46298" points="388" reactiontime="+72" swimtime="00:00:28.66" resultid="46994" heatid="50817" lane="1" entrytime="00:00:28.35" entrycourse="LCM" />
                <RESULT eventid="46310" points="396" reactiontime="+70" swimtime="00:00:32.66" resultid="46995" heatid="50860" lane="0" entrytime="00:00:36.59" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="44399" points="494" reactiontime="+76" swimtime="00:04:22.11" resultid="47000" heatid="50729" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.77" />
                    <SPLIT distance="100" swimtime="00:01:11.62" />
                    <SPLIT distance="150" swimtime="00:01:44.67" />
                    <SPLIT distance="200" swimtime="00:02:22.87" />
                    <SPLIT distance="250" swimtime="00:02:50.53" />
                    <SPLIT distance="300" swimtime="00:03:23.44" />
                    <SPLIT distance="350" swimtime="00:03:50.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="46991" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="46977" number="2" reactiontime="+16" />
                    <RELAYPOSITION athleteid="46966" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="46971" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46289" points="493" reactiontime="+64" swimtime="00:03:58.17" resultid="47002" heatid="50793" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.28" />
                    <SPLIT distance="100" swimtime="00:00:56.07" />
                    <SPLIT distance="150" swimtime="00:01:25.22" />
                    <SPLIT distance="200" swimtime="00:01:59.56" />
                    <SPLIT distance="250" swimtime="00:02:27.23" />
                    <SPLIT distance="300" swimtime="00:02:58.43" />
                    <SPLIT distance="350" swimtime="00:03:28.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="46966" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="46991" number="2" />
                    <RELAYPOSITION athleteid="46971" number="3" />
                    <RELAYPOSITION athleteid="46977" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT comment="S-1" eventid="44401" reactiontime="+67" status="DSQ" swimtime="00:04:40.62" resultid="47001" heatid="50887" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                    <SPLIT distance="100" swimtime="00:01:09.33" />
                    <SPLIT distance="150" swimtime="00:01:45.41" />
                    <SPLIT distance="200" swimtime="00:02:28.82" />
                    <SPLIT distance="250" swimtime="00:03:00.19" />
                    <SPLIT distance="300" swimtime="00:03:39.29" />
                    <SPLIT distance="350" swimtime="00:04:08.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="46996" number="1" reactiontime="+67" status="DSQ" />
                    <RELAYPOSITION athleteid="46982" number="2" reactiontime="-20" status="DSQ" />
                    <RELAYPOSITION athleteid="46960" number="3" reactiontime="+44" status="DSQ" />
                    <RELAYPOSITION athleteid="46955" number="4" reactiontime="+1" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46291" points="607" reactiontime="+59" swimtime="00:04:08.01" resultid="47003" heatid="50795" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.14" />
                    <SPLIT distance="100" swimtime="00:01:00.89" />
                    <SPLIT distance="150" swimtime="00:01:30.02" />
                    <SPLIT distance="200" swimtime="00:02:02.57" />
                    <SPLIT distance="250" swimtime="00:02:32.27" />
                    <SPLIT distance="300" swimtime="00:03:06.10" />
                    <SPLIT distance="350" swimtime="00:03:35.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="46996" number="1" reactiontime="+59" />
                    <RELAYPOSITION athleteid="46960" number="2" reactiontime="+30" />
                    <RELAYPOSITION athleteid="46982" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="46955" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02601" nation="POL" region="01" clubid="46896" name="KS WANKAN Legnica">
          <ATHLETES>
            <ATHLETE firstname="Aleksandra" lastname="Lepczak" birthdate="2006-12-08" gender="F" nation="POL" license="102601600133" swrid="5166040" athleteid="46932">
              <RESULTS>
                <RESULT eventid="44380" points="461" reactiontime="+61" swimtime="00:01:06.89" resultid="46933" heatid="50685" lane="9" entrytime="00:01:06.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44396" points="410" reactiontime="+73" swimtime="00:01:17.48" resultid="46934" heatid="50726" lane="4" entrytime="00:01:17.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="388" reactiontime="+67" swimtime="00:02:34.90" resultid="46935" heatid="50741" lane="5" entrytime="00:02:32.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.15" />
                    <SPLIT distance="100" swimtime="00:01:13.77" />
                    <SPLIT distance="150" swimtime="00:01:55.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="380" reactiontime="+73" swimtime="00:00:33.72" resultid="46936" heatid="50772" lane="7" />
                <RESULT eventid="46300" points="492" reactiontime="+66" swimtime="00:00:29.97" resultid="46937" heatid="50832" lane="0" entrytime="00:00:30.02" entrycourse="LCM" />
                <RESULT eventid="46312" points="432" reactiontime="+75" swimtime="00:00:35.69" resultid="46938" heatid="50908" lane="7" entrytime="00:00:34.41" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Sarowski" birthdate="2007-09-10" gender="M" nation="POL" license="102601700105" swrid="5192999" athleteid="46911">
              <RESULTS>
                <RESULT eventid="44378" points="442" reactiontime="+56" swimtime="00:01:01.54" resultid="46912" heatid="50672" lane="4" entrytime="00:01:01.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="362" reactiontime="+67" swimtime="00:01:12.75" resultid="46913" heatid="50722" lane="9" entrytime="00:01:12.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="395" reactiontime="+67" swimtime="00:02:19.01" resultid="46914" heatid="50736" lane="7" entrytime="00:02:17.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                    <SPLIT distance="100" swimtime="00:01:06.94" />
                    <SPLIT distance="150" swimtime="00:01:43.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="364" reactiontime="+70" swimtime="00:00:31.17" resultid="46915" heatid="50765" lane="6" entrytime="00:00:30.31" entrycourse="LCM" />
                <RESULT eventid="46298" points="404" reactiontime="+63" swimtime="00:00:28.27" resultid="46916" heatid="50816" lane="2" entrytime="00:00:29.15" entrycourse="LCM" />
                <RESULT eventid="46306" points="342" reactiontime="+66" swimtime="00:01:10.78" resultid="46917" heatid="50847" lane="6" entrytime="00:01:10.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Borys" lastname="Kaszubowski" birthdate="2008-07-07" gender="M" nation="POL" license="102601700131" swrid="5200953" athleteid="46897">
              <RESULTS>
                <RESULT eventid="44378" points="529" reactiontime="+64" swimtime="00:00:57.99" resultid="46898" heatid="50674" lane="7" entrytime="00:00:58.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="407" reactiontime="+59" swimtime="00:01:09.94" resultid="46899" heatid="50722" lane="8" entrytime="00:01:11.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="457" reactiontime="+65" swimtime="00:02:12.37" resultid="46900" heatid="50737" lane="7" entrytime="00:02:14.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                    <SPLIT distance="100" swimtime="00:01:04.98" />
                    <SPLIT distance="150" swimtime="00:01:40.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="481" reactiontime="+61" swimtime="00:00:28.42" resultid="46901" heatid="50894" lane="5" entrytime="00:00:28.51" entrycourse="LCM" />
                <RESULT eventid="46298" points="467" reactiontime="+55" swimtime="00:00:26.95" resultid="46902" heatid="50817" lane="4" entrytime="00:00:27.79" entrycourse="LCM" />
                <RESULT eventid="46306" points="474" reactiontime="+42" swimtime="00:01:03.48" resultid="46903" heatid="50848" lane="5" entrytime="00:01:03.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kacper" lastname="Kubiak" birthdate="2008-04-15" gender="M" nation="POL" license="102601700129" swrid="5334381" athleteid="46918">
              <RESULTS>
                <RESULT eventid="44378" points="291" reactiontime="+54" swimtime="00:01:10.72" resultid="46919" heatid="50667" lane="1" entrytime="00:01:10.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="256" reactiontime="+61" swimtime="00:01:21.61" resultid="46920" heatid="50719" lane="7" entrytime="00:01:24.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="261" reactiontime="+52" swimtime="00:02:39.44" resultid="46921" heatid="50733" lane="6" entrytime="00:02:40.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                    <SPLIT distance="100" swimtime="00:01:15.97" />
                    <SPLIT distance="150" swimtime="00:01:59.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="234" reactiontime="+54" swimtime="00:00:36.12" resultid="46922" heatid="50762" lane="3" entrytime="00:00:36.74" entrycourse="LCM" />
                <RESULT eventid="46298" points="272" swimtime="00:00:32.27" resultid="46923" heatid="50808" lane="4" />
                <RESULT eventid="46310" points="270" swimtime="00:00:37.11" resultid="46924" heatid="50860" lane="9" entrytime="00:00:37.04" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Szymkowicz" birthdate="2007-03-23" gender="M" nation="POL" license="102601700107" swrid="5081122" athleteid="46904">
              <RESULTS>
                <RESULT eventid="44378" points="388" reactiontime="+79" swimtime="00:01:04.27" resultid="46905" heatid="50670" lane="7" entrytime="00:01:04.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="391" reactiontime="+68" swimtime="00:01:10.89" resultid="46906" heatid="50722" lane="0" entrytime="00:01:11.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="380" reactiontime="+65" swimtime="00:02:20.81" resultid="46907" heatid="50735" lane="5" entrytime="00:02:23.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.81" />
                    <SPLIT distance="100" swimtime="00:01:08.25" />
                    <SPLIT distance="150" swimtime="00:01:45.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="379" reactiontime="+81" swimtime="00:00:30.75" resultid="46908" heatid="50765" lane="3" entrytime="00:00:30.28" entrycourse="LCM" />
                <RESULT eventid="46298" points="361" reactiontime="+75" swimtime="00:00:29.36" resultid="46909" heatid="50816" lane="9" entrytime="00:00:29.62" entrycourse="LCM" />
                <RESULT eventid="46310" points="423" reactiontime="+93" swimtime="00:00:31.97" resultid="46910" heatid="50861" lane="2" entrytime="00:00:31.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Kulas" birthdate="2007-05-12" gender="F" nation="POL" license="102601600104" swrid="5072846" athleteid="46946">
              <RESULTS>
                <RESULT eventid="44380" points="390" reactiontime="+56" swimtime="00:01:10.74" resultid="46947" heatid="50684" lane="5" entrytime="00:01:06.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44396" points="360" reactiontime="+78" swimtime="00:01:20.91" resultid="46948" heatid="50726" lane="2" entrytime="00:01:18.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="375" reactiontime="+65" swimtime="00:02:36.64" resultid="46949" heatid="50741" lane="3" entrytime="00:02:33.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.48" />
                    <SPLIT distance="100" swimtime="00:01:15.44" />
                    <SPLIT distance="150" swimtime="00:01:57.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="335" reactiontime="+66" swimtime="00:00:35.15" resultid="46950" heatid="50777" lane="2" entrytime="00:00:32.98" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliwia" lastname="Wiesiołek" birthdate="2005-01-05" gender="F" nation="POL" license="102601600091" swrid="5200942" athleteid="46925">
              <RESULTS>
                <RESULT eventid="44380" points="560" reactiontime="+65" swimtime="00:01:02.73" resultid="46926" heatid="50687" lane="7" entrytime="00:01:02.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44396" points="482" reactiontime="+63" swimtime="00:01:13.38" resultid="46927" heatid="50728" lane="8" entrytime="00:01:11.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="474" reactiontime="+67" swimtime="00:02:24.87" resultid="46928" heatid="50742" lane="2" entrytime="00:02:26.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.97" />
                    <SPLIT distance="100" swimtime="00:01:10.04" />
                    <SPLIT distance="150" swimtime="00:01:47.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="422" reactiontime="+66" swimtime="00:00:32.55" resultid="46929" heatid="50777" lane="0" entrytime="00:00:33.48" entrycourse="LCM" />
                <RESULT eventid="46300" points="566" reactiontime="+65" swimtime="00:00:28.61" resultid="46930" heatid="50834" lane="7" entrytime="00:00:28.59" entrycourse="LCM" />
                <RESULT eventid="46312" points="566" reactiontime="+61" swimtime="00:00:32.61" resultid="46931" heatid="50909" lane="9" entrytime="00:00:32.35" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="44399" points="362" reactiontime="+75" swimtime="00:04:50.84" resultid="46951" heatid="50729" lane="4" entrytime="00:04:59.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.15" />
                    <SPLIT distance="100" swimtime="00:01:09.89" />
                    <SPLIT distance="150" swimtime="00:01:50.05" />
                    <SPLIT distance="200" swimtime="00:02:35.84" />
                    <SPLIT distance="250" swimtime="00:03:05.68" />
                    <SPLIT distance="300" swimtime="00:03:40.20" />
                    <SPLIT distance="350" swimtime="00:04:13.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="46904" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="46911" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="46897" number="3" />
                    <RELAYPOSITION athleteid="46918" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46289" points="372" swimtime="00:04:21.56" resultid="46952" heatid="50793" lane="5" entrytime="00:04:13.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                    <SPLIT distance="100" swimtime="00:01:12.58" />
                    <SPLIT distance="150" swimtime="00:01:43.11" />
                    <SPLIT distance="200" swimtime="00:02:17.22" />
                    <SPLIT distance="250" swimtime="00:02:47.95" />
                    <SPLIT distance="300" swimtime="00:03:22.26" />
                    <SPLIT distance="350" swimtime="00:03:51.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="46918" number="1" />
                    <RELAYPOSITION athleteid="46904" number="2" />
                    <RELAYPOSITION athleteid="46911" number="3" />
                    <RELAYPOSITION athleteid="46897" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46314" points="381" reactiontime="+73" swimtime="00:09:37.31" resultid="46953" heatid="50870" lane="3" entrytime="00:09:34.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.10" />
                    <SPLIT distance="100" swimtime="00:01:07.12" />
                    <SPLIT distance="150" swimtime="00:01:45.03" />
                    <SPLIT distance="200" swimtime="00:02:22.72" />
                    <SPLIT distance="250" swimtime="00:02:56.83" />
                    <SPLIT distance="300" swimtime="00:03:36.59" />
                    <SPLIT distance="350" swimtime="00:04:19.00" />
                    <SPLIT distance="400" swimtime="00:05:00.99" />
                    <SPLIT distance="450" swimtime="00:05:32.41" />
                    <SPLIT distance="500" swimtime="00:06:07.97" />
                    <SPLIT distance="550" swimtime="00:06:44.94" />
                    <SPLIT distance="600" swimtime="00:07:21.67" />
                    <SPLIT distance="650" swimtime="00:07:51.81" />
                    <SPLIT distance="700" swimtime="00:08:26.71" />
                    <SPLIT distance="750" swimtime="00:09:02.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="46904" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="46918" number="2" reactiontime="+38" />
                    <RELAYPOSITION athleteid="46911" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="46897" number="4" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="08314" nation="POL" region="14" clubid="48098" name="UKS Delfin Garwolin">
          <ATHLETES>
            <ATHLETE firstname="Jakub" lastname="Sitnik" birthdate="2003-10-07" gender="M" nation="POL" license="108314700020" swrid="5120231" athleteid="48099">
              <RESULTS>
                <RESULT eventid="44378" points="500" reactiontime="+73" swimtime="00:00:59.08" resultid="48100" heatid="50673" lane="2" entrytime="00:00:59.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="528" swimtime="00:00:27.55" resultid="48101" heatid="50767" lane="9" entrytime="00:00:29.17" entrycourse="LCM" />
                <RESULT eventid="46298" points="516" reactiontime="+69" swimtime="00:00:26.06" resultid="48102" heatid="50821" lane="1" entrytime="00:00:25.73" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00304" nation="POL" region="04" clubid="47652" name="TP Zielona Góra">
          <ATHLETES>
            <ATHLETE firstname="Kajetan" lastname="Sobiechowski" birthdate="2006-12-25" gender="M" nation="POL" license="100304700483" swrid="5186690" athleteid="47653">
              <RESULTS>
                <RESULT eventid="44378" points="560" reactiontime="+64" swimtime="00:00:56.90" resultid="47654" heatid="50669" lane="4" entrytime="00:01:05.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="519" reactiontime="+72" swimtime="00:02:06.89" resultid="47655" heatid="50738" lane="2" entrytime="00:02:06.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.07" />
                    <SPLIT distance="100" swimtime="00:00:59.95" />
                    <SPLIT distance="150" swimtime="00:01:33.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="532" swimtime="00:00:27.47" resultid="47656" heatid="50767" lane="8" entrytime="00:00:28.85" entrycourse="LCM" />
                <RESULT eventid="46294" points="555" reactiontime="+71" swimtime="00:04:27.76" resultid="47657" heatid="50800" lane="7" entrytime="00:04:34.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.35" />
                    <SPLIT distance="100" swimtime="00:01:02.45" />
                    <SPLIT distance="150" swimtime="00:01:36.79" />
                    <SPLIT distance="200" swimtime="00:02:11.92" />
                    <SPLIT distance="250" swimtime="00:02:47.43" />
                    <SPLIT distance="300" swimtime="00:03:22.23" />
                    <SPLIT distance="350" swimtime="00:03:57.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="532" reactiontime="+64" swimtime="00:00:25.80" resultid="47658" heatid="50820" lane="9" entrytime="00:00:26.25" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01910" nation="POL" region="10" clubid="46584" name="KS Delfin Gdynia">
          <ATHLETES>
            <ATHLETE firstname="Adam" lastname="Zdybel" birthdate="2005-03-12" gender="M" nation="POL" license="101910700109" swrid="5030779" athleteid="46585">
              <RESULTS>
                <RESULT eventid="44378" points="696" reactiontime="+62" swimtime="00:00:52.93" resultid="46586" heatid="50677" lane="7" entrytime="00:00:52.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44386" points="623" reactiontime="+65" swimtime="00:02:09.60" resultid="46587" heatid="50705" lane="6" entrytime="00:02:18.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.74" />
                    <SPLIT distance="100" swimtime="00:01:01.62" />
                    <SPLIT distance="150" swimtime="00:01:35.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="698" reactiontime="+62" swimtime="00:01:54.94" resultid="46588" heatid="50739" lane="4" entrytime="00:01:53.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.09" />
                    <SPLIT distance="100" swimtime="00:00:56.54" />
                    <SPLIT distance="150" swimtime="00:01:26.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="575" reactiontime="+63" swimtime="00:00:26.78" resultid="46589" heatid="50758" lane="8" />
                <RESULT eventid="46285" points="629" reactiontime="+63" swimtime="00:16:56.11" resultid="46590" heatid="50789" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.70" />
                    <SPLIT distance="100" swimtime="00:01:02.67" />
                    <SPLIT distance="150" swimtime="00:01:36.08" />
                    <SPLIT distance="200" swimtime="00:02:09.49" />
                    <SPLIT distance="250" swimtime="00:02:43.14" />
                    <SPLIT distance="300" swimtime="00:03:16.90" />
                    <SPLIT distance="350" swimtime="00:03:50.51" />
                    <SPLIT distance="400" swimtime="00:04:24.61" />
                    <SPLIT distance="450" swimtime="00:04:58.75" />
                    <SPLIT distance="500" swimtime="00:05:33.15" />
                    <SPLIT distance="550" swimtime="00:06:06.98" />
                    <SPLIT distance="600" swimtime="00:06:41.16" />
                    <SPLIT distance="650" swimtime="00:07:15.36" />
                    <SPLIT distance="700" swimtime="00:07:49.92" />
                    <SPLIT distance="750" swimtime="00:08:23.99" />
                    <SPLIT distance="800" swimtime="00:08:58.93" />
                    <SPLIT distance="850" swimtime="00:09:32.85" />
                    <SPLIT distance="900" swimtime="00:10:07.45" />
                    <SPLIT distance="950" swimtime="00:10:41.38" />
                    <SPLIT distance="1000" swimtime="00:11:16.04" />
                    <SPLIT distance="1050" swimtime="00:11:50.01" />
                    <SPLIT distance="1100" swimtime="00:12:24.23" />
                    <SPLIT distance="1150" swimtime="00:12:58.36" />
                    <SPLIT distance="1200" swimtime="00:13:33.25" />
                    <SPLIT distance="1250" swimtime="00:14:07.64" />
                    <SPLIT distance="1300" swimtime="00:14:42.21" />
                    <SPLIT distance="1350" swimtime="00:15:16.62" />
                    <SPLIT distance="1400" swimtime="00:15:51.14" />
                    <SPLIT distance="1450" swimtime="00:16:24.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="730" reactiontime="+63" swimtime="00:04:04.40" resultid="46591" heatid="50800" lane="4" entrytime="00:04:05.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.67" />
                    <SPLIT distance="100" swimtime="00:00:57.96" />
                    <SPLIT distance="150" swimtime="00:01:29.12" />
                    <SPLIT distance="200" swimtime="00:02:00.30" />
                    <SPLIT distance="250" swimtime="00:02:31.55" />
                    <SPLIT distance="300" swimtime="00:03:03.12" />
                    <SPLIT distance="350" swimtime="00:03:34.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="605" reactiontime="+61" swimtime="00:00:24.72" resultid="46592" heatid="50822" lane="8" entrytime="00:00:24.67" entrycourse="LCM" />
                <RESULT eventid="46306" points="597" reactiontime="+61" swimtime="00:00:58.78" resultid="46593" heatid="50849" lane="3" entrytime="00:00:58.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03601" nation="POL" region="01" clubid="47668" name="UKP ,,TORPEDA&apos;&apos; Oleśnica">
          <ATHLETES>
            <ATHLETE firstname="Alicja" lastname="Szwabińśka" birthdate="2006-04-18" gender="F" nation="POL" license="103601600023" swrid="5043018" athleteid="47676">
              <RESULTS>
                <RESULT eventid="44380" points="555" reactiontime="+75" swimtime="00:01:02.90" resultid="47677" heatid="50685" lane="5" entrytime="00:01:05.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="418" reactiontime="+75" swimtime="00:00:32.66" resultid="47678" heatid="50771" lane="1" />
                <RESULT eventid="46296" points="540" reactiontime="+75" swimtime="00:04:50.26" resultid="47679" heatid="50804" lane="3" entrytime="00:05:01.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                    <SPLIT distance="100" swimtime="00:01:09.21" />
                    <SPLIT distance="150" swimtime="00:01:46.81" />
                    <SPLIT distance="200" swimtime="00:02:24.13" />
                    <SPLIT distance="250" swimtime="00:03:01.63" />
                    <SPLIT distance="300" swimtime="00:03:38.65" />
                    <SPLIT distance="350" swimtime="00:04:15.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="521" reactiontime="+74" swimtime="00:00:29.40" resultid="47680" heatid="50833" lane="7" entrytime="00:00:29.12" entrycourse="LCM" />
                <RESULT eventid="46312" points="490" reactiontime="+74" swimtime="00:00:34.22" resultid="47681" heatid="50907" lane="1" entrytime="00:00:36.67" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrianna" lastname="Szwabińska" birthdate="2003-07-14" gender="F" nation="POL" license="103601600018" swrid="4931148" athleteid="47669">
              <RESULTS>
                <RESULT eventid="44380" points="697" reactiontime="+67" swimtime="00:00:58.30" resultid="47670" heatid="50688" lane="4" entrytime="00:00:57.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44384" points="624" reactiontime="+68" swimtime="00:00:34.39" resultid="47671" heatid="50703" lane="7" entrytime="00:00:34.65" entrycourse="LCM" />
                <RESULT eventid="44405" points="664" reactiontime="+62" swimtime="00:02:09.47" resultid="47672" heatid="50744" lane="4" entrytime="00:02:08.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.67" />
                    <SPLIT distance="100" swimtime="00:01:03.76" />
                    <SPLIT distance="150" swimtime="00:01:37.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="540" reactiontime="+64" swimtime="00:00:30.00" resultid="47673" heatid="50779" lane="9" entrytime="00:00:30.48" entrycourse="LCM" />
                <RESULT eventid="46296" points="562" reactiontime="+71" swimtime="00:04:46.44" resultid="47674" heatid="50805" lane="1" entrytime="00:04:45.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                    <SPLIT distance="100" swimtime="00:01:06.77" />
                    <SPLIT distance="150" swimtime="00:01:42.51" />
                    <SPLIT distance="200" swimtime="00:02:18.83" />
                    <SPLIT distance="250" swimtime="00:02:55.56" />
                    <SPLIT distance="300" swimtime="00:03:33.00" />
                    <SPLIT distance="350" swimtime="00:04:10.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="694" reactiontime="+65" swimtime="00:00:26.73" resultid="47675" heatid="50835" lane="4" entrytime="00:00:26.24" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Okoń" birthdate="2007-07-10" gender="M" nation="POL" license="103601700022" swrid="5147685" athleteid="47687">
              <RESULTS>
                <RESULT eventid="44394" points="477" reactiontime="+68" swimtime="00:01:06.36" resultid="47688" heatid="50723" lane="8" entrytime="00:01:05.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="469" reactiontime="+68" swimtime="00:00:28.66" resultid="47689" heatid="50758" lane="1" />
                <RESULT eventid="44415" points="462" reactiontime="+71" swimtime="00:02:24.71" resultid="47690" heatid="50784" lane="1" entrytime="00:02:22.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                    <SPLIT distance="100" swimtime="00:01:12.66" />
                    <SPLIT distance="150" swimtime="00:01:50.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="506" reactiontime="+64" swimtime="00:00:26.24" resultid="47691" heatid="50807" lane="5" />
                <RESULT eventid="46310" points="509" reactiontime="+63" swimtime="00:00:30.04" resultid="47692" heatid="50861" lane="4" entrytime="00:00:30.71" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Okoń" birthdate="2007-07-10" gender="M" nation="POL" license="103601700021" swrid="5147682" athleteid="47682">
              <RESULTS>
                <RESULT eventid="44382" points="430" reactiontime="+68" swimtime="00:00:34.37" resultid="47683" heatid="50691" lane="3" />
                <RESULT eventid="44407" points="402" reactiontime="+73" swimtime="00:01:17.04" resultid="47684" heatid="50746" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="430" reactiontime="+71" swimtime="00:00:27.69" resultid="47685" heatid="50808" lane="7" />
                <RESULT eventid="46302" points="403" reactiontime="+75" swimtime="00:02:50.62" resultid="47686" heatid="50837" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.24" />
                    <SPLIT distance="100" swimtime="00:01:22.68" />
                    <SPLIT distance="150" swimtime="00:02:07.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01001" nation="POL" region="01" clubid="48203" name="UKS KORAL Wrocław">
          <ATHLETES>
            <ATHLETE firstname="Alicja" lastname="Orman" birthdate="2007-11-09" gender="F" nation="POL" license="101001600288" swrid="5220819" athleteid="48358">
              <RESULTS>
                <RESULT eventid="44384" points="336" reactiontime="+94" swimtime="00:00:42.25" resultid="48359" heatid="50700" lane="0" entrytime="00:00:46.10" entrycourse="LCM" />
                <RESULT eventid="44396" points="210" reactiontime="+94" swimtime="00:01:36.76" resultid="48360" heatid="50724" lane="5" entrytime="00:01:35.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44409" points="330" reactiontime="+89" swimtime="00:01:32.71" resultid="48361" heatid="50754" lane="0" entrytime="00:01:31.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46304" points="333" reactiontime="+87" swimtime="00:03:20.56" resultid="48362" heatid="50842" lane="7" entrytime="00:03:46.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.44" />
                    <SPLIT distance="100" swimtime="00:01:34.34" />
                    <SPLIT distance="150" swimtime="00:02:27.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="238" reactiontime="+87" swimtime="00:00:43.52" resultid="48363" heatid="50902" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Jastrzębski" birthdate="2007-04-19" gender="M" nation="POL" license="101001700284" swrid="5272051" athleteid="48234">
              <RESULTS>
                <RESULT eventid="44378" points="359" reactiontime="+95" swimtime="00:01:05.99" resultid="48235" heatid="50669" lane="8" entrytime="00:01:05.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="316" reactiontime="+86" swimtime="00:02:29.66" resultid="48236" heatid="50735" lane="7" entrytime="00:02:25.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                    <SPLIT distance="100" swimtime="00:01:12.77" />
                    <SPLIT distance="150" swimtime="00:01:53.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" status="DNS" swimtime="00:00:00.00" resultid="48237" heatid="50757" lane="5" />
                <RESULT eventid="46298" points="355" reactiontime="+86" swimtime="00:00:29.53" resultid="48238" heatid="50809" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nina" lastname="Duszyńska" birthdate="2007-05-28" gender="F" nation="POL" license="101001600281" swrid="5272097" athleteid="48314">
              <RESULTS>
                <RESULT eventid="44380" points="398" reactiontime="+68" swimtime="00:01:10.27" resultid="48315" heatid="50682" lane="1" entrytime="00:01:10.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44396" points="348" reactiontime="+76" swimtime="00:01:21.80" resultid="48316" heatid="50725" lane="1" entrytime="00:01:26.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="282" reactiontime="+58" swimtime="00:00:37.25" resultid="48317" heatid="50773" lane="9" />
                <RESULT eventid="46300" points="424" reactiontime="+72" swimtime="00:00:31.50" resultid="48318" heatid="50824" lane="6" />
                <RESULT eventid="46312" points="350" reactiontime="+74" swimtime="00:00:38.28" resultid="48319" heatid="50904" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martyna" lastname="Łata" birthdate="2007-08-04" gender="F" nation="POL" license="101001600287" swrid="5272093" athleteid="48287">
              <RESULTS>
                <RESULT eventid="44380" points="297" reactiontime="+91" swimtime="00:01:17.50" resultid="48288" heatid="50680" lane="6" entrytime="00:01:18.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="285" reactiontime="+78" swimtime="00:02:51.59" resultid="48289" heatid="50740" lane="8" entrytime="00:02:54.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.48" />
                    <SPLIT distance="100" swimtime="00:01:20.57" />
                    <SPLIT distance="150" swimtime="00:02:08.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="269" reactiontime="+76" swimtime="00:06:06.06" resultid="48290" heatid="50803" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.64" />
                    <SPLIT distance="100" swimtime="00:01:23.38" />
                    <SPLIT distance="150" swimtime="00:02:09.92" />
                    <SPLIT distance="200" swimtime="00:02:57.41" />
                    <SPLIT distance="250" swimtime="00:03:45.54" />
                    <SPLIT distance="300" swimtime="00:04:33.43" />
                    <SPLIT distance="350" swimtime="00:05:21.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="314" reactiontime="+71" swimtime="00:00:34.79" resultid="48291" heatid="50824" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hanna" lastname="Tamoń" birthdate="2007-08-26" gender="F" nation="POL" license="101001600246" swrid="5222173" athleteid="48274">
              <RESULTS>
                <RESULT eventid="44380" points="282" reactiontime="+69" swimtime="00:01:18.77" resultid="48275" heatid="50681" lane="1" entrytime="00:01:16.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44396" points="309" reactiontime="+68" swimtime="00:01:25.07" resultid="48276" heatid="50724" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="258" reactiontime="+65" swimtime="00:00:38.34" resultid="48277" heatid="50770" lane="2" />
                <RESULT eventid="46312" points="325" reactiontime="+80" swimtime="00:00:39.23" resultid="48278" heatid="50904" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Szczepaniak" birthdate="2006-06-10" gender="F" nation="POL" license="101001600236" swrid="5222197" athleteid="48279">
              <RESULTS>
                <RESULT eventid="44380" points="455" reactiontime="+77" swimtime="00:01:07.21" resultid="48280" heatid="50685" lane="8" entrytime="00:01:05.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="467" reactiontime="+77" swimtime="00:02:25.61" resultid="48281" heatid="50742" lane="5" entrytime="00:02:23.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                    <SPLIT distance="100" swimtime="00:01:11.30" />
                    <SPLIT distance="150" swimtime="00:01:49.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46296" points="406" reactiontime="+79" swimtime="00:05:19.28" resultid="48282" heatid="50802" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                    <SPLIT distance="100" swimtime="00:01:15.54" />
                    <SPLIT distance="150" swimtime="00:01:57.32" />
                    <SPLIT distance="200" swimtime="00:02:39.11" />
                    <SPLIT distance="250" swimtime="00:03:20.84" />
                    <SPLIT distance="300" swimtime="00:04:01.51" />
                    <SPLIT distance="350" swimtime="00:04:41.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roksana" lastname="Zima" birthdate="2007-01-23" gender="F" nation="POL" license="101001600302" swrid="5272083" athleteid="48353">
              <RESULTS>
                <RESULT eventid="44384" points="395" reactiontime="+70" swimtime="00:00:40.04" resultid="48354" heatid="50699" lane="8" />
                <RESULT eventid="44409" points="334" reactiontime="+74" swimtime="00:01:32.38" resultid="48355" heatid="50754" lane="2" entrytime="00:01:25.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="222" reactiontime="+76" swimtime="00:00:40.30" resultid="48356" heatid="50771" lane="7" />
                <RESULT eventid="46304" points="326" reactiontime="+75" swimtime="00:03:22.03" resultid="48357" heatid="50841" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.62" />
                    <SPLIT distance="100" swimtime="00:01:33.61" />
                    <SPLIT distance="150" swimtime="00:02:27.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natan" lastname="Kuc" birthdate="2007-03-11" gender="M" nation="POL" license="101001700285" swrid="5272055" athleteid="48334">
              <RESULTS>
                <RESULT eventid="44382" points="263" reactiontime="+82" swimtime="00:00:40.47" resultid="48335" heatid="50690" lane="2" />
                <RESULT eventid="44390" points="304" reactiontime="+92" swimtime="00:02:49.41" resultid="48336" heatid="50709" lane="1" entrytime="00:02:49.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                    <SPLIT distance="100" swimtime="00:01:22.62" />
                    <SPLIT distance="150" swimtime="00:02:11.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="246" reactiontime="+86" swimtime="00:01:30.77" resultid="48337" heatid="50747" lane="2" entrytime="00:01:33.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="240" swimtime="00:00:35.81" resultid="48338" heatid="50757" lane="4" />
                <RESULT eventid="46306" points="221" reactiontime="+82" swimtime="00:01:21.79" resultid="48339" heatid="50844" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natasza" lastname="Roziel" birthdate="2008-08-07" gender="F" nation="POL" license="101001600271" swrid="5318123" athleteid="48327">
              <RESULTS>
                <RESULT eventid="44380" points="427" swimtime="00:01:08.64" resultid="48328" heatid="50682" lane="4" entrytime="00:01:09.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44388" points="316" reactiontime="+92" swimtime="00:02:58.82" resultid="48329" heatid="50706" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.35" />
                    <SPLIT distance="100" swimtime="00:01:23.87" />
                    <SPLIT distance="150" swimtime="00:02:11.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44405" points="422" reactiontime="+84" swimtime="00:02:30.53" resultid="48330" heatid="50741" lane="0" entrytime="00:02:36.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                    <SPLIT distance="100" swimtime="00:01:12.37" />
                    <SPLIT distance="150" swimtime="00:01:52.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="341" reactiontime="+83" swimtime="00:00:34.95" resultid="48331" heatid="50775" lane="2" entrytime="00:00:35.98" entrycourse="LCM" />
                <RESULT eventid="46296" points="424" swimtime="00:05:14.67" resultid="48332" heatid="50803" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                    <SPLIT distance="100" swimtime="00:01:14.13" />
                    <SPLIT distance="150" swimtime="00:01:54.17" />
                    <SPLIT distance="200" swimtime="00:02:35.00" />
                    <SPLIT distance="250" swimtime="00:03:16.03" />
                    <SPLIT distance="300" swimtime="00:03:57.27" />
                    <SPLIT distance="350" swimtime="00:04:37.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46308" points="346" reactiontime="+80" swimtime="00:01:18.99" resultid="48333" heatid="50899" lane="0" entrytime="00:01:21.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olimpia" lastname="Sałapata" birthdate="2007-09-11" gender="F" nation="POL" license="101001600293" swrid="5272060" athleteid="48298">
              <RESULTS>
                <RESULT eventid="44380" points="275" reactiontime="+90" swimtime="00:01:19.47" resultid="48299" heatid="50680" lane="3" entrytime="00:01:18.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44384" points="203" reactiontime="+89" swimtime="00:00:49.97" resultid="48300" heatid="50699" lane="1" />
                <RESULT eventid="44413" points="281" reactiontime="+87" swimtime="00:00:37.28" resultid="48301" heatid="50771" lane="6" />
                <RESULT eventid="46300" points="303" reactiontime="+86" swimtime="00:00:35.24" resultid="48302" heatid="50826" lane="3" />
                <RESULT eventid="46308" points="178" swimtime="00:01:38.49" resultid="48303" heatid="50897" lane="4" entrytime="00:01:53.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Nowak" birthdate="2008-10-29" gender="M" nation="POL" license="101001700265" swrid="5341332" athleteid="48262">
              <RESULTS>
                <RESULT eventid="44378" points="275" swimtime="00:01:12.10" resultid="48263" heatid="50667" lane="8" entrytime="00:01:12.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44390" points="261" reactiontime="+78" swimtime="00:02:58.29" resultid="48264" heatid="50709" lane="9" entrytime="00:02:57.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.24" />
                    <SPLIT distance="100" swimtime="00:01:25.00" />
                    <SPLIT distance="150" swimtime="00:02:19.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="259" reactiontime="+77" swimtime="00:00:34.90" resultid="48265" heatid="50762" lane="5" entrytime="00:00:36.56" entrycourse="LCM" />
                <RESULT eventid="46298" points="274" reactiontime="+79" swimtime="00:00:32.17" resultid="48266" heatid="50813" lane="1" entrytime="00:00:33.53" entrycourse="LCM" />
                <RESULT eventid="46306" points="220" reactiontime="+79" swimtime="00:01:21.99" resultid="48267" heatid="50844" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zofia" lastname="Grządziel" birthdate="2008-04-01" gender="F" nation="POL" license="101001600282" swrid="5272085" athleteid="48364">
              <RESULTS>
                <RESULT eventid="44392" points="359" reactiontime="+66" swimtime="00:02:57.44" resultid="48365" heatid="50713" lane="5" entrytime="00:02:58.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                    <SPLIT distance="100" swimtime="00:01:24.78" />
                    <SPLIT distance="150" swimtime="00:02:15.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44409" points="343" reactiontime="+65" swimtime="00:01:31.57" resultid="48366" heatid="50754" lane="9" entrytime="00:01:33.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="295" reactiontime="+75" swimtime="00:00:36.66" resultid="48367" heatid="50774" lane="3" entrytime="00:00:38.51" entrycourse="LCM" />
                <RESULT eventid="46304" points="350" reactiontime="+81" swimtime="00:03:17.32" resultid="48368" heatid="50841" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.82" />
                    <SPLIT distance="100" swimtime="00:01:33.77" />
                    <SPLIT distance="150" swimtime="00:02:25.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46308" points="287" reactiontime="+66" swimtime="00:01:24.09" resultid="48369" heatid="50898" lane="2" entrytime="00:01:26.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Białek" birthdate="2007-06-19" gender="F" nation="POL" license="101001600279" swrid="5272061" athleteid="48304">
              <RESULTS>
                <RESULT eventid="44380" points="189" reactiontime="+79" swimtime="00:01:30.10" resultid="48305" heatid="50679" lane="4" entrytime="00:01:32.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44384" points="212" reactiontime="+98" swimtime="00:00:49.28" resultid="48306" heatid="50698" lane="2" />
                <RESULT eventid="44409" points="200" reactiontime="+98" swimtime="00:01:49.51" resultid="48307" heatid="50752" lane="6" entrytime="00:01:54.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="205" reactiontime="+87" swimtime="00:00:40.09" resultid="48308" heatid="50828" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Pniaczek" birthdate="2006-01-10" gender="F" nation="POL" license="101001600232" swrid="5222178" athleteid="48283">
              <RESULTS>
                <RESULT eventid="44380" points="411" reactiontime="+71" swimtime="00:01:09.51" resultid="48284" heatid="50684" lane="0" entrytime="00:01:07.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="343" reactiontime="+68" swimtime="00:00:34.87" resultid="48285" heatid="50771" lane="9" />
                <RESULT eventid="46300" points="441" reactiontime="+73" swimtime="00:00:31.08" resultid="48286" heatid="50824" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartek" lastname="Szczepaniak" birthdate="2007-10-19" gender="M" nation="POL" license="101001700295" swrid="5272050" athleteid="48370">
              <RESULTS>
                <RESULT eventid="44394" points="336" reactiontime="+59" swimtime="00:01:14.57" resultid="48371" heatid="50721" lane="9" entrytime="00:01:15.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="309" reactiontime="+64" swimtime="00:02:45.47" resultid="48372" heatid="50782" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.59" />
                    <SPLIT distance="100" swimtime="00:01:19.78" />
                    <SPLIT distance="150" swimtime="00:02:04.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="307" reactiontime="+84" swimtime="00:00:30.99" resultid="48373" heatid="50809" lane="3" />
                <RESULT eventid="46310" points="359" reactiontime="+61" swimtime="00:00:33.76" resultid="48374" heatid="50858" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mikołaj" lastname="Pukas" birthdate="2006-01-06" gender="M" nation="POL" license="101001700233" swrid="5222183" athleteid="48217">
              <RESULTS>
                <RESULT eventid="44378" points="411" reactiontime="+65" swimtime="00:01:03.07" resultid="48218" heatid="50671" lane="5" entrytime="00:01:02.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44390" points="360" reactiontime="+69" swimtime="00:02:40.18" resultid="48219" heatid="50710" lane="0" entrytime="00:02:36.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.91" />
                    <SPLIT distance="100" swimtime="00:01:13.43" />
                    <SPLIT distance="150" swimtime="00:02:04.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="418" reactiontime="+60" swimtime="00:01:09.30" resultid="48220" heatid="50722" lane="7" entrytime="00:01:10.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="412" reactiontime="+60" swimtime="00:02:30.31" resultid="48221" heatid="50782" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.06" />
                    <SPLIT distance="100" swimtime="00:01:14.34" />
                    <SPLIT distance="150" swimtime="00:01:53.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46285" points="348" reactiontime="+70" swimtime="00:20:37.31" resultid="48222" heatid="50789" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                    <SPLIT distance="100" swimtime="00:01:14.31" />
                    <SPLIT distance="150" swimtime="00:01:54.40" />
                    <SPLIT distance="200" swimtime="00:02:35.33" />
                    <SPLIT distance="250" swimtime="00:03:16.80" />
                    <SPLIT distance="300" swimtime="00:03:58.55" />
                    <SPLIT distance="350" swimtime="00:04:41.10" />
                    <SPLIT distance="400" swimtime="00:05:23.93" />
                    <SPLIT distance="450" swimtime="00:06:05.99" />
                    <SPLIT distance="500" swimtime="00:06:48.55" />
                    <SPLIT distance="550" swimtime="00:07:31.22" />
                    <SPLIT distance="600" swimtime="00:08:14.09" />
                    <SPLIT distance="650" swimtime="00:08:55.48" />
                    <SPLIT distance="700" swimtime="00:09:37.00" />
                    <SPLIT distance="750" swimtime="00:10:19.88" />
                    <SPLIT distance="800" swimtime="00:11:00.72" />
                    <SPLIT distance="850" swimtime="00:11:42.36" />
                    <SPLIT distance="900" swimtime="00:12:24.08" />
                    <SPLIT distance="950" swimtime="00:13:06.56" />
                    <SPLIT distance="1000" swimtime="00:13:48.20" />
                    <SPLIT distance="1050" swimtime="00:14:30.10" />
                    <SPLIT distance="1100" swimtime="00:15:11.01" />
                    <SPLIT distance="1150" swimtime="00:15:52.18" />
                    <SPLIT distance="1200" swimtime="00:16:33.12" />
                    <SPLIT distance="1250" swimtime="00:17:14.46" />
                    <SPLIT distance="1300" swimtime="00:17:56.74" />
                    <SPLIT distance="1350" swimtime="00:18:37.76" />
                    <SPLIT distance="1400" swimtime="00:19:19.52" />
                    <SPLIT distance="1450" swimtime="00:19:58.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="370" reactiontime="+70" swimtime="00:05:06.40" resultid="48223" heatid="50797" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                    <SPLIT distance="100" swimtime="00:01:11.36" />
                    <SPLIT distance="150" swimtime="00:01:50.39" />
                    <SPLIT distance="200" swimtime="00:02:29.25" />
                    <SPLIT distance="250" swimtime="00:03:09.07" />
                    <SPLIT distance="300" swimtime="00:03:49.23" />
                    <SPLIT distance="350" swimtime="00:04:28.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46306" points="294" reactiontime="+66" swimtime="00:01:14.38" resultid="48224" heatid="50847" lane="0" entrytime="00:01:12.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46310" points="406" reactiontime="+62" swimtime="00:00:32.39" resultid="48225" heatid="50857" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonina" lastname="Rasiewicz" birthdate="2007-07-05" gender="F" nation="POL" license="101001600305" swrid="5272054" athleteid="48309">
              <RESULTS>
                <RESULT eventid="44380" points="201" swimtime="00:01:28.15" resultid="48310" heatid="50680" lane="0" entrytime="00:01:25.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44384" points="194" reactiontime="+81" swimtime="00:00:50.77" resultid="48311" heatid="50698" lane="8" />
                <RESULT eventid="44409" points="198" reactiontime="+74" swimtime="00:01:49.96" resultid="48312" heatid="50752" lane="5" entrytime="00:01:50.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="241" reactiontime="+83" swimtime="00:00:38.01" resultid="48313" heatid="50827" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Szkirpan" birthdate="2007-09-13" gender="M" nation="POL" license="101001700297" swrid="5272056" athleteid="48340">
              <RESULTS>
                <RESULT eventid="44382" points="351" reactiontime="+65" swimtime="00:00:36.78" resultid="48341" heatid="50689" lane="2" />
                <RESULT eventid="44394" points="270" reactiontime="+78" swimtime="00:01:20.17" resultid="48342" heatid="50720" lane="6" entrytime="00:01:18.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="330" reactiontime="+60" swimtime="00:01:22.26" resultid="48343" heatid="50748" lane="5" entrytime="00:01:23.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46302" points="318" reactiontime="+55" swimtime="00:03:04.64" resultid="48344" heatid="50837" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.55" />
                    <SPLIT distance="100" swimtime="00:01:28.16" />
                    <SPLIT distance="150" swimtime="00:02:17.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46310" points="311" reactiontime="+62" swimtime="00:00:35.41" resultid="48345" heatid="50858" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksander" lastname="Cieszyński" birthdate="2007-11-18" gender="M" nation="POL" license="101001700280" swrid="5272086" athleteid="48239">
              <RESULTS>
                <RESULT eventid="44378" points="351" reactiontime="+77" swimtime="00:01:06.44" resultid="48240" heatid="50668" lane="5" entrytime="00:01:06.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="255" reactiontime="+77" swimtime="00:01:21.68" resultid="48241" heatid="50720" lane="0" entrytime="00:01:20.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="349" reactiontime="+70" swimtime="00:00:29.69" resultid="48242" heatid="50807" lane="7" />
                <RESULT eventid="46310" points="272" reactiontime="+77" swimtime="00:00:37.00" resultid="48243" heatid="50858" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Malinowski" birthdate="2006-11-19" gender="M" nation="POL" license="101001700230" swrid="5222179" athleteid="48204">
              <RESULTS>
                <RESULT eventid="44378" points="328" reactiontime="+77" swimtime="00:01:07.98" resultid="48205" heatid="50668" lane="3" entrytime="00:01:06.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="285" reactiontime="+73" swimtime="00:00:39.41" resultid="48206" heatid="50692" lane="9" />
                <RESULT eventid="44407" points="263" reactiontime="+73" swimtime="00:01:28.76" resultid="48207" heatid="50748" lane="0" entrytime="00:01:26.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46285" points="286" reactiontime="+75" swimtime="00:22:01.06" resultid="48208" heatid="50790" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                    <SPLIT distance="100" swimtime="00:01:16.83" />
                    <SPLIT distance="150" swimtime="00:01:59.71" />
                    <SPLIT distance="200" swimtime="00:02:43.74" />
                    <SPLIT distance="250" swimtime="00:03:27.62" />
                    <SPLIT distance="300" swimtime="00:04:11.94" />
                    <SPLIT distance="350" swimtime="00:04:57.03" />
                    <SPLIT distance="400" swimtime="00:05:42.13" />
                    <SPLIT distance="450" swimtime="00:06:27.18" />
                    <SPLIT distance="500" swimtime="00:07:12.62" />
                    <SPLIT distance="550" swimtime="00:07:57.21" />
                    <SPLIT distance="600" swimtime="00:08:42.24" />
                    <SPLIT distance="650" swimtime="00:09:25.69" />
                    <SPLIT distance="700" swimtime="00:10:10.19" />
                    <SPLIT distance="750" swimtime="00:10:55.26" />
                    <SPLIT distance="800" swimtime="00:11:40.19" />
                    <SPLIT distance="850" swimtime="00:12:25.44" />
                    <SPLIT distance="900" swimtime="00:13:10.62" />
                    <SPLIT distance="950" swimtime="00:13:55.58" />
                    <SPLIT distance="1000" swimtime="00:14:40.68" />
                    <SPLIT distance="1050" swimtime="00:15:25.79" />
                    <SPLIT distance="1100" swimtime="00:16:10.51" />
                    <SPLIT distance="1150" swimtime="00:16:55.35" />
                    <SPLIT distance="1200" swimtime="00:17:39.76" />
                    <SPLIT distance="1250" swimtime="00:18:23.83" />
                    <SPLIT distance="1300" swimtime="00:19:08.85" />
                    <SPLIT distance="1350" swimtime="00:19:52.45" />
                    <SPLIT distance="1400" swimtime="00:20:37.19" />
                    <SPLIT distance="1450" swimtime="00:21:19.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="317" reactiontime="+71" swimtime="00:00:30.65" resultid="48209" heatid="50809" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lena" lastname="Andrzejewska" birthdate="2007-09-23" gender="F" nation="POL" license="101001600278" swrid="5272067" athleteid="48292">
              <RESULTS>
                <RESULT eventid="44380" points="268" reactiontime="+60" swimtime="00:01:20.11" resultid="48293" heatid="50680" lane="2" entrytime="00:01:19.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44384" points="284" reactiontime="+54" swimtime="00:00:44.72" resultid="48294" heatid="50696" lane="4" />
                <RESULT eventid="44409" points="281" reactiontime="+67" swimtime="00:01:37.83" resultid="48295" heatid="50753" lane="2" entrytime="00:01:37.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46300" points="257" reactiontime="+70" swimtime="00:00:37.21" resultid="48296" heatid="50824" lane="1" />
                <RESULT eventid="46304" points="298" reactiontime="+65" swimtime="00:03:28.19" resultid="48297" heatid="50841" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.94" />
                    <SPLIT distance="100" swimtime="00:01:39.57" />
                    <SPLIT distance="150" swimtime="00:02:34.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Bonowicz" birthdate="2008-10-16" gender="M" nation="POL" license="101001700254" swrid="5341329" athleteid="48346">
              <RESULTS>
                <RESULT eventid="44382" points="219" reactiontime="+72" swimtime="00:00:43.01" resultid="48347" heatid="50692" lane="6" entrytime="00:00:47.91" entrycourse="LCM" />
                <RESULT eventid="44394" points="246" reactiontime="+77" swimtime="00:01:22.70" resultid="48348" heatid="50719" lane="3" entrytime="00:01:22.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="206" reactiontime="+68" swimtime="00:01:36.17" resultid="48349" heatid="50747" lane="8" entrytime="00:01:40.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44415" points="247" reactiontime="+95" swimtime="00:02:58.17" resultid="48350" heatid="50780" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.16" />
                    <SPLIT distance="100" swimtime="00:01:27.35" />
                    <SPLIT distance="150" swimtime="00:02:14.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46302" points="218" swimtime="00:03:29.46" resultid="48351" heatid="50836" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.19" />
                    <SPLIT distance="100" swimtime="00:01:41.34" />
                    <SPLIT distance="150" swimtime="00:02:36.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46310" points="230" reactiontime="+94" swimtime="00:00:39.13" resultid="48352" heatid="50857" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Rasiewicz" birthdate="2007-07-05" gender="M" nation="POL" license="101001700292" swrid="5272071" athleteid="48249">
              <RESULTS>
                <RESULT eventid="44378" points="345" reactiontime="+72" swimtime="00:01:06.88" resultid="48250" heatid="50669" lane="6" entrytime="00:01:05.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="291" reactiontime="+65" swimtime="00:02:33.90" resultid="48251" heatid="50733" lane="4" entrytime="00:02:34.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                    <SPLIT distance="100" swimtime="00:01:14.79" />
                    <SPLIT distance="150" swimtime="00:01:55.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46285" points="295" reactiontime="+87" swimtime="00:21:48.19" resultid="48252" heatid="50789" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.39" />
                    <SPLIT distance="100" swimtime="00:01:17.71" />
                    <SPLIT distance="150" swimtime="00:02:00.90" />
                    <SPLIT distance="200" swimtime="00:02:44.37" />
                    <SPLIT distance="250" swimtime="00:03:28.20" />
                    <SPLIT distance="300" swimtime="00:04:11.91" />
                    <SPLIT distance="350" swimtime="00:04:56.52" />
                    <SPLIT distance="400" swimtime="00:05:40.87" />
                    <SPLIT distance="450" swimtime="00:06:25.06" />
                    <SPLIT distance="500" swimtime="00:07:09.37" />
                    <SPLIT distance="550" swimtime="00:07:53.68" />
                    <SPLIT distance="600" swimtime="00:08:38.34" />
                    <SPLIT distance="650" swimtime="00:09:23.04" />
                    <SPLIT distance="700" swimtime="00:10:06.88" />
                    <SPLIT distance="750" swimtime="00:10:50.80" />
                    <SPLIT distance="800" swimtime="00:11:34.43" />
                    <SPLIT distance="850" swimtime="00:12:18.15" />
                    <SPLIT distance="900" swimtime="00:13:02.45" />
                    <SPLIT distance="950" swimtime="00:13:46.51" />
                    <SPLIT distance="1000" swimtime="00:14:30.54" />
                    <SPLIT distance="1050" swimtime="00:15:14.75" />
                    <SPLIT distance="1100" swimtime="00:15:58.99" />
                    <SPLIT distance="1150" swimtime="00:16:43.39" />
                    <SPLIT distance="1200" swimtime="00:17:27.00" />
                    <SPLIT distance="1250" swimtime="00:18:11.24" />
                    <SPLIT distance="1300" swimtime="00:18:55.15" />
                    <SPLIT distance="1350" swimtime="00:19:39.77" />
                    <SPLIT distance="1400" swimtime="00:20:23.68" />
                    <SPLIT distance="1450" swimtime="00:21:06.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="304" reactiontime="+56" swimtime="00:05:27.23" resultid="48253" heatid="50797" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.03" />
                    <SPLIT distance="100" swimtime="00:01:13.97" />
                    <SPLIT distance="150" swimtime="00:01:56.20" />
                    <SPLIT distance="200" swimtime="00:02:38.91" />
                    <SPLIT distance="250" swimtime="00:03:22.08" />
                    <SPLIT distance="300" swimtime="00:04:05.66" />
                    <SPLIT distance="350" swimtime="00:04:48.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="334" reactiontime="+70" swimtime="00:00:30.12" resultid="48254" heatid="50811" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emil" lastname="Bonowicz" birthdate="2006-01-20" gender="M" nation="POL" license="101001700219" swrid="5222176" athleteid="48210">
              <RESULTS>
                <RESULT eventid="44378" points="394" reactiontime="+69" swimtime="00:01:03.96" resultid="48211" heatid="50670" lane="3" entrytime="00:01:03.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="322" reactiontime="+70" swimtime="00:00:37.83" resultid="48212" heatid="50692" lane="0" />
                <RESULT eventid="44407" points="295" reactiontime="+72" swimtime="00:01:25.44" resultid="48213" heatid="50748" lane="3" entrytime="00:01:24.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46285" points="318" reactiontime="+69" swimtime="00:21:15.33" resultid="48214" heatid="50790" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                    <SPLIT distance="100" swimtime="00:01:13.98" />
                    <SPLIT distance="150" swimtime="00:01:54.91" />
                    <SPLIT distance="200" swimtime="00:02:37.30" />
                    <SPLIT distance="250" swimtime="00:03:19.89" />
                    <SPLIT distance="300" swimtime="00:04:02.69" />
                    <SPLIT distance="350" swimtime="00:04:46.07" />
                    <SPLIT distance="400" swimtime="00:05:29.20" />
                    <SPLIT distance="450" swimtime="00:06:12.67" />
                    <SPLIT distance="500" swimtime="00:06:55.95" />
                    <SPLIT distance="550" swimtime="00:07:39.69" />
                    <SPLIT distance="600" swimtime="00:08:23.10" />
                    <SPLIT distance="650" swimtime="00:09:06.19" />
                    <SPLIT distance="700" swimtime="00:09:48.82" />
                    <SPLIT distance="750" swimtime="00:10:32.63" />
                    <SPLIT distance="800" swimtime="00:11:15.88" />
                    <SPLIT distance="850" swimtime="00:11:59.55" />
                    <SPLIT distance="900" swimtime="00:12:42.84" />
                    <SPLIT distance="950" swimtime="00:13:26.04" />
                    <SPLIT distance="1000" swimtime="00:14:09.18" />
                    <SPLIT distance="1050" swimtime="00:14:52.27" />
                    <SPLIT distance="1100" swimtime="00:15:35.87" />
                    <SPLIT distance="1150" swimtime="00:16:19.02" />
                    <SPLIT distance="1200" swimtime="00:17:02.25" />
                    <SPLIT distance="1250" swimtime="00:17:45.52" />
                    <SPLIT distance="1300" swimtime="00:18:28.85" />
                    <SPLIT distance="1350" swimtime="00:19:11.26" />
                    <SPLIT distance="1400" swimtime="00:19:53.34" />
                    <SPLIT distance="1450" swimtime="00:20:34.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="347" reactiontime="+69" swimtime="00:00:29.74" resultid="48215" heatid="50809" lane="2" />
                <RESULT eventid="46302" points="292" reactiontime="+72" swimtime="00:03:10.00" resultid="48216" heatid="50838" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.10" />
                    <SPLIT distance="100" swimtime="00:01:29.81" />
                    <SPLIT distance="150" swimtime="00:02:20.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rozalia" lastname="Kwiatkowska" birthdate="2007-03-04" gender="F" nation="POL" license="101001600229" swrid="5222191" athleteid="48268">
              <RESULTS>
                <RESULT eventid="44380" points="496" reactiontime="+75" swimtime="00:01:05.32" resultid="48269" heatid="50686" lane="9" entrytime="00:01:04.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44392" points="447" reactiontime="+76" swimtime="00:02:44.87" resultid="48270" heatid="50715" lane="9" entrytime="00:02:45.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                    <SPLIT distance="100" swimtime="00:01:18.90" />
                    <SPLIT distance="150" swimtime="00:02:08.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44413" points="418" reactiontime="+75" swimtime="00:00:32.65" resultid="48271" heatid="50774" lane="2" entrytime="00:00:39.28" entrycourse="LCM" />
                <RESULT eventid="46300" points="534" reactiontime="+75" swimtime="00:00:29.17" resultid="48272" heatid="50829" lane="8" entrytime="00:00:34.11" entrycourse="LCM" />
                <RESULT eventid="46308" points="356" reactiontime="+81" swimtime="00:01:18.22" resultid="48273" heatid="50899" lane="3" entrytime="00:01:17.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Buchla" birthdate="2007-12-04" gender="M" nation="POL" license="101001700304" swrid="5272052" athleteid="48244">
              <RESULTS>
                <RESULT eventid="44378" points="266" reactiontime="+65" swimtime="00:01:12.94" resultid="48245" heatid="50665" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46285" points="238" reactiontime="+64" swimtime="00:23:23.80" resultid="48246" heatid="50790" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                    <SPLIT distance="100" swimtime="00:01:19.78" />
                    <SPLIT distance="150" swimtime="00:02:04.93" />
                    <SPLIT distance="200" swimtime="00:02:49.11" />
                    <SPLIT distance="250" swimtime="00:03:36.12" />
                    <SPLIT distance="300" swimtime="00:04:22.54" />
                    <SPLIT distance="350" swimtime="00:05:10.65" />
                    <SPLIT distance="400" swimtime="00:05:58.93" />
                    <SPLIT distance="450" swimtime="00:06:46.60" />
                    <SPLIT distance="500" swimtime="00:07:34.64" />
                    <SPLIT distance="550" swimtime="00:08:22.51" />
                    <SPLIT distance="600" swimtime="00:09:08.74" />
                    <SPLIT distance="650" swimtime="00:09:58.08" />
                    <SPLIT distance="700" swimtime="00:10:45.60" />
                    <SPLIT distance="750" swimtime="00:11:33.68" />
                    <SPLIT distance="800" swimtime="00:12:21.96" />
                    <SPLIT distance="850" swimtime="00:13:09.35" />
                    <SPLIT distance="900" swimtime="00:13:57.13" />
                    <SPLIT distance="950" swimtime="00:14:45.16" />
                    <SPLIT distance="1000" swimtime="00:15:33.73" />
                    <SPLIT distance="1050" swimtime="00:16:21.57" />
                    <SPLIT distance="1100" swimtime="00:17:09.49" />
                    <SPLIT distance="1150" swimtime="00:17:56.46" />
                    <SPLIT distance="1200" swimtime="00:18:45.07" />
                    <SPLIT distance="1250" swimtime="00:19:31.90" />
                    <SPLIT distance="1300" swimtime="00:20:19.21" />
                    <SPLIT distance="1350" swimtime="00:21:06.28" />
                    <SPLIT distance="1400" swimtime="00:21:52.88" />
                    <SPLIT distance="1450" swimtime="00:22:38.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="283" swimtime="00:00:31.83" resultid="48247" heatid="50806" lane="4" />
                <RESULT eventid="46310" points="242" reactiontime="+57" swimtime="00:00:38.51" resultid="48248" heatid="50856" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antoni" lastname="Makowiecki" birthdate="2008-06-18" gender="M" nation="POL" license="101001700264" swrid="5341297" athleteid="48255">
              <RESULTS>
                <RESULT eventid="44378" points="380" reactiontime="+79" swimtime="00:01:04.71" resultid="48256" heatid="50670" lane="9" entrytime="00:01:04.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44394" points="303" reactiontime="+80" swimtime="00:01:17.16" resultid="48257" heatid="50720" lane="4" entrytime="00:01:17.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="331" reactiontime="+79" swimtime="00:02:27.45" resultid="48258" heatid="50734" lane="9" entrytime="00:02:34.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                    <SPLIT distance="100" swimtime="00:01:10.35" />
                    <SPLIT distance="150" swimtime="00:01:50.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="265" reactiontime="+81" swimtime="00:00:34.67" resultid="48259" heatid="50762" lane="6" entrytime="00:00:38.01" entrycourse="LCM" />
                <RESULT eventid="46298" points="363" reactiontime="+74" swimtime="00:00:29.29" resultid="48260" heatid="50814" lane="7" entrytime="00:00:32.52" entrycourse="LCM" />
                <RESULT eventid="46310" points="332" reactiontime="+71" swimtime="00:00:34.64" resultid="48261" heatid="50855" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartłomiej" lastname="Kaśków" birthdate="2006-03-11" gender="M" nation="POL" license="101001700226" swrid="5222184" athleteid="48226">
              <RESULTS>
                <RESULT eventid="44378" points="497" reactiontime="+78" swimtime="00:00:59.19" resultid="48227" heatid="50663" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44382" points="466" reactiontime="+75" swimtime="00:00:33.47" resultid="48228" heatid="50690" lane="1" />
                <RESULT eventid="44390" points="363" reactiontime="+83" swimtime="00:02:39.70" resultid="48229" heatid="50708" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                    <SPLIT distance="100" swimtime="00:01:17.61" />
                    <SPLIT distance="150" swimtime="00:02:03.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44407" points="397" reactiontime="+77" swimtime="00:01:17.34" resultid="48230" heatid="50749" lane="6" entrytime="00:01:17.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46294" points="366" reactiontime="+76" swimtime="00:05:07.39" resultid="48231" heatid="50796" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="100" swimtime="00:01:08.86" />
                    <SPLIT distance="150" swimtime="00:01:48.26" />
                    <SPLIT distance="200" swimtime="00:02:28.82" />
                    <SPLIT distance="250" swimtime="00:03:10.61" />
                    <SPLIT distance="300" swimtime="00:03:52.17" />
                    <SPLIT distance="350" swimtime="00:04:31.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46298" points="487" reactiontime="+78" swimtime="00:00:26.57" resultid="48232" heatid="50810" lane="2" />
                <RESULT eventid="46302" points="380" reactiontime="+78" swimtime="00:02:54.09" resultid="48233" heatid="50837" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.59" />
                    <SPLIT distance="100" swimtime="00:01:24.62" />
                    <SPLIT distance="150" swimtime="00:02:10.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maja" lastname="Ryczek" birthdate="2007-01-30" gender="F" nation="POL" license="101001600306" swrid="5272088" athleteid="48375">
              <RESULTS>
                <RESULT eventid="44396" points="320" reactiontime="+69" swimtime="00:01:24.15" resultid="48376" heatid="50726" lane="0" entrytime="00:01:23.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44417" points="323" reactiontime="+72" swimtime="00:02:59.61" resultid="48377" heatid="50786" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.69" />
                    <SPLIT distance="100" swimtime="00:01:29.60" />
                    <SPLIT distance="150" swimtime="00:02:16.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46312" points="338" reactiontime="+76" swimtime="00:00:38.70" resultid="48378" heatid="50904" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emilia" lastname="Weselska" birthdate="2008-12-17" gender="F" nation="POL" license="101001600275" swrid="5341320" athleteid="48320">
              <RESULTS>
                <RESULT eventid="44380" points="435" reactiontime="+73" swimtime="00:01:08.20" resultid="48321" heatid="50683" lane="6" entrytime="00:01:08.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44384" points="436" reactiontime="+77" swimtime="00:00:38.75" resultid="48322" heatid="50700" lane="3" entrytime="00:00:43.79" entrycourse="LCM" />
                <RESULT eventid="44405" points="398" reactiontime="+85" swimtime="00:02:33.47" resultid="48323" heatid="50741" lane="6" entrytime="00:02:34.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.24" />
                    <SPLIT distance="100" swimtime="00:01:14.71" />
                    <SPLIT distance="150" swimtime="00:01:55.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44409" points="440" reactiontime="+74" swimtime="00:01:24.28" resultid="48324" heatid="50754" lane="3" entrytime="00:01:25.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46287" points="355" reactiontime="+76" swimtime="00:11:24.46" resultid="48325" heatid="50791" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                    <SPLIT distance="100" swimtime="00:01:18.50" />
                    <SPLIT distance="150" swimtime="00:02:01.63" />
                    <SPLIT distance="200" swimtime="00:02:45.02" />
                    <SPLIT distance="250" swimtime="00:03:28.51" />
                    <SPLIT distance="300" swimtime="00:04:12.09" />
                    <SPLIT distance="350" swimtime="00:04:55.58" />
                    <SPLIT distance="400" swimtime="00:05:39.72" />
                    <SPLIT distance="450" swimtime="00:06:23.33" />
                    <SPLIT distance="500" swimtime="00:07:07.10" />
                    <SPLIT distance="550" swimtime="00:07:50.62" />
                    <SPLIT distance="600" swimtime="00:08:34.57" />
                    <SPLIT distance="650" swimtime="00:09:17.72" />
                    <SPLIT distance="700" swimtime="00:10:00.93" />
                    <SPLIT distance="750" swimtime="00:10:43.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46304" points="456" reactiontime="+55" swimtime="00:03:00.61" resultid="48326" heatid="50841" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.60" />
                    <SPLIT distance="100" swimtime="00:01:27.37" />
                    <SPLIT distance="150" swimtime="00:02:15.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="44399" points="354" reactiontime="+91" swimtime="00:04:52.83" resultid="48379" heatid="50730" lane="1" entrytime="00:04:46.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.24" />
                    <SPLIT distance="100" swimtime="00:01:18.67" />
                    <SPLIT distance="150" swimtime="00:01:55.29" />
                    <SPLIT distance="200" swimtime="00:02:37.92" />
                    <SPLIT distance="250" swimtime="00:03:08.97" />
                    <SPLIT distance="300" swimtime="00:03:49.88" />
                    <SPLIT distance="350" swimtime="00:04:19.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="48204" number="1" reactiontime="+91" />
                    <RELAYPOSITION athleteid="48226" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="48217" number="3" reactiontime="+25" />
                    <RELAYPOSITION athleteid="48210" number="4" reactiontime="+14" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46289" points="345" reactiontime="+56" swimtime="00:04:28.20" resultid="48382" heatid="50794" lane="9" entrytime="00:04:10.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                    <SPLIT distance="100" swimtime="00:01:06.39" />
                    <SPLIT distance="150" swimtime="00:01:39.59" />
                    <SPLIT distance="200" swimtime="00:02:17.26" />
                    <SPLIT distance="250" swimtime="00:02:50.04" />
                    <SPLIT distance="300" swimtime="00:03:28.31" />
                    <SPLIT distance="350" swimtime="00:03:56.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="48217" number="1" reactiontime="+56" />
                    <RELAYPOSITION athleteid="48204" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="48210" number="3" reactiontime="+9" />
                    <RELAYPOSITION athleteid="48226" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="44399" points="326" reactiontime="+66" swimtime="00:05:01.14" resultid="48380" heatid="50730" lane="0" entrytime="00:04:53.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                    <SPLIT distance="100" swimtime="00:01:15.50" />
                    <SPLIT distance="150" swimtime="00:01:54.37" />
                    <SPLIT distance="200" swimtime="00:02:39.16" />
                    <SPLIT distance="250" swimtime="00:03:12.91" />
                    <SPLIT distance="300" swimtime="00:03:54.71" />
                    <SPLIT distance="350" swimtime="00:04:25.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="48370" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="48340" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="48234" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="48239" number="4" reactiontime="+4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46289" points="356" reactiontime="+82" swimtime="00:04:25.43" resultid="48383" heatid="50793" lane="3" entrytime="00:04:16.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                    <SPLIT distance="100" swimtime="00:01:06.40" />
                    <SPLIT distance="150" swimtime="00:01:38.10" />
                    <SPLIT distance="200" swimtime="00:02:13.60" />
                    <SPLIT distance="250" swimtime="00:02:43.94" />
                    <SPLIT distance="300" swimtime="00:03:20.13" />
                    <SPLIT distance="350" swimtime="00:03:51.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="48249" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="48234" number="2" />
                    <RELAYPOSITION athleteid="48239" number="3" />
                    <RELAYPOSITION athleteid="48340" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="44401" points="321" reactiontime="+70" swimtime="00:05:36.37" resultid="48381" heatid="50731" lane="2" entrytime="00:05:16.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.90" />
                    <SPLIT distance="100" swimtime="00:01:24.89" />
                    <SPLIT distance="150" swimtime="00:02:07.39" />
                    <SPLIT distance="200" swimtime="00:02:57.25" />
                    <SPLIT distance="250" swimtime="00:03:35.16" />
                    <SPLIT distance="300" swimtime="00:04:32.98" />
                    <SPLIT distance="350" swimtime="00:05:00.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="48375" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="48358" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="48353" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="48268" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="46291" points="377" reactiontime="+63" swimtime="00:04:50.55" resultid="48384" heatid="50795" lane="0" entrytime="00:04:35.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                    <SPLIT distance="100" swimtime="00:01:10.01" />
                    <SPLIT distance="150" swimtime="00:01:45.82" />
                    <SPLIT distance="200" swimtime="00:02:27.56" />
                    <SPLIT distance="250" swimtime="00:03:04.15" />
                    <SPLIT distance="300" swimtime="00:03:45.04" />
                    <SPLIT distance="350" swimtime="00:04:15.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="48314" number="1" reactiontime="+63" />
                    <RELAYPOSITION athleteid="48375" number="2" />
                    <RELAYPOSITION athleteid="48353" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="48268" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="06614" nation="POL" region="14" clubid="47004" name="Legia Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Jan" lastname="Marczewski" birthdate="2004-09-08" gender="M" nation="POL" license="106614700091" swrid="5403857" athleteid="47012">
              <RESULTS>
                <RESULT eventid="44382" points="411" reactiontime="+70" swimtime="00:00:34.90" resultid="47013" heatid="50694" lane="1" entrytime="00:00:34.07" entrycourse="LCM" />
                <RESULT eventid="44407" points="328" reactiontime="+71" swimtime="00:01:22.42" resultid="47014" heatid="50749" lane="0" entrytime="00:01:20.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="352" reactiontime="+69" swimtime="00:00:31.53" resultid="47015" heatid="50760" lane="4" />
                <RESULT eventid="46298" points="414" reactiontime="+66" swimtime="00:00:28.04" resultid="47016" heatid="50815" lane="8" entrytime="00:00:30.42" entrycourse="LCM" />
                <RESULT eventid="46302" status="DNS" swimtime="00:00:00.00" resultid="47017" heatid="50837" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stefan" lastname="Dobrowolski" birthdate="2005-07-31" gender="M" nation="POL" license="106614700076" swrid="5115033" athleteid="47005">
              <RESULTS>
                <RESULT eventid="44378" points="473" reactiontime="+75" swimtime="00:01:00.17" resultid="47006" heatid="50671" lane="6" entrytime="00:01:02.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44390" points="425" reactiontime="+73" swimtime="00:02:31.57" resultid="47007" heatid="50708" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                    <SPLIT distance="100" swimtime="00:01:10.95" />
                    <SPLIT distance="150" swimtime="00:01:56.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44403" points="418" reactiontime="+74" swimtime="00:02:16.37" resultid="47008" heatid="50735" lane="3" entrytime="00:02:25.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                    <SPLIT distance="100" swimtime="00:01:06.47" />
                    <SPLIT distance="150" swimtime="00:01:42.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44411" points="429" reactiontime="+72" swimtime="00:00:29.51" resultid="47009" heatid="50759" lane="2" />
                <RESULT eventid="46298" points="464" reactiontime="+75" swimtime="00:00:27.00" resultid="47010" heatid="50818" lane="1" entrytime="00:00:27.15" entrycourse="LCM" />
                <RESULT eventid="46306" points="339" reactiontime="+55" swimtime="00:01:10.95" resultid="47011" heatid="50844" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>

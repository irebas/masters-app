<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="KSP Katowice" version="11.72268">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Katowice" name="Puchar Polski Masters w Pływaniu" course="SCM" deadline="2022-05-05" hostclub="Wodnik 29 Katowice" organizer="Wodnik 29 Katowice" reservecount="2" startmethod="1" timing="AUTOMATIC" nation="POL" maxentriesathlete="4">
      <AGEDATE value="2022-05-14" type="YEAR" />
      <POOL name="Katowice" lanemin="1" lanemax="6" />
      <FACILITY city="Katowice" name="Katowice" nation="POL" street="Kościuszki" />
      <POINTTABLE pointtableid="997" name="MASTERS FINA WR" version="2022" />
      <CONTACT city="Katowice" email="zawody.jczarnecki@gmail.com" />
      <SESSIONS>
        <SESSION date="2022-05-14" daytime="10:00" endtime="13:41" number="1" warmupfrom="09:00" warmupuntil="09:45">
          <EVENTS>
            <EVENT eventid="1059" daytime="10:00" gender="F" number="1" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1061" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3607" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1062" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3108" />
                    <RANKING order="2" place="2" resultid="2919" />
                    <RANKING order="3" place="3" resultid="3052" />
                    <RANKING order="4" place="4" resultid="2243" />
                    <RANKING order="5" place="-1" resultid="3113" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1063" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2715" />
                    <RANKING order="2" place="2" resultid="3064" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1064" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2852" />
                    <RANKING order="2" place="2" resultid="3283" />
                    <RANKING order="3" place="3" resultid="2625" />
                    <RANKING order="4" place="-1" resultid="2849" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2534" />
                    <RANKING order="2" place="2" resultid="3822" />
                    <RANKING order="3" place="3" resultid="2630" />
                    <RANKING order="4" place="4" resultid="2640" />
                    <RANKING order="5" place="5" resultid="2539" />
                    <RANKING order="6" place="6" resultid="2477" />
                    <RANKING order="7" place="7" resultid="2544" />
                    <RANKING order="8" place="8" resultid="3413" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3420" />
                    <RANKING order="2" place="2" resultid="3334" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3377" />
                    <RANKING order="2" place="2" resultid="2157" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1068" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2570" />
                    <RANKING order="2" place="2" resultid="3150" />
                    <RANKING order="3" place="3" resultid="2337" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3372" />
                    <RANKING order="2" place="2" resultid="2635" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69" />
                <AGEGROUP agegroupid="1071" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3551" />
                    <RANKING order="2" place="2" resultid="3518" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1072" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2401" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1073" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3194" />
                    <RANKING order="2" place="2" resultid="3837" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4818" agemax="-1" agemin="20" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3108" />
                    <RANKING order="2" place="2" resultid="2919" />
                    <RANKING order="3" place="3" resultid="3052" />
                    <RANKING order="4" place="4" resultid="2534" />
                    <RANKING order="5" place="5" resultid="2715" />
                    <RANKING order="6" place="6" resultid="2852" />
                    <RANKING order="7" place="7" resultid="3822" />
                    <RANKING order="8" place="8" resultid="3607" />
                    <RANKING order="9" place="9" resultid="2243" />
                    <RANKING order="10" place="10" resultid="2570" />
                    <RANKING order="11" place="11" resultid="2630" />
                    <RANKING order="12" place="12" resultid="2640" />
                    <RANKING order="13" place="13" resultid="3064" />
                    <RANKING order="14" place="14" resultid="3377" />
                    <RANKING order="15" place="15" resultid="3372" />
                    <RANKING order="16" place="16" resultid="3150" />
                    <RANKING order="17" place="17" resultid="2337" />
                    <RANKING order="18" place="18" resultid="2157" />
                    <RANKING order="19" place="19" resultid="3283" />
                    <RANKING order="20" place="20" resultid="2539" />
                    <RANKING order="21" place="21" resultid="2477" />
                    <RANKING order="22" place="22" resultid="3420" />
                    <RANKING order="23" place="23" resultid="2544" />
                    <RANKING order="24" place="24" resultid="2625" />
                    <RANKING order="25" place="25" resultid="3551" />
                    <RANKING order="26" place="26" resultid="2635" />
                    <RANKING order="27" place="27" resultid="3413" />
                    <RANKING order="28" place="28" resultid="3518" />
                    <RANKING order="29" place="29" resultid="3334" />
                    <RANKING order="30" place="30" resultid="3194" />
                    <RANKING order="31" place="31" resultid="2401" />
                    <RANKING order="32" place="32" resultid="3837" />
                    <RANKING order="33" place="-1" resultid="2849" />
                    <RANKING order="34" place="-1" resultid="3113" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4664" daytime="10:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4665" daytime="10:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4666" daytime="10:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4667" daytime="10:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4668" daytime="10:05" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4669" daytime="10:10" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1102" daytime="10:10" gender="M" number="2" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1116" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3079" />
                    <RANKING order="2" place="2" resultid="3158" />
                    <RANKING order="3" place="3" resultid="2559" />
                    <RANKING order="4" place="4" resultid="2376" />
                    <RANKING order="5" place="5" resultid="2367" />
                    <RANKING order="6" place="6" resultid="3163" />
                    <RANKING order="7" place="7" resultid="2186" />
                    <RANKING order="8" place="8" resultid="2898" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1117" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2793" />
                    <RANKING order="2" place="2" resultid="3088" />
                    <RANKING order="3" place="3" resultid="3098" />
                    <RANKING order="4" place="4" resultid="3250" />
                    <RANKING order="5" place="5" resultid="2168" />
                    <RANKING order="6" place="6" resultid="3428" />
                    <RANKING order="7" place="7" resultid="3103" />
                    <RANKING order="8" place="8" resultid="2615" />
                    <RANKING order="9" place="9" resultid="2435" />
                    <RANKING order="10" place="10" resultid="3620" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1118" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3068" />
                    <RANKING order="2" place="2" resultid="3156" />
                    <RANKING order="3" place="3" resultid="3319" />
                    <RANKING order="4" place="4" resultid="2465" />
                    <RANKING order="5" place="5" resultid="3118" />
                    <RANKING order="6" place="6" resultid="2878" />
                    <RANKING order="7" place="7" resultid="2422" />
                    <RANKING order="8" place="8" resultid="3630" />
                    <RANKING order="9" place="9" resultid="2883" />
                    <RANKING order="10" place="10" resultid="2417" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1119" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2430" />
                    <RANKING order="2" place="2" resultid="2344" />
                    <RANKING order="3" place="3" resultid="3666" />
                    <RANKING order="4" place="4" resultid="3076" />
                    <RANKING order="5" place="5" resultid="2888" />
                    <RANKING order="6" place="6" resultid="2425" />
                    <RANKING order="7" place="-1" resultid="2162" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1120" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3142" />
                    <RANKING order="2" place="2" resultid="3309" />
                    <RANKING order="3" place="3" resultid="2815" />
                    <RANKING order="4" place="4" resultid="3408" />
                    <RANKING order="5" place="5" resultid="3616" />
                    <RANKING order="6" place="6" resultid="2193" />
                    <RANKING order="7" place="7" resultid="2372" />
                    <RANKING order="8" place="8" resultid="2657" />
                    <RANKING order="9" place="-1" resultid="3133" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1121" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3498" />
                    <RANKING order="2" place="2" resultid="2824" />
                    <RANKING order="3" place="3" resultid="2565" />
                    <RANKING order="4" place="4" resultid="3294" />
                    <RANKING order="5" place="5" resultid="2215" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1122" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2605" />
                    <RANKING order="2" place="2" resultid="3358" />
                    <RANKING order="3" place="3" resultid="3433" />
                    <RANKING order="4" place="4" resultid="2482" />
                    <RANKING order="5" place="5" resultid="3561" />
                    <RANKING order="6" place="6" resultid="3645" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1123" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3205" />
                    <RANKING order="2" place="2" resultid="2209" />
                    <RANKING order="3" place="3" resultid="3502" />
                    <RANKING order="4" place="4" resultid="2862" />
                    <RANKING order="5" place="5" resultid="2590" />
                    <RANKING order="6" place="6" resultid="3041" />
                    <RANKING order="7" place="7" resultid="3566" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1124" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3466" />
                    <RANKING order="2" place="2" resultid="2585" />
                    <RANKING order="3" place="3" resultid="3171" />
                    <RANKING order="4" place="4" resultid="3403" />
                    <RANKING order="5" place="5" resultid="2226" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1125" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3395" />
                    <RANKING order="2" place="2" resultid="3845" />
                    <RANKING order="3" place="3" resultid="2669" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1126" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3527" />
                    <RANKING order="2" place="2" resultid="2199" />
                    <RANKING order="3" place="3" resultid="3354" />
                    <RANKING order="4" place="4" resultid="3536" />
                    <RANKING order="5" place="5" resultid="3226" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1127" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2580" />
                    <RANKING order="2" place="2" resultid="2174" />
                    <RANKING order="3" place="3" resultid="2406" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1128" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi" />
                <AGEGROUP agegroupid="4819" agemax="-1" agemin="20" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3079" />
                    <RANKING order="2" place="2" resultid="3068" />
                    <RANKING order="3" place="3" resultid="2793" />
                    <RANKING order="4" place="4" resultid="3158" />
                    <RANKING order="5" place="5" resultid="3088" />
                    <RANKING order="6" place="6" resultid="3156" />
                    <RANKING order="7" place="7" resultid="3098" />
                    <RANKING order="8" place="8" resultid="2559" />
                    <RANKING order="9" place="9" resultid="2376" />
                    <RANKING order="10" place="10" resultid="3319" />
                    <RANKING order="11" place="11" resultid="3250" />
                    <RANKING order="12" place="12" resultid="2168" />
                    <RANKING order="13" place="13" resultid="2367" />
                    <RANKING order="14" place="14" resultid="3142" />
                    <RANKING order="15" place="15" resultid="3163" />
                    <RANKING order="16" place="16" resultid="3309" />
                    <RANKING order="17" place="17" resultid="2186" />
                    <RANKING order="18" place="18" resultid="2898" />
                    <RANKING order="19" place="19" resultid="2465" />
                    <RANKING order="20" place="19" resultid="2605" />
                    <RANKING order="21" place="21" resultid="3428" />
                    <RANKING order="22" place="22" resultid="3498" />
                    <RANKING order="23" place="23" resultid="3103" />
                    <RANKING order="24" place="24" resultid="3118" />
                    <RANKING order="25" place="25" resultid="2430" />
                    <RANKING order="26" place="26" resultid="2878" />
                    <RANKING order="27" place="27" resultid="3205" />
                    <RANKING order="28" place="28" resultid="2615" />
                    <RANKING order="29" place="29" resultid="3466" />
                    <RANKING order="30" place="30" resultid="2344" />
                    <RANKING order="31" place="31" resultid="2209" />
                    <RANKING order="32" place="32" resultid="3502" />
                    <RANKING order="33" place="33" resultid="2435" />
                    <RANKING order="34" place="34" resultid="3666" />
                    <RANKING order="35" place="35" resultid="3620" />
                    <RANKING order="36" place="36" resultid="2422" />
                    <RANKING order="37" place="37" resultid="2585" />
                    <RANKING order="38" place="38" resultid="2862" />
                    <RANKING order="39" place="39" resultid="3358" />
                    <RANKING order="40" place="40" resultid="3171" />
                    <RANKING order="41" place="41" resultid="2815" />
                    <RANKING order="42" place="42" resultid="3433" />
                    <RANKING order="43" place="43" resultid="2482" />
                    <RANKING order="44" place="44" resultid="3561" />
                    <RANKING order="45" place="45" resultid="2590" />
                    <RANKING order="46" place="46" resultid="2824" />
                    <RANKING order="47" place="47" resultid="3630" />
                    <RANKING order="48" place="48" resultid="3395" />
                    <RANKING order="49" place="49" resultid="2565" />
                    <RANKING order="50" place="50" resultid="3076" />
                    <RANKING order="51" place="51" resultid="3294" />
                    <RANKING order="52" place="52" resultid="3527" />
                    <RANKING order="53" place="53" resultid="2215" />
                    <RANKING order="54" place="54" resultid="3408" />
                    <RANKING order="55" place="55" resultid="2888" />
                    <RANKING order="56" place="56" resultid="3616" />
                    <RANKING order="57" place="57" resultid="3403" />
                    <RANKING order="58" place="58" resultid="2883" />
                    <RANKING order="59" place="59" resultid="2193" />
                    <RANKING order="60" place="59" resultid="3845" />
                    <RANKING order="61" place="61" resultid="2425" />
                    <RANKING order="62" place="62" resultid="2372" />
                    <RANKING order="63" place="63" resultid="2417" />
                    <RANKING order="64" place="64" resultid="2580" />
                    <RANKING order="65" place="65" resultid="2174" />
                    <RANKING order="66" place="66" resultid="3645" />
                    <RANKING order="67" place="67" resultid="2226" />
                    <RANKING order="68" place="68" resultid="3041" />
                    <RANKING order="69" place="69" resultid="2657" />
                    <RANKING order="70" place="70" resultid="2199" />
                    <RANKING order="71" place="71" resultid="2669" />
                    <RANKING order="72" place="72" resultid="3354" />
                    <RANKING order="73" place="73" resultid="3536" />
                    <RANKING order="74" place="74" resultid="3226" />
                    <RANKING order="75" place="75" resultid="2406" />
                    <RANKING order="76" place="76" resultid="3566" />
                    <RANKING order="77" place="-1" resultid="2162" />
                    <RANKING order="78" place="-1" resultid="3133" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4670" daytime="10:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4671" daytime="10:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4672" daytime="10:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4673" daytime="10:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4674" daytime="10:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4675" daytime="10:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4676" daytime="10:20" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4677" daytime="10:20" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4678" daytime="10:20" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4679" daytime="10:20" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4680" daytime="10:25" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4681" daytime="10:25" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="4682" daytime="10:25" number="13" order="13" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1129" daytime="10:30" gender="F" number="3" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1130" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3215" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1131" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3260" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1132" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3268" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1133" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2829" />
                    <RANKING order="2" place="2" resultid="2807" />
                    <RANKING order="3" place="3" resultid="3825" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1134" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2535" />
                    <RANKING order="2" place="2" resultid="2631" />
                    <RANKING order="3" place="-1" resultid="3584" />
                    <RANKING order="4" place="-1" resultid="3839" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1135" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49" />
                <AGEGROUP agegroupid="1136" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3378" />
                    <RANKING order="2" place="2" resultid="3852" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1137" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2699" />
                    <RANKING order="2" place="2" resultid="3329" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1138" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2450" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1139" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2310" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1140" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3552" />
                    <RANKING order="2" place="2" resultid="3519" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1141" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="1142" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4683" daytime="10:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4684" daytime="10:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4685" daytime="10:35" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1143" daytime="10:35" gender="M" number="4" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1144" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2549" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1145" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3245" />
                    <RANKING order="2" place="2" resultid="3099" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1146" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3093" />
                    <RANKING order="2" place="2" resultid="2466" />
                    <RANKING order="3" place="3" resultid="2610" />
                    <RANKING order="4" place="4" resultid="3290" />
                    <RANKING order="5" place="-1" resultid="3573" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1147" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3578" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1148" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2857" />
                    <RANKING order="2" place="2" resultid="2471" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1149" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2839" />
                    <RANKING order="2" place="2" resultid="3338" />
                    <RANKING order="3" place="3" resultid="3479" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1150" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2674" />
                    <RANKING order="2" place="2" resultid="3232" />
                    <RANKING order="3" place="3" resultid="2180" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1151" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3046" />
                    <RANKING order="2" place="-1" resultid="3456" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1152" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3272" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1153" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3484" />
                    <RANKING order="2" place="2" resultid="3556" />
                    <RANKING order="3" place="3" resultid="2393" />
                    <RANKING order="4" place="-1" resultid="3513" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1154" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3355" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1155" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3509" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1156" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2386" />
                    <RANKING order="2" place="2" resultid="2397" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4686" daytime="10:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4687" daytime="10:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4688" daytime="10:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4689" daytime="10:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4690" daytime="10:45" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1157" daytime="10:50" gender="F" number="5" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1158" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3175" />
                    <RANKING order="2" place="2" resultid="2341" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1159" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2834" />
                    <RANKING order="2" place="2" resultid="3255" />
                    <RANKING order="3" place="3" resultid="2920" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1160" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34" />
                <AGEGROUP agegroupid="1161" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2853" />
                    <RANKING order="2" place="2" resultid="2801" />
                    <RANKING order="3" place="3" resultid="3656" />
                    <RANKING order="4" place="4" resultid="2914" />
                    <RANKING order="5" place="5" resultid="3185" />
                    <RANKING order="6" place="6" resultid="3211" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1162" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3601" />
                    <RANKING order="2" place="2" resultid="3642" />
                    <RANKING order="3" place="3" resultid="2540" />
                    <RANKING order="4" place="4" resultid="2545" />
                    <RANKING order="5" place="5" resultid="3414" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1163" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3368" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1164" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3032" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1165" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2571" />
                    <RANKING order="2" place="2" resultid="2338" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1166" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3373" />
                    <RANKING order="2" place="2" resultid="3201" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1167" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69" />
                <AGEGROUP agegroupid="1168" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3523" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1169" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="1170" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4691" daytime="10:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4692" daytime="10:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4693" daytime="10:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4694" daytime="10:55" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1171" daytime="10:55" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1172" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2560" />
                    <RANKING order="2" place="2" resultid="3610" />
                    <RANKING order="3" place="3" resultid="2368" />
                    <RANKING order="4" place="4" resultid="3164" />
                    <RANKING order="5" place="5" resultid="2187" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1173" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3263" />
                    <RANKING order="2" place="2" resultid="2844" />
                    <RANKING order="3" place="3" resultid="3429" />
                    <RANKING order="4" place="4" resultid="2893" />
                    <RANKING order="5" place="5" resultid="3104" />
                    <RANKING order="6" place="6" resultid="2436" />
                    <RANKING order="7" place="7" resultid="2616" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1174" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3424" />
                    <RANKING order="2" place="2" resultid="2819" />
                    <RANKING order="3" place="3" resultid="3833" />
                    <RANKING order="4" place="4" resultid="3239" />
                    <RANKING order="5" place="5" resultid="2611" />
                    <RANKING order="6" place="6" resultid="2884" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1175" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3568" />
                    <RANKING order="2" place="2" resultid="3474" />
                    <RANKING order="3" place="3" resultid="2237" />
                    <RANKING order="4" place="4" resultid="2889" />
                    <RANKING order="5" place="5" resultid="2459" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1176" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3310" />
                    <RANKING order="2" place="2" resultid="3471" />
                    <RANKING order="3" place="3" resultid="4007" />
                    <RANKING order="4" place="4" resultid="3437" />
                    <RANKING order="5" place="5" resultid="2194" />
                    <RANKING order="6" place="6" resultid="3409" />
                    <RANKING order="7" place="-1" resultid="3134" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1177" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3488" />
                    <RANKING order="2" place="2" resultid="2332" />
                    <RANKING order="3" place="3" resultid="3138" />
                    <RANKING order="4" place="4" resultid="3278" />
                    <RANKING order="5" place="5" resultid="2825" />
                    <RANKING order="6" place="6" resultid="2529" />
                    <RANKING order="7" place="-1" resultid="2216" />
                    <RANKING order="8" place="-1" resultid="3382" />
                    <RANKING order="9" place="-1" resultid="3461" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1178" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2362" />
                    <RANKING order="2" place="2" resultid="2606" />
                    <RANKING order="3" place="3" resultid="2661" />
                    <RANKING order="4" place="4" resultid="2181" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1179" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2591" />
                    <RANKING order="2" place="2" resultid="3042" />
                    <RANKING order="3" place="3" resultid="3037" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1180" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3167" />
                    <RANKING order="2" place="2" resultid="2586" />
                    <RANKING order="3" place="3" resultid="3324" />
                    <RANKING order="4" place="4" resultid="3634" />
                    <RANKING order="5" place="5" resultid="3404" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1181" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3390" />
                    <RANKING order="2" place="-1" resultid="4816" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1182" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74" />
                <AGEGROUP agegroupid="1183" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3130" />
                    <RANKING order="2" place="2" resultid="2407" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1184" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3834" />
                    <RANKING order="2" place="2" resultid="2390" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4695" daytime="10:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4696" daytime="11:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4697" daytime="11:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4698" daytime="11:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4699" daytime="11:05" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4700" daytime="11:05" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4701" daytime="11:05" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4702" daytime="11:05" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4703" daytime="11:10" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4704" daytime="11:10" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1185" daytime="11:10" gender="F" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1186" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24" />
                <AGEGROUP agegroupid="1187" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3053" />
                    <RANKING order="2" place="2" resultid="2326" />
                    <RANKING order="3" place="3" resultid="3114" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1188" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34" />
                <AGEGROUP agegroupid="1189" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2808" />
                    <RANKING order="2" place="2" resultid="3018" />
                    <RANKING order="3" place="3" resultid="3284" />
                    <RANKING order="4" place="4" resultid="2413" />
                    <RANKING order="5" place="5" resultid="2221" />
                    <RANKING order="6" place="6" resultid="3826" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1190" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2205" />
                    <RANKING order="2" place="-1" resultid="3585" />
                    <RANKING order="3" place="-1" resultid="3840" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1191" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3659" />
                    <RANKING order="2" place="2" resultid="3421" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1192" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3539" />
                    <RANKING order="2" place="-1" resultid="2600" />
                    <RANKING order="3" place="-1" resultid="3190" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1193" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3151" />
                    <RANKING order="2" place="2" resultid="3330" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1194" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2595" />
                    <RANKING order="2" place="2" resultid="2451" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1195" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69" />
                <AGEGROUP agegroupid="1196" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74" />
                <AGEGROUP agegroupid="1197" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2402" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1198" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4705" daytime="11:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4706" daytime="11:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4707" daytime="11:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4708" daytime="11:25" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1199" daytime="11:30" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1200" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3159" />
                    <RANKING order="2" place="2" resultid="2377" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1201" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3621" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1202" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2350" />
                    <RANKING order="2" place="2" resultid="3320" />
                    <RANKING order="3" place="-1" resultid="3119" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1203" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2345" />
                    <RANKING order="2" place="2" resultid="3667" />
                    <RANKING order="3" place="-1" resultid="2164" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1204" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3314" />
                    <RANKING order="2" place="2" resultid="3617" />
                    <RANKING order="3" place="3" resultid="2373" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1205" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3499" />
                    <RANKING order="2" place="2" resultid="3339" />
                    <RANKING order="3" place="-1" resultid="3462" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1206" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3359" />
                    <RANKING order="2" place="2" resultid="3562" />
                    <RANKING order="3" place="3" resultid="3058" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1207" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3503" />
                    <RANKING order="2" place="2" resultid="3047" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1208" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3467" />
                    <RANKING order="2" place="2" resultid="2227" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1209" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3514" />
                    <RANKING order="2" place="2" resultid="3846" />
                    <RANKING order="3" place="3" resultid="2670" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1210" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2200" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1211" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2581" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1212" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2620" />
                    <RANKING order="2" place="2" resultid="3025" />
                    <RANKING order="3" place="3" resultid="2398" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4709" daytime="11:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4710" daytime="11:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4711" daytime="11:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4712" daytime="11:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4713" daytime="11:45" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1213" daytime="11:50" gender="F" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1214" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2554" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1215" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29" />
                <AGEGROUP agegroupid="1216" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3300" />
                    <RANKING order="2" place="2" resultid="3650" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1217" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2830" />
                    <RANKING order="2" place="2" resultid="3019" />
                    <RANKING order="3" place="3" resultid="2222" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1218" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2641" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1219" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3647" />
                    <RANKING order="2" place="2" resultid="3363" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1220" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54" />
                <AGEGROUP agegroupid="1221" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2700" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1222" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2636" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1223" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2311" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1224" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74" />
                <AGEGROUP agegroupid="1225" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="1226" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4714" daytime="11:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4715" daytime="11:55" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1227" daytime="12:00" gender="M" number="10" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1228" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2550" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1229" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3251" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1230" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3240" />
                    <RANKING order="2" place="2" resultid="2418" />
                    <RANKING order="3" place="-1" resultid="3574" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1231" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2238" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1232" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2858" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1233" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3295" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1234" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2649" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1235" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59" />
                <AGEGROUP agegroupid="1236" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64" />
                <AGEGROUP agegroupid="1237" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3485" />
                    <RANKING order="2" place="2" resultid="3557" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1238" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74" />
                <AGEGROUP agegroupid="1239" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="1240" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4716" daytime="12:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4717" daytime="12:05" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1241" daytime="12:10" gender="F" number="11" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1242" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24" />
                <AGEGROUP agegroupid="1243" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3109" />
                    <RANKING order="2" place="2" resultid="2327" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1244" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34" />
                <AGEGROUP agegroupid="1245" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39" />
                <AGEGROUP agegroupid="1246" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2478" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1247" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3660" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1248" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3417" />
                    <RANKING order="2" place="-1" resultid="2601" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1249" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59" />
                <AGEGROUP agegroupid="1250" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2596" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1251" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69" />
                <AGEGROUP agegroupid="1252" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74" />
                <AGEGROUP agegroupid="1253" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3533" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1254" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4718" daytime="12:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4719" daytime="12:10" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1255" daytime="12:15" gender="M" number="12" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1256" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2899" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1257" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2794" />
                    <RANKING order="2" place="2" resultid="3089" />
                    <RANKING order="3" place="3" resultid="2169" />
                    <RANKING order="4" place="-1" resultid="3246" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1258" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3069" />
                    <RANKING order="2" place="2" resultid="2820" />
                    <RANKING order="3" place="3" resultid="2351" />
                    <RANKING order="4" place="4" resultid="3626" />
                    <RANKING order="5" place="5" resultid="2879" />
                    <RANKING order="6" place="6" resultid="3291" />
                    <RANKING order="7" place="-1" resultid="3094" />
                    <RANKING order="8" place="-1" resultid="3597" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1259" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3832" />
                    <RANKING order="2" place="2" resultid="2431" />
                    <RANKING order="3" place="3" resultid="2426" />
                    <RANKING order="4" place="-1" resultid="3579" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1260" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2472" />
                    <RANKING order="2" place="2" resultid="3315" />
                    <RANKING order="3" place="-1" resultid="3143" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1261" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2333" />
                    <RANKING order="2" place="2" resultid="2530" />
                    <RANKING order="3" place="-1" resultid="2840" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1262" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3233" />
                    <RANKING order="2" place="2" resultid="2675" />
                    <RANKING order="3" place="3" resultid="2483" />
                    <RANKING order="4" place="4" resultid="3059" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1263" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2210" />
                    <RANKING order="2" place="-1" resultid="3457" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1264" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3273" />
                    <RANKING order="2" place="2" resultid="3172" />
                    <RANKING order="3" place="3" resultid="2575" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1265" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3396" />
                    <RANKING order="2" place="2" resultid="2394" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1266" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74" />
                <AGEGROUP agegroupid="1267" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="1268" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4720" daytime="12:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4721" daytime="12:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4722" daytime="12:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4723" daytime="12:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4724" daytime="12:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4725" daytime="12:25" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1269" daytime="12:30" gender="F" number="13" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1270" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2320" />
                    <RANKING order="2" place="2" resultid="3176" />
                    <RANKING order="3" place="3" resultid="2555" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1271" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2835" />
                    <RANKING order="2" place="2" resultid="3256" />
                    <RANKING order="3" place="-1" resultid="3653" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1272" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3301" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1273" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2802" />
                    <RANKING order="2" place="2" resultid="2915" />
                    <RANKING order="3" place="3" resultid="3186" />
                    <RANKING order="4" place="4" resultid="2626" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1274" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3602" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1275" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3369" />
                    <RANKING order="2" place="2" resultid="3364" />
                    <RANKING order="3" place="3" resultid="3335" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1276" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3033" />
                    <RANKING order="2" place="-1" resultid="3191" />
                    <RANKING order="3" place="-1" resultid="3540" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1277" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59" />
                <AGEGROUP agegroupid="1278" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3202" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1279" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69" />
                <AGEGROUP agegroupid="1280" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1281" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="1282" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi" />
                <AGEGROUP agegroupid="4822" agemax="-1" agemin="20" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2835" />
                    <RANKING order="2" place="2" resultid="3256" />
                    <RANKING order="3" place="3" resultid="2320" />
                    <RANKING order="4" place="4" resultid="3176" />
                    <RANKING order="5" place="5" resultid="3033" />
                    <RANKING order="6" place="6" resultid="2802" />
                    <RANKING order="7" place="7" resultid="3602" />
                    <RANKING order="8" place="8" resultid="2555" />
                    <RANKING order="9" place="9" resultid="3301" />
                    <RANKING order="10" place="10" resultid="3369" />
                    <RANKING order="11" place="11" resultid="3364" />
                    <RANKING order="12" place="12" resultid="3202" />
                    <RANKING order="13" place="13" resultid="2915" />
                    <RANKING order="14" place="14" resultid="3186" />
                    <RANKING order="15" place="15" resultid="3335" />
                    <RANKING order="16" place="16" resultid="2626" />
                    <RANKING order="17" place="17" resultid="3524" />
                    <RANKING order="18" place="-1" resultid="3191" />
                    <RANKING order="19" place="-1" resultid="3540" />
                    <RANKING order="20" place="-1" resultid="3653" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4726" daytime="12:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4727" daytime="12:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4728" daytime="12:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4729" daytime="12:45" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1283" daytime="12:50" gender="M" number="14" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1284" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3611" />
                    <RANKING order="2" place="2" resultid="3850" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1285" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3264" />
                    <RANKING order="2" place="2" resultid="2845" />
                    <RANKING order="3" place="3" resultid="2894" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1286" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3425" />
                    <RANKING order="2" place="2" resultid="3241" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1287" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3569" />
                    <RANKING order="2" place="2" resultid="3475" />
                    <RANKING order="3" place="3" resultid="2460" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1288" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44" />
                <AGEGROUP agegroupid="1289" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3480" />
                    <RANKING order="2" place="2" resultid="2711" />
                    <RANKING order="3" place="3" resultid="3279" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1290" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2363" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1291" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2863" />
                    <RANKING order="2" place="2" resultid="3038" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1292" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3168" />
                    <RANKING order="2" place="2" resultid="3325" />
                    <RANKING order="3" place="3" resultid="2576" />
                    <RANKING order="4" place="4" resultid="3635" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1293" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3391" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1294" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4820" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1295" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="1296" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3530" />
                    <RANKING order="2" place="2" resultid="2454" />
                    <RANKING order="3" place="3" resultid="2621" />
                    <RANKING order="4" place="4" resultid="3026" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4823" agemax="-1" agemin="20" name="OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3264" />
                    <RANKING order="2" place="2" resultid="3611" />
                    <RANKING order="3" place="3" resultid="2845" />
                    <RANKING order="4" place="4" resultid="3425" />
                    <RANKING order="5" place="5" resultid="2363" />
                    <RANKING order="6" place="6" resultid="3569" />
                    <RANKING order="7" place="7" resultid="3850" />
                    <RANKING order="8" place="8" resultid="3475" />
                    <RANKING order="9" place="9" resultid="3241" />
                    <RANKING order="10" place="10" resultid="3480" />
                    <RANKING order="11" place="11" resultid="2711" />
                    <RANKING order="12" place="12" resultid="2894" />
                    <RANKING order="13" place="13" resultid="3279" />
                    <RANKING order="14" place="14" resultid="2863" />
                    <RANKING order="15" place="15" resultid="3168" />
                    <RANKING order="16" place="16" resultid="3325" />
                    <RANKING order="17" place="17" resultid="3391" />
                    <RANKING order="18" place="18" resultid="2576" />
                    <RANKING order="19" place="19" resultid="3038" />
                    <RANKING order="20" place="20" resultid="3635" />
                    <RANKING order="21" place="21" resultid="3530" />
                    <RANKING order="22" place="22" resultid="2460" />
                    <RANKING order="23" place="23" resultid="2454" />
                    <RANKING order="24" place="24" resultid="4820" />
                    <RANKING order="25" place="25" resultid="2621" />
                    <RANKING order="26" place="26" resultid="3026" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4730" daytime="12:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4731" daytime="12:55" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4732" daytime="13:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4733" daytime="13:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4734" daytime="13:10" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1088" daytime="13:15" gender="F" number="15" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1089" agemax="96" agemin="80" name="Kategoria &quot;0&quot; 80-96" />
                <AGEGROUP agegroupid="1090" agemax="119" agemin="100" name="Kategoria &quot;A&quot; 100-119" />
                <AGEGROUP agegroupid="1331" agemax="159" agemin="120" name="Kategoria &quot;B&quot; 120-159" />
                <AGEGROUP agegroupid="1332" agemax="199" agemin="160" name="Kategoria &quot;C&quot; 160-199">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3662" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1333" agemax="239" agemin="200" name="Kategoria &quot;D&quot; 200-239" />
                <AGEGROUP agegroupid="1334" agemax="279" agemin="240" name="Kategoria &quot;E&quot; 240-279" />
                <AGEGROUP agegroupid="1335" agemax="-1" agemin="280" name="Kategoria &quot;F&quot; 280 +" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4735" daytime="13:15" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1325" daytime="13:20" gender="M" number="16" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1336" agemax="96" agemin="80" name="Kategoria &quot;0&quot; 80-96" />
                <AGEGROUP agegroupid="1337" agemax="119" agemin="100" name="Kategoria &quot;A&quot; 100-119">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3120" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1338" agemax="159" agemin="120" name="Kategoria &quot;B&quot; 120-159">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4811" />
                    <RANKING order="2" place="2" resultid="2439" />
                    <RANKING order="3" place="3" resultid="2902" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1339" agemax="199" agemin="160" name="Kategoria &quot;C&quot; 160-199">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3548" />
                    <RANKING order="2" place="2" resultid="3342" />
                    <RANKING order="3" place="3" resultid="2681" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1340" agemax="239" agemin="200" name="Kategoria &quot;D&quot; 200-239">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3442" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1341" agemax="279" agemin="240" name="Kategoria &quot;E&quot; 240-279" />
                <AGEGROUP agegroupid="1342" agemax="-1" agemin="280" name="Kategoria &quot;F&quot; 280 +" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4736" daytime="13:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4737" daytime="13:25" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2022-05-14" daytime="16:00" endtime="19:51" number="2" warmupfrom="15:00" warmupuntil="15:50">
          <EVENTS>
            <EVENT eventid="1329" daytime="16:00" gender="F" number="17" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1343" agemax="96" agemin="80" name="Kategoria &quot;0&quot; 80-96" />
                <AGEGROUP agegroupid="1344" agemax="119" agemin="100" name="Kategoria &quot;A&quot; 100-119" />
                <AGEGROUP agegroupid="1345" agemax="159" agemin="120" name="Kategoria &quot;B&quot; 120-159">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3663" />
                    <RANKING order="2" place="-1" resultid="2867" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1346" agemax="199" agemin="160" name="Kategoria &quot;C&quot; 160-199">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2678" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1347" agemax="239" agemin="200" name="Kategoria &quot;D&quot; 200-239">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3440" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1348" agemax="279" agemin="240" name="Kategoria &quot;E&quot; 240-279">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3224" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1349" agemax="-1" agemin="280" name="Kategoria &quot;F&quot; 280 +" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4738" daytime="16:00" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1350" daytime="16:05" gender="M" number="18" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1351" agemax="96" agemin="80" name="Kategoria &quot;0&quot; 80-96" />
                <AGEGROUP agegroupid="1352" agemax="119" agemin="100" name="Kategoria &quot;A&quot; 100-119">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3121" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1353" agemax="159" agemin="120" name="Kategoria &quot;B&quot; 120-159">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2866" />
                    <RANKING order="2" place="2" resultid="4812" />
                    <RANKING order="3" place="3" resultid="2438" />
                    <RANKING order="4" place="4" resultid="2903" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1354" agemax="199" agemin="160" name="Kategoria &quot;C&quot; 160-199">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3343" />
                    <RANKING order="2" place="-1" resultid="3223" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1355" agemax="239" agemin="200" name="Kategoria &quot;D&quot; 200-239">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2679" />
                    <RANKING order="2" place="2" resultid="3441" />
                    <RANKING order="3" place="-1" resultid="3491" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1356" agemax="279" agemin="240" name="Kategoria &quot;E&quot; 240-279">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2680" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1357" agemax="-1" agemin="280" name="Kategoria &quot;F&quot; 280 +">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3543" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4739" daytime="16:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4740" daytime="16:10" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1358" daytime="16:15" gender="F" number="19" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1366" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24" />
                <AGEGROUP agegroupid="1367" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3054" />
                    <RANKING order="2" place="2" resultid="2328" />
                    <RANKING order="3" place="3" resultid="2245" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1368" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3269" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1369" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="2850" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1370" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2536" />
                    <RANKING order="2" place="2" resultid="3643" />
                    <RANKING order="3" place="3" resultid="3603" />
                    <RANKING order="4" place="4" resultid="2642" />
                    <RANKING order="5" place="5" resultid="3182" />
                    <RANKING order="6" place="6" resultid="2479" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1371" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3649" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1372" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3418" />
                    <RANKING order="2" place="2" resultid="2158" />
                    <RANKING order="3" place="-1" resultid="2602" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1373" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2572" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1374" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3374" />
                    <RANKING order="2" place="2" resultid="2637" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1375" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69" />
                <AGEGROUP agegroupid="1376" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74" />
                <AGEGROUP agegroupid="1377" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="1378" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4741" daytime="16:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4742" daytime="16:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4743" daytime="16:15" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1379" daytime="16:20" gender="M" number="20" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1380" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3080" />
                    <RANKING order="2" place="2" resultid="3160" />
                    <RANKING order="3" place="3" resultid="2188" />
                    <RANKING order="4" place="4" resultid="2900" />
                    <RANKING order="5" place="5" resultid="2813" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1381" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2795" />
                    <RANKING order="2" place="2" resultid="3247" />
                    <RANKING order="3" place="3" resultid="3090" />
                    <RANKING order="4" place="4" resultid="2170" />
                    <RANKING order="5" place="5" resultid="3252" />
                    <RANKING order="6" place="6" resultid="2617" />
                    <RANKING order="7" place="-1" resultid="2316" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1382" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3070" />
                    <RANKING order="2" place="2" resultid="2880" />
                    <RANKING order="3" place="3" resultid="2885" />
                    <RANKING order="4" place="4" resultid="2419" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1383" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3830" />
                    <RANKING order="2" place="2" resultid="2432" />
                    <RANKING order="3" place="3" resultid="2239" />
                    <RANKING order="4" place="4" resultid="3077" />
                    <RANKING order="5" place="5" resultid="2890" />
                    <RANKING order="6" place="-1" resultid="2165" />
                    <RANKING order="7" place="-1" resultid="3580" />
                    <RANKING order="8" place="-1" resultid="3668" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1384" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3144" />
                    <RANKING order="2" place="-1" resultid="3135" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1385" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2841" />
                    <RANKING order="2" place="2" resultid="2334" />
                    <RANKING order="3" place="3" resultid="3139" />
                    <RANKING order="4" place="4" resultid="2826" />
                    <RANKING order="5" place="5" resultid="2531" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1386" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2607" />
                    <RANKING order="2" place="2" resultid="3434" />
                    <RANKING order="3" place="3" resultid="2484" />
                    <RANKING order="4" place="4" resultid="3360" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1387" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3458" />
                    <RANKING order="2" place="2" resultid="2211" />
                    <RANKING order="3" place="3" resultid="3206" />
                    <RANKING order="4" place="3" resultid="3504" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1388" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2587" />
                    <RANKING order="2" place="2" resultid="3173" />
                    <RANKING order="3" place="3" resultid="3636" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1389" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3397" />
                    <RANKING order="2" place="2" resultid="2395" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1390" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3528" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1391" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2176" />
                    <RANKING order="2" place="2" resultid="3510" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1392" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4744" daytime="16:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4745" daytime="16:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4746" daytime="16:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4747" daytime="16:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4748" daytime="16:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4749" daytime="16:25" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4750" daytime="16:25" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4751" daytime="16:25" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1393" daytime="16:30" gender="F" number="21" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1394" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3608" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1395" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3110" />
                    <RANKING order="2" place="2" resultid="2921" />
                    <RANKING order="3" place="3" resultid="3055" />
                    <RANKING order="4" place="4" resultid="2329" />
                    <RANKING order="5" place="5" resultid="3115" />
                    <RANKING order="6" place="6" resultid="2244" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1396" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2716" />
                    <RANKING order="2" place="2" resultid="3198" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1397" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2414" />
                    <RANKING order="2" place="2" resultid="3285" />
                    <RANKING order="3" place="3" resultid="2223" />
                    <RANKING order="4" place="4" resultid="3828" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1398" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2206" />
                    <RANKING order="2" place="2" resultid="3644" />
                    <RANKING order="3" place="3" resultid="2632" />
                    <RANKING order="4" place="4" resultid="3183" />
                    <RANKING order="5" place="-1" resultid="3586" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1399" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3661" />
                    <RANKING order="2" place="2" resultid="3422" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1400" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3541" />
                    <RANKING order="2" place="2" resultid="3379" />
                    <RANKING order="3" place="3" resultid="2159" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1401" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3152" />
                    <RANKING order="2" place="2" resultid="3331" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1402" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2597" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1403" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2312" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1404" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3553" />
                    <RANKING order="2" place="2" resultid="3520" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1405" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="1406" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3195" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4752" daytime="16:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4753" daytime="16:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4754" daytime="16:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4755" daytime="16:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4756" daytime="16:40" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1407" daytime="16:40" gender="M" number="22" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1408" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3081" />
                    <RANKING order="2" place="2" resultid="3161" />
                    <RANKING order="3" place="3" resultid="2378" />
                    <RANKING order="4" place="4" resultid="3165" />
                    <RANKING order="5" place="5" resultid="2901" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1409" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3091" />
                    <RANKING order="2" place="2" resultid="3105" />
                    <RANKING order="3" place="3" resultid="3622" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1410" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3071" />
                    <RANKING order="2" place="2" resultid="2352" />
                    <RANKING order="3" place="3" resultid="3321" />
                    <RANKING order="4" place="-1" resultid="2881" />
                    <RANKING order="5" place="-1" resultid="3598" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1411" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3669" />
                    <RANKING order="2" place="2" resultid="2346" />
                    <RANKING order="3" place="3" resultid="2427" />
                    <RANKING order="4" place="-1" resultid="2163" />
                    <RANKING order="5" place="-1" resultid="3476" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1412" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2816" />
                    <RANKING order="2" place="2" resultid="3618" />
                    <RANKING order="3" place="3" resultid="2195" />
                    <RANKING order="4" place="4" resultid="2374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1413" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3500" />
                    <RANKING order="2" place="2" resultid="2827" />
                    <RANKING order="3" place="3" resultid="3400" />
                    <RANKING order="4" place="4" resultid="2566" />
                    <RANKING order="5" place="5" resultid="3296" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1414" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3361" />
                    <RANKING order="2" place="2" resultid="3563" />
                    <RANKING order="3" place="3" resultid="3646" />
                    <RANKING order="4" place="4" resultid="3060" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1415" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3505" />
                    <RANKING order="2" place="2" resultid="2592" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1416" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3468" />
                    <RANKING order="2" place="2" resultid="3405" />
                    <RANKING order="3" place="3" resultid="2228" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1417" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3515" />
                    <RANKING order="2" place="2" resultid="3847" />
                    <RANKING order="3" place="3" resultid="2671" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1418" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2201" />
                    <RANKING order="2" place="2" resultid="3356" />
                    <RANKING order="3" place="-1" resultid="3228" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1419" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2582" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1420" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4757" daytime="16:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4758" daytime="16:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4759" daytime="16:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4760" daytime="16:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4761" daytime="16:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4762" daytime="16:55" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4763" daytime="16:55" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4764" daytime="16:55" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1575" daytime="17:00" gender="F" number="23" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1576" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2322" />
                    <RANKING order="2" place="2" resultid="3177" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1577" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2836" />
                    <RANKING order="2" place="2" resultid="3257" />
                    <RANKING order="3" place="-1" resultid="3654" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1578" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3302" />
                    <RANKING order="2" place="2" resultid="3651" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1579" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2854" />
                    <RANKING order="2" place="2" resultid="2803" />
                    <RANKING order="3" place="3" resultid="3657" />
                    <RANKING order="4" place="4" resultid="3187" />
                    <RANKING order="5" place="5" resultid="2627" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1580" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2541" />
                    <RANKING order="2" place="2" resultid="2546" />
                    <RANKING order="3" place="3" resultid="3415" />
                    <RANKING order="4" place="-1" resultid="3604" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1581" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3370" />
                    <RANKING order="2" place="2" resultid="3336" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1582" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3034" />
                    <RANKING order="2" place="2" resultid="3854" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1583" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2339" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1584" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3203" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1585" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69" />
                <AGEGROUP agegroupid="1586" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3525" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1587" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3534" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1588" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4765" daytime="17:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4766" daytime="17:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4767" daytime="17:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4768" daytime="17:10" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1589" daytime="17:10" gender="M" number="24" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1590" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2561" />
                    <RANKING order="2" place="2" resultid="3612" />
                    <RANKING order="3" place="3" resultid="2369" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1591" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3265" />
                    <RANKING order="2" place="2" resultid="2846" />
                    <RANKING order="3" place="3" resultid="3430" />
                    <RANKING order="4" place="4" resultid="2895" />
                    <RANKING order="5" place="5" resultid="2618" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1592" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3426" />
                    <RANKING order="2" place="2" resultid="3627" />
                    <RANKING order="3" place="3" resultid="3242" />
                    <RANKING order="4" place="4" resultid="2420" />
                    <RANKING order="5" place="-1" resultid="2821" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1593" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3570" />
                    <RANKING order="2" place="2" resultid="2240" />
                    <RANKING order="3" place="3" resultid="2461" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1594" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3311" />
                    <RANKING order="2" place="2" resultid="3472" />
                    <RANKING order="3" place="3" resultid="3438" />
                    <RANKING order="4" place="4" resultid="3410" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1595" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3489" />
                    <RANKING order="2" place="2" resultid="3481" />
                    <RANKING order="3" place="3" resultid="3280" />
                    <RANKING order="4" place="4" resultid="2217" />
                    <RANKING order="5" place="-1" resultid="3384" />
                    <RANKING order="6" place="-1" resultid="3463" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1596" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2364" />
                    <RANKING order="2" place="2" resultid="2676" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1597" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2864" />
                    <RANKING order="2" place="2" resultid="3043" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1598" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3169" />
                    <RANKING order="2" place="2" resultid="3326" />
                    <RANKING order="3" place="3" resultid="2577" />
                    <RANKING order="4" place="-1" resultid="3637" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1599" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3392" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1600" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74" />
                <AGEGROUP agegroupid="1601" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2410" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1602" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3531" />
                    <RANKING order="2" place="2" resultid="2455" />
                    <RANKING order="3" place="3" resultid="2622" />
                    <RANKING order="4" place="4" resultid="3028" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4769" daytime="17:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4770" daytime="17:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4771" daytime="17:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4772" daytime="17:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4773" daytime="17:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4774" daytime="17:25" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4775" daytime="17:25" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1421" daytime="17:30" gender="F" number="25" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1422" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3208" />
                    <RANKING order="2" place="2" resultid="2556" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1423" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29" />
                <AGEGROUP agegroupid="1424" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34" />
                <AGEGROUP agegroupid="1425" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2809" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1426" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3587" />
                    <RANKING order="2" place="-1" resultid="3841" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1427" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49" />
                <AGEGROUP agegroupid="1428" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54" />
                <AGEGROUP agegroupid="1429" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3332" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1430" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64" />
                <AGEGROUP agegroupid="1431" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69" />
                <AGEGROUP agegroupid="1432" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74" />
                <AGEGROUP agegroupid="1433" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="1434" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4776" daytime="17:30" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1435" daytime="17:35" gender="M" number="26" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1436" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2551" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1437" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3248" />
                    <RANKING order="2" place="2" resultid="3100" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1438" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3095" />
                    <RANKING order="2" place="2" resultid="2467" />
                    <RANKING order="3" place="-1" resultid="3575" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1439" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39" />
                <AGEGROUP agegroupid="1440" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2473" />
                    <RANKING order="2" place="2" resultid="2859" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1441" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3340" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1442" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3234" />
                    <RANKING order="2" place="2" resultid="2182" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1443" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3048" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1444" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3274" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1445" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3486" />
                    <RANKING order="2" place="2" resultid="3558" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1446" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3506" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1447" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="1448" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2391" />
                    <RANKING order="2" place="2" resultid="2399" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4777" daytime="17:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4778" daytime="17:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4779" daytime="17:45" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1449" daytime="17:50" gender="F" number="27" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1450" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24" />
                <AGEGROUP agegroupid="1451" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29" />
                <AGEGROUP agegroupid="1452" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34" />
                <AGEGROUP agegroupid="1453" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39" />
                <AGEGROUP agegroupid="1454" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2480" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1455" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3365" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1456" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54" />
                <AGEGROUP agegroupid="1457" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59" />
                <AGEGROUP agegroupid="1458" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2598" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1459" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69" />
                <AGEGROUP agegroupid="1460" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74" />
                <AGEGROUP agegroupid="1461" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="1462" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4780" daytime="17:50" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1463" daytime="17:55" gender="M" number="28" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1464" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3613" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1465" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29" />
                <AGEGROUP agegroupid="1466" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3628" />
                    <RANKING order="2" place="2" resultid="4824" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1467" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3477" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1468" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3316" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1469" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2712" />
                    <RANKING order="2" place="-1" resultid="3482" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1470" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2485" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1471" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3039" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1472" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2578" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1473" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69" />
                <AGEGROUP agegroupid="1474" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74" />
                <AGEGROUP agegroupid="1475" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="1476" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4781" daytime="17:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4782" daytime="18:00" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1477" daytime="18:05" gender="F" number="29" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1478" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3178" />
                    <RANKING order="2" place="2" resultid="2557" />
                    <RANKING order="3" place="3" resultid="2323" />
                    <RANKING order="4" place="4" resultid="3216" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1479" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3111" />
                    <RANKING order="2" place="2" resultid="2922" />
                    <RANKING order="3" place="3" resultid="2837" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1480" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3303" />
                    <RANKING order="2" place="2" resultid="3065" />
                    <RANKING order="3" place="3" resultid="3652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1481" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2831" />
                    <RANKING order="2" place="2" resultid="2855" />
                    <RANKING order="3" place="3" resultid="2804" />
                    <RANKING order="4" place="4" resultid="3020" />
                    <RANKING order="5" place="5" resultid="2224" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1482" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2643" />
                    <RANKING order="2" place="2" resultid="2542" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1483" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3648" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1484" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54" />
                <AGEGROUP agegroupid="1485" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2573" />
                    <RANKING order="2" place="2" resultid="2340" />
                    <RANKING order="3" place="3" resultid="2701" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1486" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3375" />
                    <RANKING order="2" place="2" resultid="2638" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1487" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69" />
                <AGEGROUP agegroupid="1488" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74" />
                <AGEGROUP agegroupid="1489" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79" />
                <AGEGROUP agegroupid="1490" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4783" daytime="18:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4784" daytime="18:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4785" daytime="18:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4786" daytime="18:10" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1491" daytime="18:15" gender="M" number="30" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1492" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2562" />
                    <RANKING order="2" place="2" resultid="2370" />
                    <RANKING order="3" place="3" resultid="2189" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1493" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2796" />
                    <RANKING order="2" place="2" resultid="3253" />
                    <RANKING order="3" place="3" resultid="2171" />
                    <RANKING order="4" place="4" resultid="3431" />
                    <RANKING order="5" place="5" resultid="3106" />
                    <RANKING order="6" place="6" resultid="2896" />
                    <RANKING order="7" place="-1" resultid="2317" />
                    <RANKING order="8" place="-1" resultid="2437" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1494" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2822" />
                    <RANKING order="2" place="2" resultid="3322" />
                    <RANKING order="3" place="3" resultid="2612" />
                    <RANKING order="4" place="4" resultid="3631" />
                    <RANKING order="5" place="-1" resultid="2423" />
                    <RANKING order="6" place="-1" resultid="2886" />
                    <RANKING order="7" place="-1" resultid="3576" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1495" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2891" />
                    <RANKING order="2" place="2" resultid="2428" />
                    <RANKING order="3" place="3" resultid="2462" />
                    <RANKING order="4" place="-1" resultid="2433" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1496" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2860" />
                    <RANKING order="2" place="2" resultid="3411" />
                    <RANKING order="3" place="3" resultid="2196" />
                    <RANKING order="4" place="4" resultid="2658" />
                    <RANKING order="5" place="-1" resultid="3136" />
                    <RANKING order="6" place="-1" resultid="3145" />
                    <RANKING order="7" place="-1" resultid="3312" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1497" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2335" />
                    <RANKING order="2" place="2" resultid="3281" />
                    <RANKING order="3" place="3" resultid="2532" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1498" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2365" />
                    <RANKING order="2" place="2" resultid="2608" />
                    <RANKING order="3" place="3" resultid="2650" />
                    <RANKING order="4" place="4" resultid="3435" />
                    <RANKING order="5" place="5" resultid="3564" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1499" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3459" />
                    <RANKING order="2" place="2" resultid="2212" />
                    <RANKING order="3" place="3" resultid="2593" />
                    <RANKING order="4" place="4" resultid="3044" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1500" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3327" />
                    <RANKING order="2" place="2" resultid="3406" />
                    <RANKING order="3" place="-1" resultid="3469" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1501" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3393" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1502" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3229" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1503" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2177" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1504" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2456" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4787" daytime="18:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4788" daytime="18:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4789" daytime="18:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4790" daytime="18:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4791" daytime="18:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4792" daytime="18:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4793" daytime="18:30" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4794" daytime="18:30" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1505" daytime="18:35" gender="F" number="31" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1506" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3213" />
                    <RANKING order="2" place="2" resultid="3217" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1507" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3180" />
                    <RANKING order="2" place="2" resultid="3261" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1508" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3270" />
                    <RANKING order="2" place="2" resultid="3066" />
                    <RANKING order="3" place="-1" resultid="3199" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1509" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2832" />
                    <RANKING order="2" place="2" resultid="3827" />
                    <RANKING order="3" place="3" resultid="2628" />
                    <RANKING order="4" place="4" resultid="3188" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1510" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2537" />
                    <RANKING order="2" place="2" resultid="2633" />
                    <RANKING order="3" place="3" resultid="2547" />
                    <RANKING order="4" place="-1" resultid="3842" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1511" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49" />
                <AGEGROUP agegroupid="1512" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3380" />
                    <RANKING order="2" place="-1" resultid="2603" />
                    <RANKING order="3" place="-1" resultid="3853" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1513" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3153" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1514" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64" />
                <AGEGROUP agegroupid="1515" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69" />
                <AGEGROUP agegroupid="1516" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3554" />
                    <RANKING order="2" place="2" resultid="3521" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1517" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2403" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1518" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3196" />
                    <RANKING order="2" place="2" resultid="3838" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4795" daytime="18:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4796" daytime="18:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4797" daytime="18:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4798" daytime="18:40" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1519" daytime="18:45" gender="M" number="32" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1520" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2552" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1521" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3101" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1522" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3096" />
                    <RANKING order="2" place="2" resultid="2468" />
                    <RANKING order="3" place="3" resultid="2613" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1523" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3831" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1524" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2474" />
                    <RANKING order="2" place="2" resultid="3439" />
                    <RANKING order="3" place="3" resultid="2659" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1525" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2842" />
                    <RANKING order="2" place="2" resultid="3341" />
                    <RANKING order="3" place="3" resultid="2218" />
                    <RANKING order="4" place="4" resultid="2567" />
                    <RANKING order="5" place="-1" resultid="3140" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1526" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2677" />
                    <RANKING order="2" place="2" resultid="2662" />
                    <RANKING order="3" place="3" resultid="2183" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1527" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3049" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1528" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3275" />
                    <RANKING order="2" place="2" resultid="2588" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1529" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3398" />
                    <RANKING order="2" place="2" resultid="2396" />
                    <RANKING order="3" place="3" resultid="3848" />
                    <RANKING order="4" place="4" resultid="2672" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1530" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3537" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1531" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3511" />
                    <RANKING order="2" place="2" resultid="2408" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1532" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2392" />
                    <RANKING order="2" place="2" resultid="2400" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4799" daytime="18:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4800" daytime="18:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4801" daytime="18:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4802" daytime="18:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4803" daytime="18:50" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1533" daytime="18:50" gender="F" number="33" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1534" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3209" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1535" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3116" />
                    <RANKING order="2" place="2" resultid="3655" />
                    <RANKING order="3" place="-1" resultid="3258" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1536" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34" />
                <AGEGROUP agegroupid="1537" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2810" />
                    <RANKING order="2" place="2" resultid="3021" />
                    <RANKING order="3" place="3" resultid="3286" />
                    <RANKING order="4" place="4" resultid="2415" />
                    <RANKING order="5" place="5" resultid="3658" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1538" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2207" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1539" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3366" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1540" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3542" />
                    <RANKING order="2" place="2" resultid="3035" />
                    <RANKING order="3" place="-1" resultid="3192" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1541" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2702" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1542" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64" />
                <AGEGROUP agegroupid="1543" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2313" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1544" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74" />
                <AGEGROUP agegroupid="1545" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2404" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1546" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi" />
                <AGEGROUP agegroupid="4813" agemax="-1" agemin="20" name="Kategoria OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2207" />
                    <RANKING order="2" place="2" resultid="3116" />
                    <RANKING order="3" place="3" resultid="3542" />
                    <RANKING order="4" place="4" resultid="3209" />
                    <RANKING order="5" place="5" resultid="2810" />
                    <RANKING order="6" place="6" resultid="3035" />
                    <RANKING order="7" place="7" resultid="3021" />
                    <RANKING order="8" place="8" resultid="3286" />
                    <RANKING order="9" place="9" resultid="2415" />
                    <RANKING order="10" place="10" resultid="2702" />
                    <RANKING order="11" place="11" resultid="3366" />
                    <RANKING order="12" place="12" resultid="3658" />
                    <RANKING order="13" place="13" resultid="3655" />
                    <RANKING order="14" place="14" resultid="2313" />
                    <RANKING order="15" place="15" resultid="2404" />
                    <RANKING order="16" place="-1" resultid="3192" />
                    <RANKING order="17" place="-1" resultid="3258" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4804" daytime="18:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4805" daytime="19:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4806" daytime="19:05" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1547" daytime="19:15" gender="M" number="34" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1548" agemax="24" agemin="20" name="Kategoria &quot;0&quot; 20-24">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2379" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1549" agemax="29" agemin="25" name="Kategoria &quot;A&quot; 25-29">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2847" />
                    <RANKING order="2" place="2" resultid="3623" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1550" agemax="34" agemin="30" name="Kategoria &quot;B&quot; 30-34">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2353" />
                    <RANKING order="2" place="2" resultid="3293" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1551" agemax="39" agemin="35" name="Kategoria &quot;C&quot; 35-39">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1552" agemax="44" agemin="40" name="Kategoria &quot;D&quot; 40-44">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3317" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1553" agemax="49" agemin="45" name="Kategoria &quot;E&quot; 45-49">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2713" />
                    <RANKING order="2" place="2" resultid="3297" />
                    <RANKING order="3" place="3" resultid="3401" />
                    <RANKING order="4" place="-1" resultid="3385" />
                    <RANKING order="5" place="-1" resultid="3464" />
                    <RANKING order="6" place="-1" resultid="3490" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1554" agemax="54" agemin="50" name="Kategoria &quot;F&quot; 50-54">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3235" />
                    <RANKING order="2" place="2" resultid="3061" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1555" agemax="59" agemin="55" name="Kategoria &quot;G&quot; 55-59">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="2865" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1556" agemax="64" agemin="60" name="Kategoria &quot;H&quot; 60-64">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2229" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1557" agemax="69" agemin="65" name="Kategoria &quot;I&quot; 65-69">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3559" />
                    <RANKING order="2" place="2" resultid="3516" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1558" agemax="74" agemin="70" name="Kategoria &quot;J&quot; 70-74">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2202" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1559" agemax="79" agemin="75" name="Kategoria &quot;K&quot; 75-79">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1560" agemax="-1" agemin="80" name="Kategoria &quot;L&quot; 80 i starsi">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2623" />
                    <RANKING order="2" place="2" resultid="3029" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4814" agemax="-1" agemin="20" name="Kategoria OPEN">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2847" />
                    <RANKING order="2" place="2" resultid="2379" />
                    <RANKING order="3" place="3" resultid="2353" />
                    <RANKING order="4" place="4" resultid="3623" />
                    <RANKING order="5" place="5" resultid="3317" />
                    <RANKING order="6" place="6" resultid="2713" />
                    <RANKING order="7" place="7" resultid="3235" />
                    <RANKING order="8" place="8" resultid="2347" />
                    <RANKING order="9" place="9" resultid="3293" />
                    <RANKING order="10" place="10" resultid="3297" />
                    <RANKING order="11" place="11" resultid="3559" />
                    <RANKING order="12" place="12" resultid="3516" />
                    <RANKING order="13" place="13" resultid="3401" />
                    <RANKING order="14" place="14" resultid="3061" />
                    <RANKING order="15" place="15" resultid="2229" />
                    <RANKING order="16" place="16" resultid="2583" />
                    <RANKING order="17" place="17" resultid="2202" />
                    <RANKING order="18" place="18" resultid="2623" />
                    <RANKING order="19" place="19" resultid="3029" />
                    <RANKING order="20" place="-1" resultid="2865" />
                    <RANKING order="21" place="-1" resultid="3385" />
                    <RANKING order="22" place="-1" resultid="3464" />
                    <RANKING order="23" place="-1" resultid="3490" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4807" daytime="19:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4808" daytime="19:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4809" daytime="19:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4810" daytime="19:40" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="ZILSVK" nation="SVK" clubid="3632" name="PSK Žilina">
          <ATHLETES>
            <ATHLETE firstname="Juraj" lastname="Jaroš" birthdate="1962-06-22" gender="M" nation="SVK" athleteid="3633">
              <RESULTS>
                <RESULT eventid="1171" points="436" swimtime="00:00:41.54" resultid="3634" heatid="4699" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1283" points="330" swimtime="00:03:40.37" resultid="3635" heatid="4731" lane="3" late="yes" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.28" />
                    <SPLIT distance="100" swimtime="00:01:42.47" />
                    <SPLIT distance="150" swimtime="00:02:40.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="398" swimtime="00:00:36.42" resultid="3636" heatid="4746" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1589" status="DNS" swimtime="00:00:00.00" resultid="3637" heatid="4770" lane="3" entrytime="00:01:35.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIEBED" nation="POL" region="11" clubid="2191" name="Zawodnik Niezrzeszony Będzin">
          <ATHLETES>
            <ATHLETE firstname="Robert" lastname="Bomba" birthdate="1978-08-01" gender="M" nation="POL" athleteid="2192">
              <RESULTS>
                <RESULT eventid="1102" points="260" swimtime="00:00:35.65" resultid="2193" heatid="4672" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1171" points="273" swimtime="00:00:43.28" resultid="2194" heatid="4696" lane="3" entrytime="00:00:49.00" />
                <RESULT eventid="1407" points="244" swimtime="00:01:19.49" resultid="2195" heatid="4760" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="188" swimtime="00:01:39.28" resultid="2196" heatid="4789" lane="3" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00611" nation="POL" region="11" clubid="3022" name="AZS AWF Katowice">
          <CONTACT city="Katowice" email="m.skora@awf.katowice.pl" name="Michał Skóra" phone="501370222" state="ŚLĄSK" street="Mikołowska 72a" zip="40-065" />
          <ATHLETES>
            <ATHLETE firstname="Jan" lastname="Ślężyński" birthdate="1931-04-27" gender="M" nation="POL" license="100611700315" athleteid="3023">
              <RESULTS>
                <RESULT eventid="1199" points="143" swimtime="00:06:36.20" resultid="3025" heatid="4709" lane="4" entrytime="00:05:03.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:25.66" />
                    <SPLIT distance="100" swimtime="00:03:11.58" />
                    <SPLIT distance="150" swimtime="00:04:58.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1283" points="178" swimtime="00:07:45.30" resultid="3026" heatid="4731" lane="6" entrytime="00:05:23.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:55.61" />
                    <SPLIT distance="100" swimtime="00:03:53.58" />
                    <SPLIT distance="150" swimtime="00:05:52.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1589" points="158" swimtime="00:03:35.58" resultid="3028" heatid="4769" lane="3" entrytime="00:02:43.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:46.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="135" swimtime="00:15:05.38" resultid="3029" heatid="4807" lane="3" entrytime="00:10:46.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:42.13" />
                    <SPLIT distance="100" swimtime="00:03:37.21" />
                    <SPLIT distance="150" swimtime="00:05:32.83" />
                    <SPLIT distance="200" swimtime="00:07:26.26" />
                    <SPLIT distance="250" swimtime="00:09:19.02" />
                    <SPLIT distance="300" swimtime="00:11:15.20" />
                    <SPLIT distance="350" swimtime="00:13:16.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="RMKRYB" nation="POL" region="11" clubid="3638" name="RMKS Rybnik">
          <ATHLETES>
            <ATHLETE firstname="Anna" lastname="Duda" birthdate="1981-04-15" gender="F" nation="POL" license="101911600104" athleteid="3639">
              <RESULTS>
                <RESULT eventid="1157" points="525" swimtime="00:00:39.87" resultid="3642" heatid="4693" lane="2" entrytime="00:00:40.00" />
                <RESULT eventid="1358" points="713" swimtime="00:00:31.56" resultid="3643" heatid="4743" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="1393" points="621" swimtime="00:01:06.89" resultid="3644" heatid="4755" lane="3" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1059" points="712" swimtime="00:00:29.14" resultid="3822" heatid="4668" lane="3" entrytime="00:00:28.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Henzel" birthdate="1971-09-20" gender="M" nation="POL" license="501911700174" athleteid="3641">
              <RESULTS>
                <RESULT eventid="1102" points="269" swimtime="00:00:36.20" resultid="3645" heatid="4670" lane="6" />
                <RESULT eventid="1407" points="304" swimtime="00:01:16.61" resultid="3646" heatid="4757" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SENRYD" nation="POL" region="11" clubid="2381" name="Rydułtowska Akademia Aktywnego Seniora 60+" shortname="Akademia Aktywnego Seniora 60+">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Lippa" birthdate="1946-02-02" gender="F" nation="POL" athleteid="2385">
              <RESULTS>
                <RESULT eventid="1059" points="60" swimtime="00:01:28.43" resultid="2401" heatid="4664" lane="4" />
                <RESULT eventid="1185" points="92" swimtime="00:06:20.00" resultid="2402" heatid="4705" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.04" />
                    <SPLIT distance="100" swimtime="00:03:03.59" />
                    <SPLIT distance="150" swimtime="00:04:42.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1505" points="66" swimtime="00:01:36.44" resultid="2403" heatid="4795" lane="6" />
                <RESULT eventid="1533" points="101" swimtime="00:13:10.96" resultid="2404" heatid="4804" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:22.88" />
                    <SPLIT distance="100" swimtime="00:03:02.22" />
                    <SPLIT distance="150" swimtime="00:04:43.85" />
                    <SPLIT distance="200" swimtime="00:06:27.83" />
                    <SPLIT distance="250" swimtime="00:08:11.07" />
                    <SPLIT distance="300" swimtime="00:09:50.22" />
                    <SPLIT distance="350" swimtime="00:11:31.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Władysław" lastname="Szurek" birthdate="1940-05-26" gender="M" nation="POL" athleteid="2384">
              <RESULTS>
                <RESULT eventid="1143" points="33" swimtime="00:04:18.55" resultid="2397" heatid="4686" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:57.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1199" points="52" swimtime="00:07:03.71" resultid="2398" heatid="4709" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:27.21" />
                    <SPLIT distance="100" swimtime="00:03:13.16" />
                    <SPLIT distance="150" swimtime="00:05:08.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1435" points="35" swimtime="00:09:35.56" resultid="2399" heatid="4777" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:05.76" />
                    <SPLIT distance="100" swimtime="00:04:33.01" />
                    <SPLIT distance="150" swimtime="00:07:03.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1519" points="28" swimtime="00:02:04.64" resultid="2400" heatid="4799" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rudolf" lastname="Bugla" birthdate="1940-05-16" gender="M" nation="POL" athleteid="2383">
              <RESULTS>
                <RESULT eventid="1143" points="112" swimtime="00:02:52.88" resultid="2386" heatid="4686" lane="4" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="150" swimtime="00:01:17.94" resultid="2390" heatid="4695" lane="4" />
                <RESULT eventid="1435" points="118" swimtime="00:06:21.74" resultid="2391" heatid="4777" lane="4" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:30.61" />
                    <SPLIT distance="100" swimtime="00:03:08.42" />
                    <SPLIT distance="150" swimtime="00:04:45.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1519" points="105" swimtime="00:01:20.06" resultid="2392" heatid="4799" lane="4" entrytime="00:00:59.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Ciecior" birthdate="1953-11-24" gender="M" nation="POL" athleteid="2382">
              <RESULTS>
                <RESULT eventid="1143" points="369" swimtime="00:01:34.35" resultid="2393" heatid="4687" lane="3" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1255" points="228" swimtime="00:01:47.08" resultid="2394" heatid="4721" lane="1" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="364" swimtime="00:00:40.11" resultid="2395" heatid="4744" lane="2" entrytime="00:00:41.00" />
                <RESULT eventid="1519" points="389" swimtime="00:00:41.57" resultid="2396" heatid="4801" lane="1" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="05201" nation="POL" region="01" clubid="2219" name="KS Just Swim Jelenia Góra">
          <CONTACT city="Jelenia Góra" email="marcin.binasiewicz@justswim.pl" name="Binasiewicz Marcin" phone="509071929" state="DOLN" zip="58506" />
          <ATHLETES>
            <ATHLETE firstname="Marek" lastname="Lipka" birthdate="1958-06-05" gender="M" nation="POL" athleteid="2225">
              <RESULTS>
                <RESULT eventid="1102" points="322" swimtime="00:00:36.33" resultid="2226" heatid="4671" lane="3" entrytime="00:00:37.20" />
                <RESULT eventid="1199" points="243" swimtime="00:03:14.93" resultid="2227" heatid="4710" lane="5" entrytime="00:03:10.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.24" />
                    <SPLIT distance="100" swimtime="00:01:31.31" />
                    <SPLIT distance="150" swimtime="00:02:23.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="286" swimtime="00:01:24.77" resultid="2228" heatid="4758" lane="3" entrytime="00:01:20.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="272" swimtime="00:06:56.57" resultid="2229" heatid="4808" lane="2" entrytime="00:06:40.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.66" />
                    <SPLIT distance="100" swimtime="00:01:36.35" />
                    <SPLIT distance="150" swimtime="00:02:28.92" />
                    <SPLIT distance="200" swimtime="00:03:22.30" />
                    <SPLIT distance="250" swimtime="00:04:16.99" />
                    <SPLIT distance="300" swimtime="00:05:11.24" />
                    <SPLIT distance="350" swimtime="00:06:04.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Lara" birthdate="1985-06-16" gender="F" nation="POL" athleteid="2220">
              <RESULTS>
                <RESULT eventid="1185" points="284" swimtime="00:03:07.32" resultid="2221" heatid="4705" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.99" />
                    <SPLIT distance="100" swimtime="00:01:30.95" />
                    <SPLIT distance="150" swimtime="00:02:18.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="265" swimtime="00:03:34.41" resultid="2222" heatid="4714" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.51" />
                    <SPLIT distance="100" swimtime="00:01:50.34" />
                    <SPLIT distance="150" swimtime="00:02:45.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="229" swimtime="00:01:29.87" resultid="2223" heatid="4752" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1477" points="244" swimtime="00:01:41.09" resultid="2224" heatid="4783" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WATWAR" nation="POL" region="14" clubid="2817" name="Water Squad Warszawa">
          <CONTACT city="Warszawa" email="agnieszka.kaczmarek85@gmail.com" name="Kaczmarek" phone="531799855" state="MAZOW" street="Borkow" zip="04-786" />
          <ATHLETES>
            <ATHLETE firstname="Agata" lastname="Korc" birthdate="1986-03-27" gender="F" nation="POL" athleteid="2848">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="2849" heatid="4669" lane="3" entrytime="00:00:26.50" />
                <RESULT eventid="1358" status="DNS" swimtime="00:00:00.00" resultid="2850" heatid="4743" lane="3" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrian" lastname="Kulisz" birthdate="1977-06-16" gender="M" nation="POL" athleteid="2823">
              <RESULTS>
                <RESULT eventid="1102" points="405" swimtime="00:00:30.89" resultid="2824" heatid="4675" lane="1" entrytime="00:00:31.00" />
                <RESULT eventid="1171" points="343" swimtime="00:00:40.93" resultid="2825" heatid="4699" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="1379" points="388" swimtime="00:00:33.44" resultid="2826" heatid="4747" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1407" points="401" swimtime="00:01:07.81" resultid="2827" heatid="4761" lane="5" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Rowinski" birthdate="1990-07-12" gender="M" nation="POL" athleteid="2818">
              <RESULTS>
                <RESULT eventid="1171" points="656" swimtime="00:00:30.75" resultid="2819" heatid="4704" lane="4" entrytime="00:00:29.06" />
                <RESULT eventid="1255" points="591" swimtime="00:01:02.49" resultid="2820" heatid="4724" lane="3" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1589" status="DNS" swimtime="00:00:00.00" resultid="2821" heatid="4775" lane="5" entrytime="00:01:07.50" />
                <RESULT eventid="1491" points="568" swimtime="00:01:04.34" resultid="2822" heatid="4794" lane="2" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Veronica" lastname="Campbell-Żemier" birthdate="1986-04-20" gender="F" nation="POL" athleteid="2851">
              <RESULTS>
                <RESULT eventid="1059" points="652" swimtime="00:00:28.95" resultid="2852" heatid="4664" lane="5" />
                <RESULT eventid="1157" points="639" swimtime="00:00:36.76" resultid="2853" heatid="4691" lane="1" />
                <RESULT eventid="1575" points="595" swimtime="00:01:22.14" resultid="2854" heatid="4765" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1477" points="562" swimtime="00:01:16.56" resultid="2855" heatid="4783" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Kosmider" birthdate="1966-03-01" gender="M" nation="POL" athleteid="2861">
              <RESULTS>
                <RESULT eventid="1102" points="524" swimtime="00:00:30.23" resultid="2862" heatid="4676" lane="3" entrytime="00:00:29.00" />
                <RESULT eventid="1283" points="475" swimtime="00:03:03.11" resultid="2863" heatid="4732" lane="2" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.25" />
                    <SPLIT distance="100" swimtime="00:01:28.69" />
                    <SPLIT distance="150" swimtime="00:02:15.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1589" points="459" swimtime="00:01:23.30" resultid="2864" heatid="4773" lane="2" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" status="DNS" swimtime="00:00:00.00" resultid="2865" heatid="4810" lane="6" entrytime="00:05:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karol" lastname="Żemier" birthdate="1982-11-09" gender="M" nation="POL" athleteid="2856">
              <RESULTS>
                <RESULT eventid="1143" points="638" swimtime="00:01:03.73" resultid="2857" heatid="4686" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="690" swimtime="00:02:21.96" resultid="2858" heatid="4716" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.44" />
                    <SPLIT distance="100" swimtime="00:01:05.84" />
                    <SPLIT distance="150" swimtime="00:01:47.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1435" points="593" swimtime="00:02:27.38" resultid="2859" heatid="4777" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.67" />
                    <SPLIT distance="100" swimtime="00:01:11.31" />
                    <SPLIT distance="150" swimtime="00:01:50.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="684" swimtime="00:01:04.60" resultid="2860" heatid="4787" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Kaczmarek" birthdate="1985-05-07" gender="F" nation="POL" athleteid="2828">
              <RESULTS>
                <RESULT eventid="1129" points="580" swimtime="00:01:12.46" resultid="2829" heatid="4685" lane="5" entrytime="00:01:11.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="579" swimtime="00:02:45.17" resultid="2830" heatid="4715" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.25" />
                    <SPLIT distance="100" swimtime="00:01:17.19" />
                    <SPLIT distance="150" swimtime="00:02:05.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1477" points="626" swimtime="00:01:13.83" resultid="2831" heatid="4786" lane="5" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1505" points="561" swimtime="00:00:33.51" resultid="2832" heatid="4798" lane="4" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arkadiusz" lastname="Aptewicz" birthdate="1993-12-20" gender="M" nation="POL" athleteid="2843">
              <RESULTS>
                <RESULT eventid="1171" points="656" swimtime="00:00:31.07" resultid="2844" heatid="4704" lane="1" entrytime="00:00:30.50" />
                <RESULT eventid="1283" points="656" swimtime="00:02:26.80" resultid="2845" heatid="4734" lane="3" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                    <SPLIT distance="100" swimtime="00:01:10.31" />
                    <SPLIT distance="150" swimtime="00:01:47.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1589" points="600" swimtime="00:01:08.92" resultid="2846" heatid="4775" lane="6" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="753" swimtime="00:04:15.92" resultid="2847" heatid="4810" lane="3" entrytime="00:04:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.59" />
                    <SPLIT distance="100" swimtime="00:01:02.00" />
                    <SPLIT distance="150" swimtime="00:01:34.82" />
                    <SPLIT distance="200" swimtime="00:02:07.91" />
                    <SPLIT distance="250" swimtime="00:02:41.04" />
                    <SPLIT distance="300" swimtime="00:03:13.74" />
                    <SPLIT distance="350" swimtime="00:03:45.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Szyszkowska" birthdate="1996-11-05" gender="F" nation="POL" athleteid="2833">
              <RESULTS>
                <RESULT eventid="1157" points="669" swimtime="00:00:34.87" resultid="2834" heatid="4694" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1269" points="727" swimtime="00:02:44.95" resultid="2835" heatid="4729" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                    <SPLIT distance="100" swimtime="00:01:20.01" />
                    <SPLIT distance="150" swimtime="00:02:02.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1575" points="689" swimtime="00:01:15.67" resultid="2836" heatid="4768" lane="3" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1477" points="672" swimtime="00:01:10.56" resultid="2837" heatid="4786" lane="2" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Kaczmarek" birthdate="1977-06-25" gender="M" nation="POL" athleteid="2838">
              <RESULTS>
                <RESULT eventid="1143" points="844" swimtime="00:01:00.31" resultid="2839" heatid="4690" lane="3" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1255" status="DNS" swimtime="00:00:00.00" resultid="2840" heatid="4725" lane="2" entrytime="00:00:57.50" />
                <RESULT eventid="1379" points="840" swimtime="00:00:25.84" resultid="2841" heatid="4751" lane="2" entrytime="00:00:25.50" />
                <RESULT eventid="1519" points="916" swimtime="00:00:27.01" resultid="2842" heatid="4803" lane="4" entrytime="00:00:26.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1350" points="717" swimtime="00:01:49.99" resultid="2866" heatid="4740" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.39" />
                    <SPLIT distance="100" swimtime="00:00:57.64" />
                    <SPLIT distance="150" swimtime="00:01:25.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2838" number="1" />
                    <RELAYPOSITION athleteid="2818" number="2" />
                    <RELAYPOSITION athleteid="2856" number="3" />
                    <RELAYPOSITION athleteid="2843" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1325" points="710" swimtime="00:03:52.55" resultid="3548" heatid="4737" lane="2" entrytime="00:03:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.21" />
                    <SPLIT distance="100" swimtime="00:00:56.25" />
                    <SPLIT distance="150" swimtime="00:01:22.90" />
                    <SPLIT distance="200" swimtime="00:01:53.01" />
                    <SPLIT distance="250" swimtime="00:02:24.07" />
                    <SPLIT distance="300" swimtime="00:02:57.89" />
                    <SPLIT distance="350" swimtime="00:03:24.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2838" number="1" />
                    <RELAYPOSITION athleteid="2856" number="2" />
                    <RELAYPOSITION athleteid="2861" number="3" />
                    <RELAYPOSITION athleteid="2843" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1329" status="DNS" swimtime="00:00:00.00" resultid="2867" heatid="4738" lane="3" entrytime="00:02:05.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2828" number="1" />
                    <RELAYPOSITION athleteid="2851" number="2" />
                    <RELAYPOSITION athleteid="2848" number="3" />
                    <RELAYPOSITION athleteid="2833" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="NIEGOR" nation="POL" region="04" clubid="2791" name="Zawodnik Niezrzeszony Gorzów Wlkp." shortname="Zawodnik Niezrzeszony Gorzów W">
          <ATHLETES>
            <ATHLETE firstname="Bartłomiej" lastname="Karpisz" birthdate="1993-04-17" gender="M" nation="POL" athleteid="2792">
              <RESULTS>
                <RESULT eventid="1102" points="694" swimtime="00:00:24.04" resultid="2793" heatid="4682" lane="2" entrytime="00:00:24.00" />
                <RESULT eventid="1255" points="772" swimtime="00:00:56.02" resultid="2794" heatid="4725" lane="3" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="778" swimtime="00:00:25.17" resultid="2795" heatid="4751" lane="3" entrytime="00:00:25.00" />
                <RESULT eventid="1491" points="776" swimtime="00:00:57.43" resultid="2796" heatid="4794" lane="3" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZSWRO" nation="POL" region="01" clubid="3050" name="KS AZS AWF Wrocław">
          <CONTACT city="Wrocław" email="andrzwejklarowicz@gmail.com" name="Klarowicz" phone="661443902" state="DOLNO" street="Paderewskiego 35" zip="51-612" />
          <ATHLETES>
            <ATHLETE firstname="Dominika" lastname="Sasin" birthdate="1994-05-29" gender="F" nation="POL" license="100201600097" athleteid="3051">
              <RESULTS>
                <RESULT eventid="1059" points="734" swimtime="00:00:27.71" resultid="3052" heatid="4669" lane="5" entrytime="00:00:27.20" />
                <RESULT eventid="1185" points="712" swimtime="00:02:13.69" resultid="3053" heatid="4708" lane="3" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.18" />
                    <SPLIT distance="100" swimtime="00:01:04.31" />
                    <SPLIT distance="150" swimtime="00:01:39.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="722" swimtime="00:00:29.14" resultid="3054" heatid="4743" lane="4" entrytime="00:00:28.70" />
                <RESULT eventid="1393" points="740" swimtime="00:01:00.18" resultid="3055" heatid="4756" lane="3" entrytime="00:00:58.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TROPUL" nation="POL" region="03" clubid="2709" name="UKS TRÓJKA Puławy">
          <CONTACT city="Puławy" name="Gogacz" phone="506694816" state="LUBEL" />
          <ATHLETES>
            <ATHLETE firstname="Sebastian" lastname="Gogacz" birthdate="1976-10-28" gender="M" nation="POL" license="501203700057" athleteid="2710">
              <RESULTS>
                <RESULT eventid="1283" points="477" swimtime="00:02:53.34" resultid="2711" heatid="4733" lane="6" entrytime="00:02:51.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.09" />
                    <SPLIT distance="100" swimtime="00:01:24.03" />
                    <SPLIT distance="150" swimtime="00:02:09.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="548" swimtime="00:02:32.74" resultid="2712" heatid="4782" lane="2" entrytime="00:02:35.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                    <SPLIT distance="100" swimtime="00:01:12.76" />
                    <SPLIT distance="150" swimtime="00:01:52.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="507" swimtime="00:05:04.79" resultid="2713" heatid="4807" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.71" />
                    <SPLIT distance="100" swimtime="00:01:14.03" />
                    <SPLIT distance="150" swimtime="00:01:52.81" />
                    <SPLIT distance="200" swimtime="00:02:31.70" />
                    <SPLIT distance="250" swimtime="00:03:10.43" />
                    <SPLIT distance="300" swimtime="00:03:48.98" />
                    <SPLIT distance="350" swimtime="00:04:27.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MUZGI" nation="POL" region="05" clubid="2717" name="MUKS Zgierz">
          <CONTACT city="ZGIERZ" email="roman.wiczel@gmail.com" name="WICZEL" phone="691-928-922" state="ŁÓDZK" street="ANDRZEJA 14" zip="95-100" />
          <ATHLETES>
            <ATHLETE firstname="Małgorzata" lastname="Ścibiorek" birthdate="1971-09-12" gender="F" nation="POL" license="502805600026" athleteid="3416">
              <RESULTS>
                <RESULT eventid="1241" points="783" swimtime="00:01:12.57" resultid="3417" heatid="4719" lane="4" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="714" swimtime="00:00:32.73" resultid="3418" heatid="4743" lane="6" entrytime="00:00:32.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Sypniewski" birthdate="1957-02-01" gender="M" nation="POL" license="102805700035" athleteid="3389">
              <RESULTS>
                <RESULT eventid="1171" points="475" swimtime="00:00:41.66" resultid="3390" heatid="4698" lane="2" entrytime="00:00:41.00" entrycourse="SCM" />
                <RESULT eventid="1283" points="414" swimtime="00:03:30.38" resultid="3391" heatid="4731" lane="4" entrytime="00:03:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.11" />
                    <SPLIT distance="100" swimtime="00:01:39.90" />
                    <SPLIT distance="150" swimtime="00:02:35.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1589" points="433" swimtime="00:01:34.91" resultid="3392" heatid="4771" lane="1" entrytime="00:01:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="450" swimtime="00:01:25.41" resultid="3393" heatid="4789" lane="2" entrytime="00:01:26.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zdzisław" lastname="Jasiński" birthdate="1960-07-23" gender="M" nation="POL" license="502805700027" athleteid="3402">
              <RESULTS>
                <RESULT eventid="1102" points="357" swimtime="00:00:35.09" resultid="3403" heatid="4674" lane="1" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1171" points="317" swimtime="00:00:46.22" resultid="3404" heatid="4697" lane="3" entrytime="00:00:43.00" entrycourse="SCM" />
                <RESULT eventid="1407" points="359" swimtime="00:01:18.63" resultid="3405" heatid="4759" lane="3" entrytime="00:01:19.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="317" swimtime="00:01:34.21" resultid="3406" heatid="4790" lane="1" entrytime="00:01:23.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Klarecka" birthdate="1977-06-06" gender="F" nation="POL" license="502805600" athleteid="3362">
              <RESULTS>
                <RESULT eventid="1213" points="254" swimtime="00:03:43.60" resultid="3363" heatid="4714" lane="4" entrytime="00:03:39.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.43" />
                    <SPLIT distance="100" swimtime="00:01:52.98" />
                    <SPLIT distance="150" swimtime="00:02:53.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1269" points="333" swimtime="00:03:47.86" resultid="3364" heatid="4727" lane="4" entrytime="00:03:47.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.31" />
                    <SPLIT distance="100" swimtime="00:01:49.86" />
                    <SPLIT distance="150" swimtime="00:02:48.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="232" swimtime="00:03:53.01" resultid="3365" heatid="4780" lane="4" entrytime="00:03:46.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.93" />
                    <SPLIT distance="100" swimtime="00:01:49.73" />
                    <SPLIT distance="150" swimtime="00:02:52.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1533" points="268" swimtime="00:06:50.92" resultid="3366" heatid="4804" lane="3" entrytime="00:07:00.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.33" />
                    <SPLIT distance="100" swimtime="00:01:37.64" />
                    <SPLIT distance="150" swimtime="00:02:29.85" />
                    <SPLIT distance="200" swimtime="00:03:22.97" />
                    <SPLIT distance="250" swimtime="00:04:16.24" />
                    <SPLIT distance="300" swimtime="00:05:09.71" />
                    <SPLIT distance="350" swimtime="00:06:02.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Morozowski" birthdate="1973-05-09" gender="M" nation="POL" license="102805700051" athleteid="3381">
              <RESULTS>
                <RESULT eventid="1171" status="DNS" swimtime="00:00:00.00" resultid="3382" heatid="4699" lane="2" entrytime="00:00:39.30" entrycourse="SCM" />
                <RESULT eventid="1283" swimtime="00:00:00.00" resultid="3383" entrytime="00:03:27.10" entrycourse="SCM" />
                <RESULT eventid="1589" status="DNS" swimtime="00:00:00.00" resultid="3384" heatid="4771" lane="4" entrytime="00:01:29.22" entrycourse="SCM" />
                <RESULT eventid="1547" status="DNS" swimtime="00:00:00.00" resultid="3385" heatid="4809" lane="1" entrytime="00:05:58.59" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Matczak" birthdate="1989-08-12" gender="M" nation="POL" license="502805700" athleteid="3423">
              <RESULTS>
                <RESULT eventid="1171" points="678" swimtime="00:00:30.41" resultid="3424" heatid="4704" lane="5" entrytime="00:00:30.02" entrycourse="SCM" />
                <RESULT eventid="1283" points="679" swimtime="00:02:29.21" resultid="3425" heatid="4734" lane="1" entrytime="00:02:39.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                    <SPLIT distance="100" swimtime="00:01:11.69" />
                    <SPLIT distance="150" swimtime="00:01:50.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1589" points="704" swimtime="00:01:06.43" resultid="3426" heatid="4775" lane="1" entrytime="00:01:07.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek-Maciej" lastname="Dziedziczak" birthdate="1977-02-04" gender="M" nation="POL" license="502805700" athleteid="3399">
              <RESULTS>
                <RESULT eventid="1407" points="361" swimtime="00:01:10.23" resultid="3400" heatid="4760" lane="1" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="257" swimtime="00:06:22.44" resultid="3401" heatid="4808" lane="6" entrytime="00:08:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                    <SPLIT distance="100" swimtime="00:01:21.91" />
                    <SPLIT distance="150" swimtime="00:02:09.78" />
                    <SPLIT distance="200" swimtime="00:02:59.71" />
                    <SPLIT distance="250" swimtime="00:03:50.32" />
                    <SPLIT distance="300" swimtime="00:04:42.31" />
                    <SPLIT distance="350" swimtime="00:05:34.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robert" lastname="Szalbierz" birthdate="1968-08-06" gender="M" nation="POL" license="502805700034" athleteid="3432">
              <RESULTS>
                <RESULT eventid="1102" points="443" swimtime="00:00:30.68" resultid="3433" heatid="4676" lane="6" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="1379" points="443" swimtime="00:00:33.44" resultid="3434" heatid="4747" lane="1" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1491" points="405" swimtime="00:01:18.00" resultid="3435" heatid="4790" lane="3" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Wiśniewska" birthdate="1981-02-02" gender="F" nation="POL" license="502805600123" athleteid="3412">
              <RESULTS>
                <RESULT eventid="1059" points="122" swimtime="00:00:52.46" resultid="3413" heatid="4665" lane="4" entrytime="00:00:52.00" entrycourse="SCM" />
                <RESULT eventid="1157" points="139" swimtime="00:01:02.07" resultid="3414" heatid="4691" lane="4" entrytime="00:01:02.00" entrycourse="SCM" />
                <RESULT eventid="1575" points="132" swimtime="00:02:17.30" resultid="3415" heatid="4765" lane="4" entrytime="00:02:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Węgrzycka" birthdate="1977-01-26" gender="F" nation="POL" license="502805600056" athleteid="3419">
              <RESULTS>
                <RESULT eventid="1059" points="259" swimtime="00:00:41.24" resultid="3420" heatid="4666" lane="5" entrytime="00:00:39.00" entrycourse="SCM" />
                <RESULT eventid="1185" points="164" swimtime="00:03:50.13" resultid="3421" heatid="4706" lane="5" entrytime="00:03:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.72" />
                    <SPLIT distance="100" swimtime="00:01:46.96" />
                    <SPLIT distance="150" swimtime="00:02:48.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="160" swimtime="00:01:46.63" resultid="3422" heatid="4753" lane="1" entrytime="00:01:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Justyna" lastname="Barańska" birthdate="1977-05-01" gender="F" nation="POL" license="502805600055" athleteid="3367">
              <RESULTS>
                <RESULT eventid="1157" points="343" swimtime="00:00:47.14" resultid="3368" heatid="4693" lane="6" entrytime="00:00:44.00" entrycourse="SCM" />
                <RESULT eventid="1269" points="373" swimtime="00:03:39.49" resultid="3369" heatid="4727" lane="3" entrytime="00:03:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.18" />
                    <SPLIT distance="100" swimtime="00:01:48.29" />
                    <SPLIT distance="150" swimtime="00:02:45.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1575" points="311" swimtime="00:01:44.29" resultid="3370" heatid="4767" lane="1" entrytime="00:01:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Urszula" lastname="Mróz" birthdate="1962-03-03" gender="F" nation="POL" license="502805600024" athleteid="3371">
              <RESULTS>
                <RESULT eventid="1059" points="591" swimtime="00:00:33.96" resultid="3372" heatid="4667" lane="2" entrytime="00:00:33.60" entrycourse="SCM" />
                <RESULT eventid="1157" points="575" swimtime="00:00:44.60" resultid="3373" heatid="4693" lane="1" entrytime="00:00:43.30" entrycourse="SCM" />
                <RESULT eventid="1358" points="623" swimtime="00:00:36.57" resultid="3374" heatid="4742" lane="1" entrytime="00:00:34.60" entrycourse="SCM" />
                <RESULT eventid="1477" points="588" swimtime="00:01:26.18" resultid="3375" heatid="4785" lane="1" entrytime="00:01:21.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jarosław" lastname="Woźniak" birthdate="1980-09-30" gender="M" nation="POL" license="502805700" athleteid="3407">
              <RESULTS>
                <RESULT eventid="1102" points="288" swimtime="00:00:34.46" resultid="3408" heatid="4673" lane="1" entrytime="00:00:34.00" entrycourse="SCM" />
                <RESULT eventid="1171" points="242" swimtime="00:00:45.00" resultid="3409" heatid="4698" lane="6" entrytime="00:00:43.00" entrycourse="SCM" />
                <RESULT eventid="1589" points="234" swimtime="00:01:39.69" resultid="3410" heatid="4770" lane="2" entrytime="00:01:43.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="210" swimtime="00:01:35.73" resultid="3411" heatid="4789" lane="6" entrytime="00:01:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Rembowska-Świeboda" birthdate="1968-06-27" gender="F" nation="POL" license="102805600031" athleteid="3376">
              <RESULTS>
                <RESULT eventid="1059" points="474" swimtime="00:00:33.70" resultid="3377" heatid="4667" lane="5" entrytime="00:00:34.90" entrycourse="SCM" />
                <RESULT eventid="1129" points="501" swimtime="00:01:22.94" resultid="3378" heatid="4684" lane="4" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="466" swimtime="00:01:15.56" resultid="3379" heatid="4754" lane="1" entrytime="00:01:19.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1505" points="505" swimtime="00:00:38.00" resultid="3380" heatid="4797" lane="5" entrytime="00:00:38.90" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Włodzimierz" lastname="Przytulski" birthdate="1957-01-09" gender="M" nation="POL" license="502805700049" athleteid="3394">
              <RESULTS>
                <RESULT eventid="1102" points="503" swimtime="00:00:31.97" resultid="3395" heatid="4675" lane="6" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1255" points="475" swimtime="00:01:23.77" resultid="3396" heatid="4721" lane="2" entrytime="00:01:21.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="560" swimtime="00:00:34.76" resultid="3397" heatid="4747" lane="6" entrytime="00:00:33.05" entrycourse="SCM" />
                <RESULT eventid="1519" points="511" swimtime="00:00:37.95" resultid="3398" heatid="4801" lane="5" entrytime="00:00:37.50" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Gołębiowski" birthdate="1996-05-20" gender="M" nation="POL" license="502805700" athleteid="3427">
              <RESULTS>
                <RESULT eventid="1102" points="502" swimtime="00:00:26.77" resultid="3428" heatid="4678" lane="1" entrytime="00:00:28.00" entrycourse="SCM" />
                <RESULT eventid="1171" points="503" swimtime="00:00:33.94" resultid="3429" heatid="4702" lane="4" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1589" points="434" swimtime="00:01:16.79" resultid="3430" heatid="4773" lane="5" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="461" swimtime="00:01:08.33" resultid="3431" heatid="4789" lane="4" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Gajda" birthdate="1978-02-23" gender="M" nation="POL" license="502805700059" athleteid="3436">
              <RESULTS>
                <RESULT eventid="1171" points="359" swimtime="00:00:39.49" resultid="3437" heatid="4698" lane="3" entrytime="00:00:40.47" entrycourse="SCM" />
                <RESULT eventid="1589" points="273" swimtime="00:01:34.66" resultid="3438" heatid="4771" lane="2" entrytime="00:01:30.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1519" points="339" swimtime="00:00:36.54" resultid="3439" heatid="4801" lane="3" entrytime="00:00:35.39" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1350" points="538" swimtime="00:02:14.50" resultid="3441" heatid="4739" lane="3" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.32" />
                    <SPLIT distance="100" swimtime="00:01:07.46" />
                    <SPLIT distance="150" swimtime="00:01:43.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3394" number="1" />
                    <RELAYPOSITION athleteid="3423" number="2" />
                    <RELAYPOSITION athleteid="3389" number="3" />
                    <RELAYPOSITION athleteid="3436" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1325" points="376" swimtime="00:05:05.05" resultid="3442" heatid="4736" lane="3" entrytime="00:05:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                    <SPLIT distance="100" swimtime="00:01:12.25" />
                    <SPLIT distance="150" swimtime="00:01:50.57" />
                    <SPLIT distance="200" swimtime="00:02:33.10" />
                    <SPLIT distance="250" swimtime="00:03:09.53" />
                    <SPLIT distance="300" swimtime="00:03:51.33" />
                    <SPLIT distance="350" swimtime="00:04:27.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3432" number="1" />
                    <RELAYPOSITION athleteid="3402" number="2" />
                    <RELAYPOSITION athleteid="3389" number="3" />
                    <RELAYPOSITION athleteid="3436" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1329" points="599" swimtime="00:02:30.07" resultid="3440" heatid="4738" lane="2" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                    <SPLIT distance="100" swimtime="00:01:23.84" />
                    <SPLIT distance="150" swimtime="00:01:56.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3376" number="1" />
                    <RELAYPOSITION athleteid="3367" number="2" />
                    <RELAYPOSITION athleteid="3416" number="3" />
                    <RELAYPOSITION athleteid="3371" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="EXTOBO" nation="POL" region="15" clubid="2197" name="KS EXTREME TEAM Oborniki">
          <CONTACT city="Oborniki" email="JANWOL2212@GMAIL.COM" name="WOLNIEWICZ" phone="791064667" state="WIELK" street="CZARNKOWSKA 84" zip="64-600" />
          <ATHLETES>
            <ATHLETE firstname="Janusz" lastname="Wolniewicz" birthdate="1948-12-22" gender="M" nation="POL" athleteid="2198">
              <RESULTS>
                <RESULT eventid="1102" points="336" swimtime="00:00:38.68" resultid="2199" heatid="4672" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="1199" points="209" swimtime="00:03:40.57" resultid="2200" heatid="4710" lane="1" entrytime="00:03:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.88" />
                    <SPLIT distance="100" swimtime="00:01:46.81" />
                    <SPLIT distance="150" swimtime="00:02:44.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="286" swimtime="00:01:33.60" resultid="2201" heatid="4758" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="229" swimtime="00:08:05.55" resultid="2202" heatid="4808" lane="1" entrytime="00:07:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.31" />
                    <SPLIT distance="100" swimtime="00:01:53.10" />
                    <SPLIT distance="150" swimtime="00:02:54.76" />
                    <SPLIT distance="200" swimtime="00:03:57.76" />
                    <SPLIT distance="250" swimtime="00:05:00.70" />
                    <SPLIT distance="300" swimtime="00:06:03.92" />
                    <SPLIT distance="350" swimtime="00:07:06.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIEKRA" nation="POL" region="06" clubid="2314" name="Zawodnik Niezrzeszony Kraków">
          <ATHLETES>
            <ATHLETE firstname="Szymon" lastname="Klimkowski" birthdate="1994-02-07" gender="M" nation="POL" athleteid="2315">
              <RESULTS>
                <RESULT eventid="1379" status="DNS" swimtime="00:00:00.00" resultid="2316" heatid="4746" lane="4" entrytime="00:00:33.47" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="2317" heatid="4789" lane="5" entrytime="00:01:26.29" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Wesołowski" birthdate="1971-12-10" gender="M" nation="POL" athleteid="3352">
              <RESULTS>
                <RESULT eventid="1102" points="459" swimtime="00:00:30.32" resultid="3358" heatid="4673" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="1199" points="361" swimtime="00:02:40.98" resultid="3359" heatid="4711" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                    <SPLIT distance="100" swimtime="00:01:16.68" />
                    <SPLIT distance="150" swimtime="00:01:59.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="376" swimtime="00:00:35.32" resultid="3360" heatid="4745" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="1407" points="445" swimtime="00:01:07.42" resultid="3361" heatid="4761" lane="4" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bogdan" lastname="Szczurek" birthdate="1952-02-07" gender="M" nation="POL" athleteid="3353">
              <RESULTS>
                <RESULT eventid="1102" points="182" swimtime="00:00:47.41" resultid="3354" heatid="4670" lane="3" entrytime="00:00:50.00" />
                <RESULT eventid="1143" points="182" swimtime="00:02:06.15" resultid="3355" heatid="4686" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="153" swimtime="00:01:55.44" resultid="3356" heatid="4758" lane="2" entrytime="00:01:55.00" />
                <RESULT eventid="1435" points="176" swimtime="00:04:36.50" resultid="3506" heatid="4777" lane="3" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.49" />
                    <SPLIT distance="100" swimtime="00:02:14.06" />
                    <SPLIT distance="150" swimtime="00:03:26.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00211" nation="POL" region="11" clubid="3230" name="KS Górnik Radlin">
          <CONTACT city="Radlin" name="Cymerman, Jakub" state="ŚLĄSK" />
          <ATHLETES>
            <ATHLETE firstname="Ryszard" lastname="Kubica" birthdate="1972-02-22" gender="M" nation="POL" license="100211700343" athleteid="3231">
              <RESULTS>
                <RESULT eventid="1143" points="416" swimtime="00:01:17.60" resultid="3232" heatid="4688" lane="2" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1255" points="440" swimtime="00:01:14.63" resultid="3233" heatid="4722" lane="5" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1435" points="388" swimtime="00:02:54.33" resultid="3234" heatid="4778" lane="5" entrytime="00:02:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.25" />
                    <SPLIT distance="100" swimtime="00:01:24.83" />
                    <SPLIT distance="150" swimtime="00:02:10.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="390" swimtime="00:05:34.61" resultid="3235" heatid="4809" lane="4" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                    <SPLIT distance="100" swimtime="00:01:17.85" />
                    <SPLIT distance="150" swimtime="00:02:00.78" />
                    <SPLIT distance="200" swimtime="00:02:44.24" />
                    <SPLIT distance="250" swimtime="00:03:27.70" />
                    <SPLIT distance="300" swimtime="00:04:10.84" />
                    <SPLIT distance="350" swimtime="00:04:53.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="JUVBIA" nation="POL" region="09" clubid="2203" name="MKS JUVENIA Białystok">
          <CONTACT city="Białystok" email="wzmasters@wp.pl" name="Żmiejko" phone="797309140" />
          <ATHLETES>
            <ATHLETE firstname="Dominika" lastname="Michalik" birthdate="1979-01-01" gender="F" nation="POL" athleteid="2204">
              <RESULTS>
                <RESULT eventid="1185" points="654" swimtime="00:02:24.33" resultid="2205" heatid="4708" lane="4" entrytime="00:02:19.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                    <SPLIT distance="100" swimtime="00:01:08.87" />
                    <SPLIT distance="150" swimtime="00:01:46.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="656" swimtime="00:01:05.69" resultid="2206" heatid="4756" lane="6" entrytime="00:01:04.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1533" points="616" swimtime="00:05:07.58" resultid="2207" heatid="4806" lane="4" entrytime="00:04:56.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="100" swimtime="00:01:15.95" />
                    <SPLIT distance="150" swimtime="00:01:55.37" />
                    <SPLIT distance="200" swimtime="00:02:34.78" />
                    <SPLIT distance="250" swimtime="00:03:14.12" />
                    <SPLIT distance="300" swimtime="00:03:53.86" />
                    <SPLIT distance="350" swimtime="00:04:31.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Żmiejko" birthdate="1963-01-01" gender="M" nation="POL" athleteid="2208">
              <RESULTS>
                <RESULT eventid="1102" points="611" swimtime="00:00:28.72" resultid="2209" heatid="4677" lane="4" entrytime="00:00:28.75" />
                <RESULT eventid="1255" points="597" swimtime="00:01:11.00" resultid="2210" heatid="4722" lane="2" entrytime="00:01:10.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="611" swimtime="00:00:31.14" resultid="2211" heatid="4748" lane="2" entrytime="00:00:30.95" />
                <RESULT eventid="1491" points="591" swimtime="00:01:13.03" resultid="2212" heatid="4792" lane="6" entrytime="00:01:11.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIEWAR" nation="POL" region="14" clubid="2235" name="Zawodnik Niezrzeszony Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Tobiasz" lastname="Jankowski" birthdate="1983-05-12" gender="M" nation="POL" athleteid="2236">
              <RESULTS>
                <RESULT eventid="1171" points="325" swimtime="00:00:38.78" resultid="2237" heatid="4699" lane="6" entrytime="00:00:40.00" />
                <RESULT eventid="1227" points="279" swimtime="00:03:03.46" resultid="2238" heatid="4716" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                    <SPLIT distance="100" swimtime="00:01:27.33" />
                    <SPLIT distance="150" swimtime="00:02:20.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="304" swimtime="00:00:34.37" resultid="2239" heatid="4745" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1589" points="339" swimtime="00:01:26.37" resultid="2240" heatid="4771" lane="3" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIEKAT" nation="POL" region="11" clubid="2457" name="Zawodnik Niezrzeszony Katowice">
          <ATHLETES>
            <ATHLETE firstname="Łukasz" lastname="Rogoziński" birthdate="1986-02-16" gender="M" nation="POL" athleteid="2458">
              <RESULTS>
                <RESULT eventid="1171" points="132" swimtime="00:00:52.38" resultid="2459" heatid="4695" lane="3" />
                <RESULT eventid="1283" points="136" swimtime="00:04:23.40" resultid="2460" heatid="4730" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.67" />
                    <SPLIT distance="100" swimtime="00:02:04.72" />
                    <SPLIT distance="150" swimtime="00:03:12.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1589" points="127" swimtime="00:01:59.90" resultid="2461" heatid="4769" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="84" swimtime="00:02:05.32" resultid="2462" heatid="4787" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Opałko" birthdate="1999-07-06" gender="F" nation="POL" athleteid="2553">
              <RESULTS>
                <RESULT eventid="1213" swimtime="00:02:47.97" resultid="2554" heatid="4715" lane="4" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.20" />
                    <SPLIT distance="100" swimtime="00:01:17.61" />
                    <SPLIT distance="150" swimtime="00:02:05.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1269" swimtime="00:03:07.28" resultid="2555" heatid="4728" lane="4" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.98" />
                    <SPLIT distance="100" swimtime="00:01:27.98" />
                    <SPLIT distance="150" swimtime="00:02:17.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1421" swimtime="00:02:56.71" resultid="2556" heatid="4776" lane="2" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.51" />
                    <SPLIT distance="100" swimtime="00:01:24.53" />
                    <SPLIT distance="150" swimtime="00:02:10.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1477" swimtime="00:01:16.24" resultid="2557" heatid="4786" lane="6" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Władyka" birthdate="2002-04-20" gender="M" nation="POL" athleteid="2558">
              <RESULTS>
                <RESULT eventid="1102" swimtime="00:00:25.30" resultid="2559" heatid="4682" lane="5" entrytime="00:00:24.22" />
                <RESULT eventid="1171" swimtime="00:00:29.77" resultid="2560" heatid="4704" lane="3" entrytime="00:00:28.05" />
                <RESULT eventid="1589" swimtime="00:01:05.24" resultid="2561" heatid="4775" lane="3" entrytime="00:01:01.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" swimtime="00:01:02.47" resultid="2562" heatid="4794" lane="4" entrytime="00:00:59.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksander" lastname="Ludynia" birthdate="1979-10-23" gender="M" nation="POL" athleteid="2814">
              <RESULTS>
                <RESULT eventid="1102" points="410" swimtime="00:00:30.63" resultid="2815" heatid="4676" lane="1" entrytime="00:00:29.90" />
                <RESULT eventid="1407" points="363" swimtime="00:01:09.56" resultid="2816" heatid="4761" lane="3" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Tokarski" birthdate="1996-07-12" gender="M" nation="POL" athleteid="3262">
              <RESULTS>
                <RESULT eventid="1171" points="845" swimtime="00:00:28.55" resultid="3263" heatid="4704" lane="6" entrytime="00:00:31.00" />
                <RESULT eventid="1283" points="707" swimtime="00:02:23.21" resultid="3264" heatid="4734" lane="2" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                    <SPLIT distance="100" swimtime="00:01:09.12" />
                    <SPLIT distance="150" swimtime="00:01:47.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1589" points="776" swimtime="00:01:03.27" resultid="3265" heatid="4774" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominika" lastname="Karpińska" birthdate="1991-07-26" gender="F" nation="POL" athleteid="2714">
              <RESULTS>
                <RESULT eventid="1059" points="668" swimtime="00:00:28.79" resultid="2715" heatid="4668" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1393" points="647" swimtime="00:01:03.29" resultid="2716" heatid="4755" lane="2" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiesław" lastname="Majcher" birthdate="1950-09-19" gender="M" nation="POL" athleteid="3225">
              <RESULTS>
                <RESULT eventid="1102" points="129" swimtime="00:00:53.25" resultid="3226" heatid="4670" lane="1" />
                <RESULT eventid="1407" status="DNS" swimtime="00:00:00.00" resultid="3228" heatid="4757" lane="2" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="3229" heatid="4787" lane="4" />
                <RESULT eventid="1283" points="131" swimtime="00:05:46.18" resultid="4820" heatid="4732" lane="1" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.65" />
                    <SPLIT distance="100" swimtime="00:02:43.97" />
                    <SPLIT distance="150" swimtime="00:04:14.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Korzuchowski" birthdate="1999-10-16" gender="M" nation="POL" athleteid="2548">
              <RESULTS>
                <RESULT eventid="1143" swimtime="00:01:08.65" resultid="2549" heatid="4690" lane="6" entrytime="00:01:07.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" swimtime="00:02:38.19" resultid="2550" heatid="4717" lane="2" entrytime="00:02:37.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.41" />
                    <SPLIT distance="100" swimtime="00:01:09.52" />
                    <SPLIT distance="150" swimtime="00:02:00.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1435" swimtime="00:02:35.10" resultid="2551" heatid="4778" lane="3" entrytime="00:02:35.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                    <SPLIT distance="100" swimtime="00:01:16.04" />
                    <SPLIT distance="150" swimtime="00:01:56.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1519" swimtime="00:00:30.65" resultid="2552" heatid="4802" lane="3" entrytime="00:00:31.51" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIEZOR" nation="POL" region="11" clubid="2463" name="Zawodnik Niezrzeszony Żory">
          <ATHLETES>
            <ATHLETE firstname="Krzysztof" lastname="Drózd" birthdate="1992-12-02" gender="M" nation="POL" athleteid="2464">
              <RESULTS>
                <RESULT eventid="1102" points="521" swimtime="00:00:26.76" resultid="2465" heatid="4679" lane="3" entrytime="00:00:26.43" />
                <RESULT eventid="1143" points="414" swimtime="00:01:10.53" resultid="2466" heatid="4689" lane="5" entrytime="00:01:10.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1435" points="339" swimtime="00:02:43.82" resultid="2467" heatid="4777" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.33" />
                    <SPLIT distance="100" swimtime="00:01:18.72" />
                    <SPLIT distance="150" swimtime="00:02:01.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1519" points="403" swimtime="00:00:32.30" resultid="2468" heatid="4802" lane="4" entrytime="00:00:31.67" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LEGWAR" nation="POL" region="14" clubid="3843" name="Legia Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Bogdan" lastname="Dubiński" birthdate="1953-05-05" gender="M" nation="POL" athleteid="3844">
              <RESULTS>
                <RESULT eventid="1102" points="363" swimtime="00:00:35.65" resultid="3845" heatid="4672" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="1199" points="306" swimtime="00:03:09.24" resultid="3846" heatid="4709" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.56" />
                    <SPLIT distance="100" swimtime="00:01:27.41" />
                    <SPLIT distance="150" swimtime="00:02:19.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="357" swimtime="00:01:21.47" resultid="3847" heatid="4759" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1519" points="326" swimtime="00:00:44.10" resultid="3848" heatid="4801" lane="6" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIEPOL" nation="POL" region="12" clubid="2241" name="Zawodnik Niezrzeszony Połaniec">
          <ATHLETES>
            <ATHLETE firstname="Anna" lastname="Gad" birthdate="1997-05-26" gender="F" nation="POL" athleteid="2242">
              <RESULTS>
                <RESULT eventid="1059" points="565" swimtime="00:00:30.24" resultid="2243" heatid="4668" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1393" points="532" swimtime="00:01:07.19" resultid="2244" heatid="4755" lane="4" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="464" swimtime="00:00:33.77" resultid="2245" heatid="4742" lane="2" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ISWBIA" nation="POL" region="09" clubid="3131" name="iSwim Białystok">
          <CONTACT city="Białystok" email="biuro@iswim.bialystok.pl" name="Sebastian Humbla" phone="535309915" state="PODLA" street="Wierzbowa 3c" zip="15-743" />
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Daszuta" birthdate="1973-03-12" gender="M" nation="POL" athleteid="3137">
              <RESULTS>
                <RESULT eventid="1171" points="555" swimtime="00:00:34.86" resultid="3138" heatid="4702" lane="5" entrytime="00:00:33.50" />
                <RESULT eventid="1379" points="521" swimtime="00:00:30.30" resultid="3139" heatid="4748" lane="3" entrytime="00:00:29.50" />
                <RESULT eventid="1519" status="DNS" swimtime="00:00:00.00" resultid="3140" heatid="4802" lane="5" entrytime="00:00:33.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Świderski" birthdate="1979-02-13" gender="M" nation="POL" athleteid="3141">
              <RESULTS>
                <RESULT eventid="1102" points="663" swimtime="00:00:26.09" resultid="3142" heatid="4681" lane="1" entrytime="00:00:25.40" />
                <RESULT eventid="1255" status="DNS" swimtime="00:00:00.00" resultid="3143" heatid="4724" lane="1" entrytime="00:01:01.79" />
                <RESULT eventid="1379" points="653" swimtime="00:00:27.82" resultid="3144" heatid="4750" lane="5" entrytime="00:00:27.48" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="3145" heatid="4794" lane="5" entrytime="00:01:03.43" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sebastian" lastname="Humbla" birthdate="1979-01-29" gender="M" nation="POL" athleteid="3132">
              <RESULTS>
                <RESULT eventid="1102" status="DNS" swimtime="00:00:00.00" resultid="3133" heatid="4680" lane="3" entrytime="00:00:25.50" />
                <RESULT eventid="1171" status="DNS" swimtime="00:00:00.00" resultid="3134" heatid="4702" lane="2" entrytime="00:00:33.20" />
                <RESULT eventid="1379" status="DNS" swimtime="00:00:00.00" resultid="3135" heatid="4750" lane="1" entrytime="00:00:27.70" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="3136" heatid="4793" lane="1" entrytime="00:01:07.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elżbieta" lastname="Piwowarczyk" birthdate="1966-01-06" gender="F" nation="POL" athleteid="3149">
              <RESULTS>
                <RESULT eventid="1059" points="467" swimtime="00:00:35.84" resultid="3150" heatid="4667" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="1185" points="431" swimtime="00:02:56.88" resultid="3151" heatid="4707" lane="1" entrytime="00:02:56.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                    <SPLIT distance="100" swimtime="00:01:23.83" />
                    <SPLIT distance="150" swimtime="00:02:10.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="436" swimtime="00:01:19.91" resultid="3152" heatid="4753" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1505" status="DNS" swimtime="00:00:00.00" resultid="3153" heatid="4796" lane="4" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00111" nation="POL" region="11" clubid="2486" name="UKS TRÓJKA Częstochowa">
          <CONTACT city="Częstochowa" email="trojkaczestochowa@o2.pl" name="Gawda" phone="511181791" state="ŚLĄSK" street="Schillera 5" zip="42-200" />
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Gajda" birthdate="1995-04-23" gender="M" nation="POL" license="100111700062" athleteid="3087">
              <RESULTS>
                <RESULT eventid="1102" points="646" swimtime="00:00:24.62" resultid="3088" heatid="4681" lane="3" entrytime="00:00:24.46" />
                <RESULT eventid="1255" points="664" swimtime="00:00:58.88" resultid="3089" heatid="4725" lane="6" entrytime="00:00:59.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="667" swimtime="00:00:26.49" resultid="3090" heatid="4750" lane="3" entrytime="00:00:26.02" />
                <RESULT eventid="1407" points="621" swimtime="00:00:55.59" resultid="3091" heatid="4764" lane="1" entrytime="00:00:54.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrian" lastname="Kozioł" birthdate="1990-08-26" gender="M" nation="POL" license="100111700090" athleteid="3117">
              <RESULTS>
                <RESULT eventid="1102" points="476" swimtime="00:00:27.58" resultid="3118" heatid="4678" lane="3" entrytime="00:00:27.45" />
                <RESULT eventid="1199" status="DNS" swimtime="00:00:00.00" resultid="3119" heatid="4712" lane="5" entrytime="00:02:26.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szymon" lastname="Warwas" birthdate="1995-07-13" gender="M" nation="POL" athleteid="3097">
              <RESULTS>
                <RESULT eventid="1102" points="605" swimtime="00:00:25.16" resultid="3098" heatid="4682" lane="4" entrytime="00:00:23.50" />
                <RESULT eventid="1143" points="495" swimtime="00:01:06.94" resultid="3099" heatid="4690" lane="4" entrytime="00:00:58.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1435" points="396" swimtime="00:02:38.30" resultid="3100" heatid="4779" lane="3" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                    <SPLIT distance="100" swimtime="00:01:14.96" />
                    <SPLIT distance="150" swimtime="00:01:56.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1519" points="516" swimtime="00:00:29.55" resultid="3101" heatid="4803" lane="3" entrytime="00:00:26.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktoria" lastname="Musik" birthdate="1997-08-04" gender="F" nation="POL" license="100111600053" athleteid="3107">
              <RESULTS>
                <RESULT eventid="1059" points="790" swimtime="00:00:27.04" resultid="3108" heatid="4669" lane="4" entrytime="00:00:26.74" />
                <RESULT eventid="1241" points="602" swimtime="00:01:08.82" resultid="3109" heatid="4719" lane="3" entrytime="00:01:07.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="766" swimtime="00:00:59.49" resultid="3110" heatid="4756" lane="2" entrytime="00:00:59.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1477" points="708" swimtime="00:01:09.33" resultid="3111" heatid="4786" lane="3" entrytime="00:01:07.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Krogulec" birthdate="1991-07-31" gender="M" nation="POL" athleteid="3092">
              <RESULTS>
                <RESULT eventid="1143" points="458" swimtime="00:01:08.20" resultid="3093" heatid="4689" lane="3" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1255" status="DNS" swimtime="00:00:00.00" resultid="3094" heatid="4723" lane="2" entrytime="00:01:06.45" />
                <RESULT eventid="1435" points="415" swimtime="00:02:33.06" resultid="3095" heatid="4779" lane="1" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                    <SPLIT distance="100" swimtime="00:01:13.84" />
                    <SPLIT distance="150" swimtime="00:01:53.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1519" points="429" swimtime="00:00:31.64" resultid="3096" heatid="4803" lane="6" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Kurek" birthdate="1994-07-11" gender="M" nation="POL" license="100111700097" athleteid="3102">
              <RESULTS>
                <RESULT eventid="1102" points="480" swimtime="00:00:27.17" resultid="3103" heatid="4678" lane="5" entrytime="00:00:27.73" />
                <RESULT eventid="1171" points="432" swimtime="00:00:35.71" resultid="3104" heatid="4701" lane="1" entrytime="00:00:35.20" />
                <RESULT eventid="1407" points="478" swimtime="00:01:00.64" resultid="3105" heatid="4762" lane="2" entrytime="00:01:01.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="424" swimtime="00:01:10.27" resultid="3106" heatid="4792" lane="3" entrytime="00:01:08.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sonia" lastname="Nowak" birthdate="1996-05-23" gender="F" nation="POL" license="100111600092" athleteid="3112">
              <RESULTS>
                <RESULT eventid="1059" status="DNS" swimtime="00:00:00.00" resultid="3113" heatid="4668" lane="5" entrytime="00:00:30.29" />
                <RESULT eventid="1185" points="548" swimtime="00:02:25.87" resultid="3114" heatid="4708" lane="2" entrytime="00:02:29.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                    <SPLIT distance="100" swimtime="00:01:11.79" />
                    <SPLIT distance="150" swimtime="00:01:49.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="533" swimtime="00:01:07.13" resultid="3115" heatid="4755" lane="5" entrytime="00:01:05.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1533" points="559" swimtime="00:05:10.48" resultid="3116" heatid="4806" lane="2" entrytime="00:05:09.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                    <SPLIT distance="100" swimtime="00:01:17.31" />
                    <SPLIT distance="150" swimtime="00:01:57.42" />
                    <SPLIT distance="200" swimtime="00:02:37.26" />
                    <SPLIT distance="250" swimtime="00:03:16.98" />
                    <SPLIT distance="300" swimtime="00:03:56.59" />
                    <SPLIT distance="350" swimtime="00:04:34.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1325" points="679" swimtime="00:03:52.65" resultid="3120" heatid="4737" lane="3" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.72" />
                    <SPLIT distance="100" swimtime="00:01:00.28" />
                    <SPLIT distance="150" swimtime="00:01:29.69" />
                    <SPLIT distance="200" swimtime="00:02:02.40" />
                    <SPLIT distance="250" swimtime="00:02:28.45" />
                    <SPLIT distance="300" swimtime="00:02:58.49" />
                    <SPLIT distance="350" swimtime="00:03:24.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3102" number="1" />
                    <RELAYPOSITION athleteid="3092" number="2" />
                    <RELAYPOSITION athleteid="3097" number="3" />
                    <RELAYPOSITION athleteid="3087" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1350" points="610" swimtime="00:01:56.69" resultid="3121" heatid="4740" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                    <SPLIT distance="100" swimtime="00:01:06.23" />
                    <SPLIT distance="150" swimtime="00:01:31.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3092" number="1" />
                    <RELAYPOSITION athleteid="3102" number="2" />
                    <RELAYPOSITION athleteid="3087" number="3" />
                    <RELAYPOSITION athleteid="3097" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="03315" nation="POL" region="15" clubid="2563" name="KU AZS UAM Poznań">
          <CONTACT city="Poznań" email="swimteamuam@gmail.com" name="Sterczyński" phone="693840114" state="WIELK" />
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Juszkiewicz" birthdate="1974-05-10" gender="M" nation="POL" athleteid="2564">
              <RESULTS>
                <RESULT eventid="1102" points="355" swimtime="00:00:32.26" resultid="2565" heatid="4674" lane="4" entrytime="00:00:31.63" />
                <RESULT eventid="1407" points="324" swimtime="00:01:12.79" resultid="2566" heatid="4760" lane="2" entrytime="00:01:12.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1519" points="203" swimtime="00:00:44.66" resultid="2567" heatid="4800" lane="5" entrytime="00:00:46.13" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIESLU" nation="POL" region="14" clubid="2912" name="Zawodnik Niezrzeszony Słupno">
          <ATHLETES>
            <ATHLETE firstname="Katarzyna" lastname="Miaśkiewicz" birthdate="1984-12-16" gender="F" nation="POL" athleteid="2913">
              <RESULTS>
                <RESULT eventid="1157" points="251" swimtime="00:00:50.18" resultid="2914" heatid="4692" lane="6" entrytime="00:00:51.10" />
                <RESULT eventid="1269" points="252" swimtime="00:03:58.35" resultid="2915" heatid="4727" lane="5" entrytime="00:04:02.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.85" />
                    <SPLIT distance="100" swimtime="00:01:50.19" />
                    <SPLIT distance="150" swimtime="00:02:53.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00408" nation="POL" region="08" clubid="3298" name="UKS DELFIN MASTERS Tarnobrzeg">
          <CONTACT city="TARNOBRZEG" email="piotr.michalik@i-bs.pl" name="MICHALIK ANGELIKA" state="PODKA" street="SKALNA GÓRA 8/21" street2="TARNOBRZEG" zip="39-400" />
          <ATHLETES>
            <ATHLETE firstname="Patrycja" lastname="Urbaniak" birthdate="1991-03-03" gender="F" nation="POL" license="500408600214" athleteid="3299">
              <RESULTS>
                <RESULT eventid="1213" points="463" swimtime="00:02:52.49" resultid="3300" heatid="4715" lane="2" entrytime="00:02:50.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                    <SPLIT distance="100" swimtime="00:01:20.75" />
                    <SPLIT distance="150" swimtime="00:02:10.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1269" points="421" swimtime="00:03:16.12" resultid="3301" heatid="4729" lane="1" entrytime="00:03:05.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.35" />
                    <SPLIT distance="100" swimtime="00:01:33.82" />
                    <SPLIT distance="150" swimtime="00:02:24.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1575" points="390" swimtime="00:01:31.67" resultid="3302" heatid="4768" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1477" points="471" swimtime="00:01:20.34" resultid="3303" heatid="4786" lane="1" entrytime="00:01:15.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00811" nation="POL" region="11" clubid="2342" name="MKS Pałac Młodzieży Katowice">
          <ATHLETES>
            <ATHLETE firstname="Małgorzata" lastname="Mądry" birthdate="1966-07-14" gender="F" nation="POL" athleteid="2698">
              <RESULTS>
                <RESULT eventid="1129" points="313" swimtime="00:01:38.90" resultid="2699" heatid="4683" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="370" swimtime="00:03:25.86" resultid="2700" heatid="4714" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.02" />
                    <SPLIT distance="100" swimtime="00:01:39.51" />
                    <SPLIT distance="150" swimtime="00:02:39.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1477" points="426" swimtime="00:01:31.82" resultid="2701" heatid="4783" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1533" points="330" swimtime="00:06:41.32" resultid="2702" heatid="4804" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.69" />
                    <SPLIT distance="100" swimtime="00:01:31.28" />
                    <SPLIT distance="150" swimtime="00:02:20.24" />
                    <SPLIT distance="200" swimtime="00:03:10.93" />
                    <SPLIT distance="250" swimtime="00:04:02.75" />
                    <SPLIT distance="300" swimtime="00:04:56.09" />
                    <SPLIT distance="350" swimtime="00:05:49.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Błażej" lastname="Kornaga" birthdate="1986-09-01" gender="M" nation="POL" athleteid="2343">
              <RESULTS>
                <RESULT eventid="1102" points="424" swimtime="00:00:28.66" resultid="2344" heatid="4676" lane="5" entrytime="00:00:29.73" />
                <RESULT eventid="1199" points="383" swimtime="00:02:29.24" resultid="2345" heatid="4711" lane="5" entrytime="00:02:45.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.78" />
                    <SPLIT distance="100" swimtime="00:01:13.36" />
                    <SPLIT distance="150" swimtime="00:01:52.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="386" swimtime="00:01:05.49" resultid="2346" heatid="4761" lane="6" entrytime="00:01:11.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="324" swimtime="00:05:46.36" resultid="2347" heatid="4807" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                    <SPLIT distance="100" swimtime="00:01:21.77" />
                    <SPLIT distance="150" swimtime="00:02:06.22" />
                    <SPLIT distance="200" swimtime="00:02:51.37" />
                    <SPLIT distance="250" swimtime="00:03:35.35" />
                    <SPLIT distance="300" swimtime="00:04:21.55" />
                    <SPLIT distance="350" swimtime="00:05:05.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIEGLI" nation="POL" region="11" clubid="2166" name="Zawodnik Niezrzeszony Gliwice">
          <ATHLETES>
            <ATHLETE firstname="Jerzy" lastname="Marciniszko" birthdate="1944-11-23" gender="M" nation="POL" athleteid="2405">
              <RESULTS>
                <RESULT eventid="1102" points="90" swimtime="00:01:04.12" resultid="2406" heatid="4670" lane="2" entrytime="00:01:05.96" />
                <RESULT eventid="1171" points="207" swimtime="00:01:04.80" resultid="2407" heatid="4696" lane="1" />
                <RESULT eventid="1519" points="82" swimtime="00:01:17.91" resultid="2408" heatid="4799" lane="1" />
                <RESULT eventid="1589" points="131" swimtime="00:02:48.32" resultid="2410" heatid="4769" lane="4" entrytime="00:02:49.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:22.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Musiałowski" birthdate="1995-08-21" gender="M" nation="POL" athleteid="2167">
              <RESULTS>
                <RESULT eventid="1102" points="557" swimtime="00:00:25.86" resultid="2168" heatid="4680" lane="1" entrytime="00:00:26.00" />
                <RESULT eventid="1255" points="584" swimtime="00:01:01.48" resultid="2169" heatid="4724" lane="2" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="621" swimtime="00:00:27.14" resultid="2170" heatid="4749" lane="3" entrytime="00:00:28.00" />
                <RESULT eventid="1491" points="476" swimtime="00:01:07.61" resultid="2171" heatid="4793" lane="2" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NESKAT" nation="POL" region="11" clubid="2213" name="NESSE Kozak Team Katowice">
          <ATHLETES>
            <ATHLETE firstname="Wojciech" lastname="Wodyński" birthdate="1977-03-01" gender="M" nation="POL" athleteid="2214">
              <RESULTS>
                <RESULT eventid="1102" points="300" swimtime="00:00:34.12" resultid="2215" heatid="4673" lane="3" entrytime="00:00:33.88" />
                <RESULT comment="K14 - Pływak wykonał kopnięcie nóg w płaszczyźnie pionowej w dół (z wyjątkiem jednego ruchu po starcie i nawrocie)." eventid="1171" status="DSQ" swimtime="00:00:42.32" resultid="2216" heatid="4698" lane="5" entrytime="00:00:41.15" />
                <RESULT eventid="1589" points="267" swimtime="00:01:36.67" resultid="2217" heatid="4771" lane="5" entrytime="00:01:31.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1519" points="222" swimtime="00:00:43.29" resultid="2218" heatid="4800" lane="3" entrytime="00:00:43.58" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KORKRA" nation="POL" region="06" clubid="2568" name="KORONA 1919 Kraków">
          <CONTACT city="Kraków" name="Mariola Kuliś" phone="500677133" state="MAŁOP" />
          <ATHLETES>
            <ATHLETE firstname="Bogusław" lastname="Kwiatkowski" birthdate="1956-07-24" gender="M" nation="POL" athleteid="2668">
              <RESULTS>
                <RESULT eventid="1102" points="158" swimtime="00:00:47.07" resultid="2669" heatid="4670" lane="4" entrytime="00:00:50.00" />
                <RESULT eventid="1199" points="124" swimtime="00:04:16.05" resultid="2670" heatid="4709" lane="3" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.95" />
                    <SPLIT distance="100" swimtime="00:01:58.80" />
                    <SPLIT distance="150" swimtime="00:03:09.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="131" swimtime="00:01:53.83" resultid="2671" heatid="4758" lane="5" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1519" points="130" swimtime="00:00:59.96" resultid="2672" heatid="4799" lane="2" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Leńczowska" birthdate="1982-01-15" gender="F" nation="POL" athleteid="2629">
              <RESULTS>
                <RESULT eventid="1059" points="538" swimtime="00:00:32.00" resultid="2630" heatid="4668" lane="6" entrytime="00:00:31.25" />
                <RESULT eventid="1129" points="477" swimtime="00:01:20.93" resultid="2631" heatid="4684" lane="3" entrytime="00:01:19.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="483" swimtime="00:01:12.77" resultid="2632" heatid="4754" lane="4" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1505" points="494" swimtime="00:00:36.52" resultid="2633" heatid="4797" lane="2" entrytime="00:00:36.45" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Mleczko" birthdate="1947-08-26" gender="M" nation="POL" athleteid="2579">
              <RESULTS>
                <RESULT eventid="1102" points="506" swimtime="00:00:36.02" resultid="2580" heatid="4672" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1199" points="395" swimtime="00:03:20.34" resultid="2581" heatid="4710" lane="2" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.41" />
                    <SPLIT distance="100" swimtime="00:01:40.89" />
                    <SPLIT distance="150" swimtime="00:02:31.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="401" swimtime="00:01:27.89" resultid="2582" heatid="4759" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="337" swimtime="00:07:32.58" resultid="2583" heatid="4808" lane="5" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.49" />
                    <SPLIT distance="100" swimtime="00:01:48.51" />
                    <SPLIT distance="150" swimtime="00:02:46.70" />
                    <SPLIT distance="200" swimtime="00:03:44.98" />
                    <SPLIT distance="250" swimtime="00:04:43.35" />
                    <SPLIT distance="300" swimtime="00:05:40.87" />
                    <SPLIT distance="350" swimtime="00:06:37.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Próchniewicz" birthdate="1978-02-18" gender="M" nation="POL" athleteid="2656">
              <RESULTS>
                <RESULT eventid="1102" points="208" swimtime="00:00:38.41" resultid="2657" heatid="4671" lane="5" entrytime="00:00:38.00" />
                <RESULT eventid="1491" points="124" swimtime="00:01:54.22" resultid="2658" heatid="4787" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1519" points="126" swimtime="00:00:50.76" resultid="2659" heatid="4800" lane="4" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Waga" birthdate="1940-07-04" gender="M" nation="POL" athleteid="2619">
              <RESULTS>
                <RESULT eventid="1199" points="197" swimtime="00:04:32.12" resultid="2620" heatid="4709" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.16" />
                    <SPLIT distance="100" swimtime="00:02:07.68" />
                    <SPLIT distance="150" swimtime="00:03:17.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1283" points="151" swimtime="00:06:17.81" resultid="2621" heatid="4730" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:30.84" />
                    <SPLIT distance="100" swimtime="00:03:08.71" />
                    <SPLIT distance="150" swimtime="00:04:46.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1589" points="153" swimtime="00:02:51.64" resultid="2622" heatid="4769" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:22.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="231" swimtime="00:09:12.86" resultid="2623" heatid="4807" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.57" />
                    <SPLIT distance="100" swimtime="00:02:15.46" />
                    <SPLIT distance="150" swimtime="00:03:27.34" />
                    <SPLIT distance="200" swimtime="00:04:38.94" />
                    <SPLIT distance="250" swimtime="00:05:49.47" />
                    <SPLIT distance="300" swimtime="00:06:58.94" />
                    <SPLIT distance="350" swimtime="00:08:07.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Weronika" lastname="Zygmuntowicz" birthdate="1982-10-17" gender="F" nation="POL" athleteid="2639">
              <RESULTS>
                <RESULT eventid="1059" points="480" swimtime="00:00:33.23" resultid="2640" heatid="4667" lane="3" entrytime="00:00:32.50" />
                <RESULT eventid="1213" points="377" swimtime="00:03:12.63" resultid="2641" heatid="4715" lane="5" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.35" />
                    <SPLIT distance="100" swimtime="00:01:27.61" />
                    <SPLIT distance="150" swimtime="00:02:25.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="444" swimtime="00:00:36.96" resultid="2642" heatid="4742" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1477" points="381" swimtime="00:01:28.52" resultid="2643" heatid="4785" lane="6" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Orlewicz-Musiał" birthdate="1960-05-29" gender="F" nation="POL" athleteid="2634">
              <RESULTS>
                <RESULT eventid="1059" points="178" swimtime="00:00:50.62" resultid="2635" heatid="4666" lane="6" entrytime="00:00:50.00" />
                <RESULT eventid="1213" points="171" swimtime="00:04:42.59" resultid="2636" heatid="4714" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.35" />
                    <SPLIT distance="100" swimtime="00:02:15.40" />
                    <SPLIT distance="150" swimtime="00:03:39.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="130" swimtime="00:01:01.60" resultid="2637" heatid="4741" lane="6" />
                <RESULT eventid="1477" points="155" swimtime="00:02:14.45" resultid="2638" heatid="4783" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Janeczko" birthdate="1972-12-23" gender="F" nation="POL" athleteid="2599">
              <RESULTS>
                <RESULT eventid="1185" status="DNS" swimtime="00:00:00.00" resultid="2600" heatid="4706" lane="3" entrytime="00:03:10.00" />
                <RESULT eventid="1241" status="DNS" swimtime="00:00:00.00" resultid="2601" heatid="4719" lane="1" entrytime="00:01:45.00" />
                <RESULT eventid="1358" status="DNS" swimtime="00:00:00.00" resultid="2602" heatid="4741" lane="3" entrytime="00:00:39.00" />
                <RESULT eventid="1505" status="DNS" swimtime="00:00:00.00" resultid="2603" heatid="4796" lane="3" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Pycia" birthdate="1966-03-21" gender="M" nation="POL" athleteid="2589">
              <RESULTS>
                <RESULT eventid="1102" points="497" swimtime="00:00:30.76" resultid="2590" heatid="4675" lane="4" entrytime="00:00:30.30" />
                <RESULT eventid="1171" points="394" swimtime="00:00:39.85" resultid="2591" heatid="4699" lane="3" entrytime="00:00:38.30" />
                <RESULT eventid="1407" points="492" swimtime="00:01:08.79" resultid="2592" heatid="4761" lane="2" entrytime="00:01:08.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="401" swimtime="00:01:23.12" resultid="2593" heatid="4790" lane="2" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariola" lastname="Kuliś" birthdate="1966-07-27" gender="F" nation="POL" athleteid="2569">
              <RESULTS>
                <RESULT eventid="1059" points="745" swimtime="00:00:30.67" resultid="2570" heatid="4668" lane="1" entrytime="00:00:30.87" />
                <RESULT eventid="1157" points="785" swimtime="00:00:38.11" resultid="2571" heatid="4693" lane="3" entrytime="00:00:38.20" />
                <RESULT eventid="1358" points="714" swimtime="00:00:32.88" resultid="2572" heatid="4742" lane="3" entrytime="00:00:33.65" />
                <RESULT eventid="1477" points="676" swimtime="00:01:18.72" resultid="2573" heatid="4785" lane="3" entrytime="00:01:17.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Borek" birthdate="1991-01-01" gender="M" nation="POL" athleteid="2609">
              <RESULTS>
                <RESULT eventid="1143" points="370" swimtime="00:01:13.25" resultid="2610" heatid="4689" lane="1" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="376" swimtime="00:00:37.03" resultid="2611" heatid="4700" lane="3" entrytime="00:00:36.00" />
                <RESULT eventid="1491" points="400" swimtime="00:01:12.33" resultid="2612" heatid="4791" lane="3" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1519" points="345" swimtime="00:00:34.01" resultid="2613" heatid="4802" lane="1" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulina" lastname="Bielańska" birthdate="1984-04-20" gender="F" nation="POL" athleteid="2624">
              <RESULTS>
                <RESULT eventid="1059" points="145" swimtime="00:00:47.75" resultid="2625" heatid="4664" lane="3" />
                <RESULT eventid="1269" points="137" swimtime="00:04:52.16" resultid="2626" heatid="4726" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.25" />
                    <SPLIT distance="100" swimtime="00:02:22.12" />
                    <SPLIT distance="150" swimtime="00:03:38.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1575" points="123" swimtime="00:02:18.99" resultid="2627" heatid="4765" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1505" points="133" swimtime="00:00:54.15" resultid="2628" heatid="4795" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Jawień" birthdate="1971-06-11" gender="M" nation="POL" athleteid="2673">
              <RESULTS>
                <RESULT eventid="1143" points="424" swimtime="00:01:17.13" resultid="2674" heatid="4688" lane="4" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1255" points="431" swimtime="00:01:15.18" resultid="2675" heatid="4722" lane="6" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1589" points="482" swimtime="00:01:22.01" resultid="2676" heatid="4772" lane="5" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1519" points="442" swimtime="00:00:35.05" resultid="2677" heatid="4802" lane="6" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Waldemar" lastname="Piszczek" birthdate="1962-11-10" gender="M" nation="POL" athleteid="2584">
              <RESULTS>
                <RESULT eventid="1102" points="568" swimtime="00:00:30.06" resultid="2585" heatid="4675" lane="5" entrytime="00:00:30.50" />
                <RESULT eventid="1171" points="627" swimtime="00:00:36.82" resultid="2586" heatid="4700" lane="5" entrytime="00:00:37.00" />
                <RESULT eventid="1379" points="607" swimtime="00:00:31.62" resultid="2587" heatid="4748" lane="1" entrytime="00:00:31.50" />
                <RESULT eventid="1519" points="566" swimtime="00:00:35.59" resultid="2588" heatid="4801" lane="2" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Damian" lastname="Jośko" birthdate="1994-07-25" gender="M" nation="POL" athleteid="2614">
              <RESULTS>
                <RESULT eventid="1102" points="425" swimtime="00:00:28.31" resultid="2615" heatid="4678" lane="6" entrytime="00:00:28.00" />
                <RESULT eventid="1171" points="409" swimtime="00:00:36.35" resultid="2616" heatid="4700" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="1379" points="323" swimtime="00:00:33.75" resultid="2617" heatid="4747" lane="4" entrytime="00:00:32.50" />
                <RESULT eventid="1589" points="313" swimtime="00:01:25.66" resultid="2618" heatid="4772" lane="2" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Macierzewska" birthdate="1960-04-20" gender="F" nation="POL" athleteid="2594">
              <RESULTS>
                <RESULT eventid="1185" points="499" swimtime="00:02:51.40" resultid="2595" heatid="4707" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.10" />
                    <SPLIT distance="100" swimtime="00:01:23.92" />
                    <SPLIT distance="150" swimtime="00:02:09.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1241" points="486" swimtime="00:01:30.93" resultid="2596" heatid="4719" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="502" swimtime="00:01:18.78" resultid="2597" heatid="4754" lane="5" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1449" points="469" swimtime="00:03:27.49" resultid="2598" heatid="4780" lane="3" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.23" />
                    <SPLIT distance="100" swimtime="00:01:36.39" />
                    <SPLIT distance="150" swimtime="00:02:33.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mirosław" lastname="Wożniak" birthdate="1969-08-22" gender="M" nation="POL" athleteid="2648">
              <RESULTS>
                <RESULT eventid="1227" points="422" swimtime="00:02:48.54" resultid="2649" heatid="4717" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.93" />
                    <SPLIT distance="100" swimtime="00:01:17.73" />
                    <SPLIT distance="150" swimtime="00:02:07.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="463" swimtime="00:01:14.56" resultid="2650" heatid="4791" lane="4" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Janusz" lastname="Toporski" birthdate="1959-10-20" gender="M" nation="POL" athleteid="2574">
              <RESULTS>
                <RESULT eventid="1255" points="173" swimtime="00:01:48.06" resultid="2575" heatid="4720" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1283" points="376" swimtime="00:03:31.00" resultid="2576" heatid="4731" lane="5" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.29" />
                    <SPLIT distance="100" swimtime="00:01:44.86" />
                    <SPLIT distance="150" swimtime="00:02:38.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1589" points="322" swimtime="00:01:41.42" resultid="2577" heatid="4770" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="195" swimtime="00:04:01.81" resultid="2578" heatid="4781" lane="1" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.58" />
                    <SPLIT distance="100" swimtime="00:01:58.21" />
                    <SPLIT distance="150" swimtime="00:03:00.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariusz" lastname="Baranik" birthdate="1969-06-29" gender="M" nation="POL" athleteid="2604">
              <RESULTS>
                <RESULT eventid="1102" points="667" swimtime="00:00:26.76" resultid="2605" heatid="4679" lane="2" entrytime="00:00:26.70" />
                <RESULT eventid="1171" points="593" swimtime="00:00:35.37" resultid="2606" heatid="4701" lane="4" entrytime="00:00:34.50" />
                <RESULT eventid="1379" points="665" swimtime="00:00:29.20" resultid="2607" heatid="4748" lane="4" entrytime="00:00:29.60" />
                <RESULT eventid="1491" points="559" swimtime="00:01:10.03" resultid="2608" heatid="4792" lane="5" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Liszkowski" birthdate="1972-07-17" gender="M" nation="POL" athleteid="2660">
              <RESULTS>
                <RESULT eventid="1171" points="453" swimtime="00:00:38.68" resultid="2661" heatid="4699" lane="4" entrytime="00:00:39.00" />
                <RESULT eventid="1519" points="423" swimtime="00:00:35.55" resultid="2662" heatid="4801" lane="4" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1350" points="545" swimtime="00:02:13.98" resultid="2679" heatid="4740" lane="1" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                    <SPLIT distance="100" swimtime="00:01:14.44" />
                    <SPLIT distance="150" swimtime="00:01:46.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2648" number="1" />
                    <RELAYPOSITION athleteid="2673" number="2" />
                    <RELAYPOSITION athleteid="2660" number="3" />
                    <RELAYPOSITION athleteid="2604" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1325" points="422" swimtime="00:04:36.62" resultid="2681" heatid="4737" lane="5" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                    <SPLIT distance="100" swimtime="00:01:10.16" />
                    <SPLIT distance="150" swimtime="00:01:41.54" />
                    <SPLIT distance="200" swimtime="00:02:17.00" />
                    <SPLIT distance="250" swimtime="00:02:50.27" />
                    <SPLIT distance="300" swimtime="00:03:26.63" />
                    <SPLIT distance="350" swimtime="00:03:59.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2614" number="1" />
                    <RELAYPOSITION athleteid="2648" number="2" />
                    <RELAYPOSITION athleteid="2589" number="3" />
                    <RELAYPOSITION athleteid="2673" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1350" points="239" swimtime="00:03:03.83" resultid="2680" heatid="4739" lane="2" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.52" />
                    <SPLIT distance="100" swimtime="00:01:49.08" />
                    <SPLIT distance="150" swimtime="00:02:27.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2668" number="1" />
                    <RELAYPOSITION athleteid="2574" number="2" />
                    <RELAYPOSITION athleteid="2589" number="3" />
                    <RELAYPOSITION athleteid="2579" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1329" points="552" swimtime="00:02:27.34" resultid="2678" heatid="4738" lane="4" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                    <SPLIT distance="100" swimtime="00:01:14.80" />
                    <SPLIT distance="150" swimtime="00:01:51.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2629" number="1" />
                    <RELAYPOSITION athleteid="2569" number="2" />
                    <RELAYPOSITION athleteid="2639" number="3" />
                    <RELAYPOSITION athleteid="2594" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SIEKRA" nation="POL" region="06" clubid="2805" name="Stowarzyszenie Siemacha Kraków">
          <CONTACT city="Kraków" email="pajka@poczta.onet.eu" name="Palmowska- Latuszek" phone="500044884" state="MAŁOP" />
          <ATHLETES>
            <ATHLETE firstname="Paulina" lastname="Palmowska- Latuszek" birthdate="1985-08-01" gender="F" nation="POL" license="503706600141" athleteid="2806">
              <RESULTS>
                <RESULT eventid="1129" points="515" swimtime="00:01:15.40" resultid="2807" heatid="4685" lane="1" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1185" points="538" swimtime="00:02:31.35" resultid="2808" heatid="4708" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.21" />
                    <SPLIT distance="100" swimtime="00:01:12.97" />
                    <SPLIT distance="150" swimtime="00:01:52.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1421" points="536" swimtime="00:02:44.14" resultid="2809" heatid="4776" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.77" />
                    <SPLIT distance="100" swimtime="00:01:19.94" />
                    <SPLIT distance="150" swimtime="00:02:02.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1533" points="511" swimtime="00:05:28.36" resultid="2810" heatid="4806" lane="1" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                    <SPLIT distance="100" swimtime="00:01:18.00" />
                    <SPLIT distance="150" swimtime="00:01:59.50" />
                    <SPLIT distance="200" swimtime="00:02:41.25" />
                    <SPLIT distance="250" swimtime="00:03:23.02" />
                    <SPLIT distance="300" swimtime="00:04:05.00" />
                    <SPLIT distance="350" swimtime="00:04:46.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DELTAR" nation="POL" region="08" clubid="2475" name="UKS Delfin Tarnobrzeg">
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Kunicki" birthdate="1972-03-14" gender="M" nation="POL" athleteid="2481">
              <RESULTS>
                <RESULT eventid="1102" points="442" swimtime="00:00:30.69" resultid="2482" heatid="4675" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1255" points="354" swimtime="00:01:20.25" resultid="2483" heatid="4721" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="434" swimtime="00:00:33.66" resultid="2484" heatid="4746" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1463" points="293" swimtime="00:03:14.52" resultid="2485" heatid="4781" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.51" />
                    <SPLIT distance="100" swimtime="00:01:33.98" />
                    <SPLIT distance="150" swimtime="00:02:24.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Tobiasz" birthdate="1979-02-01" gender="F" nation="POL" athleteid="2476">
              <RESULTS>
                <RESULT eventid="1059" points="282" swimtime="00:00:39.69" resultid="2477" heatid="4666" lane="1" entrytime="00:00:45.00" />
                <RESULT eventid="1241" points="176" swimtime="00:01:50.02" resultid="2478" heatid="4718" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="212" swimtime="00:00:47.29" resultid="2479" heatid="4741" lane="1" entrytime="00:00:47.00" />
                <RESULT eventid="1449" points="190" swimtime="00:04:04.64" resultid="2480" heatid="4780" lane="2" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.57" />
                    <SPLIT distance="100" swimtime="00:01:56.58" />
                    <SPLIT distance="150" swimtime="00:03:00.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DWOCZE" nation="POL" region="11" clubid="3056" name="UKS Dwójeczka Częstochowa">
          <CONTACT city="Częstochowa" email="klub.uks.2@wp.pl" name="Maciejewski" phone="668306689" state="ŚLĄS" street="Baczyńskiego 2a" zip="42-224" />
          <ATHLETES>
            <ATHLETE firstname="Ireneusz" lastname="Stachurski" birthdate="1969-07-22" gender="M" nation="POL" license="107311700001" athleteid="3057">
              <RESULTS>
                <RESULT eventid="1199" points="295" swimtime="00:02:52.20" resultid="3058" heatid="4711" lane="6" entrytime="00:02:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.61" />
                    <SPLIT distance="100" swimtime="00:01:21.05" />
                    <SPLIT distance="150" swimtime="00:02:06.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1255" points="164" swimtime="00:01:43.68" resultid="3059" heatid="4721" lane="6" entrytime="00:01:41.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="285" swimtime="00:01:18.23" resultid="3060" heatid="4760" lane="6" entrytime="00:01:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="257" swimtime="00:06:24.59" resultid="3061" heatid="4807" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.75" />
                    <SPLIT distance="100" swimtime="00:01:27.15" />
                    <SPLIT distance="150" swimtime="00:02:17.24" />
                    <SPLIT distance="200" swimtime="00:03:07.70" />
                    <SPLIT distance="250" swimtime="00:03:58.74" />
                    <SPLIT distance="300" swimtime="00:04:49.63" />
                    <SPLIT distance="350" swimtime="00:05:39.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOTSTA" nation="POL" region="08" clubid="2330" name="MOTYL MOSIR Stalowa Wola">
          <CONTACT city="Stalowa Wola" email="petecka.m@gmail.com" name="Petecka" phone="602829589" street="al. Jana Pawła II 13/59" zip="37-450" />
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Petecka" birthdate="1967-04-17" gender="F" nation="POL" license="100908600388" athleteid="2336">
              <RESULTS>
                <RESULT eventid="1059" points="454" swimtime="00:00:36.18" resultid="2337" heatid="4666" lane="2" entrytime="00:00:38.99" />
                <RESULT eventid="1157" points="392" swimtime="00:00:48.01" resultid="2338" heatid="4692" lane="4" entrytime="00:00:47.99" />
                <RESULT eventid="1575" points="423" swimtime="00:01:43.02" resultid="2339" heatid="4767" lane="6" entrytime="00:01:41.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1477" points="427" swimtime="00:01:31.71" resultid="2340" heatid="4784" lane="4" entrytime="00:01:29.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arkadiusz" lastname="Berwecki" birthdate="1973-01-14" gender="M" nation="POL" license="100908700263" athleteid="2331">
              <RESULTS>
                <RESULT eventid="1171" points="595" swimtime="00:00:34.07" resultid="2332" heatid="4696" lane="4" entrytime="00:00:49.99" />
                <RESULT eventid="1255" points="682" swimtime="00:01:02.56" resultid="2333" heatid="4724" lane="6" entrytime="00:01:01.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="644" swimtime="00:00:28.23" resultid="2334" heatid="4750" lane="6" entrytime="00:00:27.79" />
                <RESULT eventid="1491" points="674" swimtime="00:01:05.79" resultid="2335" heatid="4794" lane="6" entrytime="00:01:04.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WETZAB" nation="POL" region="11" clubid="3507" name="WETERAN Zabrze">
          <CONTACT city="Zabrze" email="weteranzabrze.prv.pl" name="BOSOWSKI  WŁODZIMIERZ" state="ŚLĄSK" street="ŚW.JANA  4A/4" zip="41-803" />
          <ATHLETES>
            <ATHLETE firstname="Włodzimierz" lastname="Bosowski" birthdate="1948-05-22" gender="M" nation="POL" license="102611700014" athleteid="3535">
              <RESULTS>
                <RESULT eventid="1102" points="162" swimtime="00:00:49.35" resultid="3536" heatid="4671" lane="6" entrytime="00:00:39.50" />
                <RESULT eventid="1519" points="96" swimtime="00:01:12.28" resultid="3537" heatid="4800" lane="1" entrytime="00:00:47.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiesław" lastname="Kornicki" birthdate="1949-01-28" gender="M" nation="POL" license="102611700015" athleteid="3526">
              <RESULTS>
                <RESULT eventid="1102" points="504" swimtime="00:00:33.78" resultid="3527" heatid="4673" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="1379" points="426" swimtime="00:00:39.24" resultid="3528" heatid="4745" lane="5" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Fecica" birthdate="1940-11-29" gender="M" nation="POL" license="102611700018" athleteid="3529">
              <RESULTS>
                <RESULT eventid="1283" points="580" swimtime="00:04:01.41" resultid="3530" heatid="4731" lane="2" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.23" />
                    <SPLIT distance="100" swimtime="00:01:55.47" />
                    <SPLIT distance="150" swimtime="00:02:59.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1589" points="535" swimtime="00:01:53.06" resultid="3531" heatid="4770" lane="5" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beata" lastname="Sulewska" birthdate="1972-11-02" gender="F" nation="POL" license="102611600016" athleteid="3538">
              <RESULTS>
                <RESULT eventid="1185" points="659" swimtime="00:02:30.24" resultid="3539" heatid="4708" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                    <SPLIT distance="100" swimtime="00:01:13.56" />
                    <SPLIT distance="150" swimtime="00:01:52.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1269" status="DNS" swimtime="00:00:00.00" resultid="3540" heatid="4729" lane="6" entrytime="00:03:07.00" />
                <RESULT eventid="1393" points="583" swimtime="00:01:10.13" resultid="3541" heatid="4755" lane="6" entrytime="00:01:09.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1533" points="621" swimtime="00:05:21.06" resultid="3542" heatid="4806" lane="5" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.52" />
                    <SPLIT distance="100" swimtime="00:01:17.33" />
                    <SPLIT distance="150" swimtime="00:01:57.72" />
                    <SPLIT distance="200" swimtime="00:02:38.76" />
                    <SPLIT distance="250" swimtime="00:03:19.83" />
                    <SPLIT distance="300" swimtime="00:04:00.79" />
                    <SPLIT distance="350" swimtime="00:04:42.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Twardysko" birthdate="1956-01-16" gender="M" nation="POL" license="502011603019" athleteid="3512">
              <RESULTS>
                <RESULT comment="O1 - Pływak wystartował po komendzie na miejsca i zajęciu pozycji nieruchomej, a przed sygnałem startu." eventid="1143" status="DSQ" swimtime="00:01:33.56" resultid="3513" heatid="4687" lane="5" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1199" points="376" swimtime="00:02:56.70" resultid="3514" heatid="4710" lane="4" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                    <SPLIT distance="100" swimtime="00:01:20.42" />
                    <SPLIT distance="150" swimtime="00:02:06.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="393" swimtime="00:01:18.91" resultid="3515" heatid="4759" lane="4" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="357" swimtime="00:06:17.80" resultid="3516" heatid="4808" lane="3" entrytime="00:06:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.69" />
                    <SPLIT distance="100" swimtime="00:01:25.81" />
                    <SPLIT distance="150" swimtime="00:02:13.34" />
                    <SPLIT distance="200" swimtime="00:03:02.24" />
                    <SPLIT distance="250" swimtime="00:03:51.83" />
                    <SPLIT distance="300" swimtime="00:04:41.45" />
                    <SPLIT distance="350" swimtime="00:05:31.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krystyna" lastname="Fecica" birthdate="1943-03-12" gender="F" nation="POL" license="102611600019" athleteid="3532">
              <RESULTS>
                <RESULT eventid="1241" points="409" swimtime="00:02:01.33" resultid="3533" heatid="4718" lane="4" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1575" points="457" swimtime="00:02:05.25" resultid="3534" heatid="4766" lane="5" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Teresa" lastname="Żylińska" birthdate="1950-10-13" gender="F" nation="POL" license="102611600029" athleteid="3517">
              <RESULTS>
                <RESULT eventid="1059" points="232" swimtime="00:00:52.69" resultid="3518" heatid="4665" lane="2" entrytime="00:00:52.50" />
                <RESULT eventid="1129" points="178" swimtime="00:02:16.15" resultid="3519" heatid="4683" lane="2" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="197" swimtime="00:02:00.76" resultid="3520" heatid="4752" lane="5" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1505" points="180" swimtime="00:01:02.28" resultid="3521" heatid="4796" lane="6" entrytime="00:01:02.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernard" lastname="Poloczek" birthdate="1947-02-25" gender="M" nation="POL" license="102611700032" athleteid="3508">
              <RESULTS>
                <RESULT eventid="1143" points="379" swimtime="00:01:42.34" resultid="3509" heatid="4687" lane="2" entrytime="00:01:40.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="371" swimtime="00:00:44.67" resultid="3510" heatid="4744" lane="1" entrytime="00:00:43.52" />
                <RESULT eventid="1519" points="435" swimtime="00:00:44.69" resultid="3511" heatid="4800" lane="2" entrytime="00:00:45.67" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Genowefa" lastname="Drużyńska" birthdate="1951-02-18" gender="F" nation="POL" license="102611600033" athleteid="3522">
              <RESULTS>
                <RESULT eventid="1157" points="308" swimtime="00:01:03.38" resultid="3523" heatid="4691" lane="2" entrytime="00:01:05.00" />
                <RESULT eventid="1269" points="228" swimtime="00:05:34.65" resultid="3524" heatid="4726" lane="4" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.22" />
                    <SPLIT distance="100" swimtime="00:02:41.84" />
                    <SPLIT distance="150" swimtime="00:04:09.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1575" points="207" swimtime="00:02:38.76" resultid="3525" heatid="4765" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="280" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1350" swimtime="00:03:04.11" resultid="3543" heatid="4739" lane="4" entrytime="00:02:57.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.37" />
                    <SPLIT distance="100" swimtime="00:01:32.55" />
                    <SPLIT distance="150" swimtime="00:02:14.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3512" number="1" />
                    <RELAYPOSITION athleteid="3529" number="2" />
                    <RELAYPOSITION athleteid="3526" number="3" />
                    <RELAYPOSITION athleteid="3535" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="TEAKRA" nation="POL" region="06" clubid="2411" name="JK TEAM Kraków">
          <CONTACT city="Kraków" name="Joanna Kwatera" phone="790611187" state="MAŁOP" />
          <ATHLETES>
            <ATHLETE firstname="Ryszard" lastname="Zając" birthdate="1984-01-01" gender="M" nation="POL" athleteid="2424">
              <RESULTS>
                <RESULT eventid="1102" points="220" swimtime="00:00:35.68" resultid="2425" heatid="4672" lane="3" entrytime="00:00:34.50" />
                <RESULT eventid="1255" points="106" swimtime="00:01:51.38" resultid="2426" heatid="4720" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="215" swimtime="00:01:19.60" resultid="2427" heatid="4759" lane="2" entrytime="00:01:19.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="174" swimtime="00:01:38.34" resultid="2428" heatid="4788" lane="2" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agata" lastname="Jasik" birthdate="1984-01-01" gender="F" nation="POL" athleteid="2412">
              <RESULTS>
                <RESULT eventid="1185" points="301" swimtime="00:03:03.63" resultid="2413" heatid="4707" lane="5" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.67" />
                    <SPLIT distance="100" swimtime="00:01:25.72" />
                    <SPLIT distance="150" swimtime="00:02:14.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="331" swimtime="00:01:19.47" resultid="2414" heatid="4754" lane="6" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1533" points="296" swimtime="00:06:33.95" resultid="2415" heatid="4804" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                    <SPLIT distance="100" swimtime="00:01:28.11" />
                    <SPLIT distance="150" swimtime="00:02:17.41" />
                    <SPLIT distance="200" swimtime="00:03:08.43" />
                    <SPLIT distance="250" swimtime="00:04:00.20" />
                    <SPLIT distance="300" swimtime="00:04:51.80" />
                    <SPLIT distance="350" swimtime="00:05:44.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Wolak" birthdate="1987-01-01" gender="M" nation="POL" athleteid="2429">
              <RESULTS>
                <RESULT eventid="1102" points="468" swimtime="00:00:27.73" resultid="2430" heatid="4678" lane="4" entrytime="00:00:27.50" />
                <RESULT eventid="1255" points="392" swimtime="00:01:12.09" resultid="2431" heatid="4720" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="448" swimtime="00:00:30.21" resultid="2432" heatid="4748" lane="5" entrytime="00:00:31.50" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="2433" heatid="4787" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Jania" birthdate="1988-01-01" gender="M" nation="POL" athleteid="2416">
              <RESULTS>
                <RESULT eventid="1102" points="216" swimtime="00:00:35.87" resultid="2417" heatid="4673" lane="4" entrytime="00:00:34.00" />
                <RESULT eventid="1227" points="186" swimtime="00:03:24.88" resultid="2418" heatid="4716" lane="2" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.82" />
                    <SPLIT distance="100" swimtime="00:01:37.99" />
                    <SPLIT distance="150" swimtime="00:02:35.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="184" swimtime="00:00:40.23" resultid="2419" heatid="4745" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="1589" points="213" swimtime="00:01:39.00" resultid="2420" heatid="4771" lane="6" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karol" lastname="Głowacz" birthdate="1997-01-01" gender="M" nation="POL" athleteid="2434">
              <RESULTS>
                <RESULT eventid="1102" points="385" swimtime="00:00:29.24" resultid="2435" heatid="4677" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="1171" points="430" swimtime="00:00:35.75" resultid="2436" heatid="4701" lane="3" entrytime="00:00:34.00" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="2437" heatid="4791" lane="6" entrytime="00:01:18.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Hełpa" birthdate="1990-01-01" gender="M" nation="POL" athleteid="2421">
              <RESULTS>
                <RESULT eventid="1102" points="376" swimtime="00:00:29.84" resultid="2422" heatid="4677" lane="2" entrytime="00:00:29.00" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="2423" heatid="4791" lane="1" entrytime="00:01:15.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1350" points="322" swimtime="00:02:23.62" resultid="2438" heatid="4740" lane="6" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.71" />
                    <SPLIT distance="100" swimtime="00:01:13.58" />
                    <SPLIT distance="150" swimtime="00:01:55.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2421" number="1" />
                    <RELAYPOSITION athleteid="2434" number="2" />
                    <RELAYPOSITION athleteid="2424" number="3" />
                    <RELAYPOSITION athleteid="2429" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1325" points="395" swimtime="00:04:37.31" resultid="2439" heatid="4736" lane="4" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.42" />
                    <SPLIT distance="100" swimtime="00:01:07.15" />
                    <SPLIT distance="150" swimtime="00:01:38.09" />
                    <SPLIT distance="200" swimtime="00:02:13.41" />
                    <SPLIT distance="250" swimtime="00:02:51.32" />
                    <SPLIT distance="300" swimtime="00:03:34.52" />
                    <SPLIT distance="350" swimtime="00:04:04.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2434" number="1" />
                    <RELAYPOSITION athleteid="2421" number="2" />
                    <RELAYPOSITION athleteid="2424" number="3" />
                    <RELAYPOSITION athleteid="2429" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MOOST" nation="POL" region="12" clubid="2172" name="MOSiR Ostrowiec Świętokrzyski">
          <CONTACT city="Ostrowiec Świętokrzyski" email="basen@mosir.ostrowiec.pl" name="Różalski Józef" phone="510-600-865" state="ŚWIĘT" />
          <ATHLETES>
            <ATHLETE firstname="Józef" lastname="Różalski" birthdate="1945-03-28" gender="M" nation="POL" license="501012700001" athleteid="2173">
              <RESULTS>
                <RESULT eventid="1102" points="505" swimtime="00:00:36.04" resultid="2174" heatid="4671" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1379" points="407" swimtime="00:00:43.29" resultid="2176" heatid="4744" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1491" points="377" swimtime="00:01:47.42" resultid="2177" heatid="4788" lane="5" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="428" swimtime="00:00:50.89" resultid="3130" heatid="4696" lane="2" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIERUD" nation="POL" region="11" clubid="2811" name="Zawodnik Niezrzeszony Ruda Śląska" shortname="Zawodnik Niezrzeszony Ruda Ślą">
          <ATHLETES>
            <ATHLETE firstname="Adam" lastname="Miler" birthdate="2002-11-13" gender="M" nation="POL" athleteid="2812">
              <RESULTS>
                <RESULT eventid="1379" swimtime="00:00:34.78" resultid="2813" heatid="4746" lane="5" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KAPZDZ" nation="POL" region="07" clubid="3582" name="Grupa KAPIJA Sport Zdzieszowice" shortname="Grupa KAPIJA Sport Zdzieszowic">
          <CONTACT city="Zdzieszowice" email="dejot.swim@gmai.com" name="Dawid" phone="505127695" state="OPOLS" street="Jajuga" zip="47-330" />
          <ATHLETES>
            <ATHLETE firstname="Katarzyna" lastname="Gniot" birthdate="1980-09-23" gender="F" nation="POL" athleteid="3583">
              <RESULTS>
                <RESULT eventid="1129" status="DNS" swimtime="00:00:00.00" resultid="3584" heatid="4683" lane="3" entrytime="00:02:00.00" />
                <RESULT eventid="1185" status="DNS" swimtime="00:00:00.00" resultid="3585" heatid="4706" lane="1" entrytime="00:03:40.00" />
                <RESULT eventid="1393" status="DNS" swimtime="00:00:00.00" resultid="3586" heatid="4753" lane="6" entrytime="00:01:40.00" />
                <RESULT eventid="1421" status="DNS" swimtime="00:00:00.00" resultid="3587" heatid="4776" lane="6" entrytime="00:03:50.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06711" nation="POL" region="11" clubid="2348" name="UKS DRAGON Będzin">
          <CONTACT city="Będzin" name="Kot Marek" state="ŚLĄSK" />
          <ATHLETES>
            <ATHLETE firstname="Emil" lastname="Strumiński" birthdate="1988-05-18" gender="M" nation="POL" license="306711700032" athleteid="2349">
              <RESULTS>
                <RESULT eventid="1199" points="617" swimtime="00:02:04.67" resultid="2350" heatid="4713" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.27" />
                    <SPLIT distance="100" swimtime="00:01:00.92" />
                    <SPLIT distance="150" swimtime="00:01:33.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1255" points="579" swimtime="00:01:02.91" resultid="2351" heatid="4724" lane="5" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="586" swimtime="00:00:56.52" resultid="2352" heatid="4764" lane="6" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="567" swimtime="00:04:40.27" resultid="2353" heatid="4810" lane="2" entrytime="00:04:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.39" />
                    <SPLIT distance="100" swimtime="00:01:06.08" />
                    <SPLIT distance="150" swimtime="00:01:42.14" />
                    <SPLIT distance="200" swimtime="00:02:18.61" />
                    <SPLIT distance="250" swimtime="00:02:55.37" />
                    <SPLIT distance="300" swimtime="00:03:31.32" />
                    <SPLIT distance="350" swimtime="00:04:07.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MASGDY" nation="POL" region="10" clubid="2448" name="Gdynia Masters">
          <CONTACT city="Gdynia" email="kasiiamysiak@gmail.com" name="Mysiak" />
          <ATHLETES>
            <ATHLETE firstname="Zuzanna" lastname="Drążkiewicz" birthdate="1961-01-01" gender="F" nation="POL" athleteid="2449">
              <RESULTS>
                <RESULT eventid="1129" points="71" swimtime="00:02:54.92" resultid="2450" heatid="4683" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1185" points="78" swimtime="00:05:17.57" resultid="2451" heatid="4705" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.01" />
                    <SPLIT distance="100" swimtime="00:02:32.70" />
                    <SPLIT distance="150" swimtime="00:03:56.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Skwarło" birthdate="1939-01-01" gender="M" nation="POL" athleteid="2452">
              <RESULTS>
                <RESULT eventid="1283" points="289" swimtime="00:05:04.58" resultid="2454" heatid="4731" lane="1" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.29" />
                    <SPLIT distance="100" swimtime="00:02:27.68" />
                    <SPLIT distance="150" swimtime="00:03:49.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1589" points="281" swimtime="00:02:20.11" resultid="2455" heatid="4770" lane="6" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="201" swimtime="00:02:24.53" resultid="2456" heatid="4788" lane="6" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="397" swimtime="00:00:56.37" resultid="3834" heatid="4696" lane="5" entrytime="00:00:56.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SWIUKR" nation="UKR" clubid="3589" name="Ukraine Swim Team">
          <ATHLETES>
            <ATHLETE firstname="Iryna" lastname="Oriekhova" birthdate="1988-05-19" gender="F" nation="UKR" athleteid="3591">
              <RESULTS>
                <RESULT eventid="1213" points="301" swimtime="00:03:18.96" resultid="3650" heatid="4714" lane="3" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.07" />
                    <SPLIT distance="100" swimtime="00:01:36.29" />
                    <SPLIT distance="150" swimtime="00:02:31.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1575" points="272" swimtime="00:01:43.41" resultid="3651" heatid="4766" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1477" points="297" swimtime="00:01:33.66" resultid="3652" heatid="4784" lane="5" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yevgeniya" lastname="Motrych " birthdate="1983-11-07" gender="F" nation="UKR" athleteid="3593">
              <RESULTS>
                <RESULT eventid="1157" points="289" swimtime="00:00:47.87" resultid="3656" heatid="4692" lane="3" entrytime="00:00:45.00" />
                <RESULT eventid="1575" points="283" swimtime="00:01:45.17" resultid="3657" heatid="4767" lane="5" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1533" points="244" swimtime="00:07:00.15" resultid="3658" heatid="4805" lane="6" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.06" />
                    <SPLIT distance="100" swimtime="00:01:34.70" />
                    <SPLIT distance="150" swimtime="00:02:28.14" />
                    <SPLIT distance="200" swimtime="00:03:22.45" />
                    <SPLIT distance="250" swimtime="00:04:17.15" />
                    <SPLIT distance="300" swimtime="00:05:12.89" />
                    <SPLIT distance="350" swimtime="00:06:07.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tatsiana" lastname.en="Turtsevich" birthdate="1974-06-22" gender="F" nameprefix="Turtsevich" nation="UKR" athleteid="3590">
              <RESULTS>
                <RESULT eventid="1213" points="418" swimtime="00:03:09.25" resultid="3647" heatid="4715" lane="1" entrytime="00:03:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.39" />
                    <SPLIT distance="100" swimtime="00:01:28.31" />
                    <SPLIT distance="150" swimtime="00:02:26.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1477" points="438" swimtime="00:01:26.42" resultid="3648" heatid="4784" lane="3" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="446" swimtime="00:00:37.33" resultid="3649" heatid="4741" lane="2" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nataliia" lastname="Boryshkevych" birthdate="1976-04-15" gender="F" nation="UKR" athleteid="3594">
              <RESULTS>
                <RESULT eventid="1185" points="584" swimtime="00:02:30.68" resultid="3659" heatid="4708" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.91" />
                    <SPLIT distance="100" swimtime="00:01:13.16" />
                    <SPLIT distance="150" swimtime="00:01:52.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1241" points="369" swimtime="00:01:28.48" resultid="3660" heatid="4719" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="583" swimtime="00:01:09.28" resultid="3661" heatid="4754" lane="3" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valeriia" lastname="Khokhol" birthdate="1996-08-21" gender="F" nation="UKR" athleteid="3592">
              <RESULTS>
                <RESULT eventid="1269" status="DNS" swimtime="00:00:00.00" resultid="3653" heatid="4728" lane="2" entrytime="00:03:10.00" />
                <RESULT eventid="1575" status="DNS" swimtime="00:00:00.00" resultid="3654" heatid="4767" lane="2" entrytime="00:01:30.00" />
                <RESULT eventid="1533" points="176" swimtime="00:07:36.74" resultid="3655" heatid="4805" lane="2" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.27" />
                    <SPLIT distance="100" swimtime="00:01:45.22" />
                    <SPLIT distance="150" swimtime="00:02:44.05" />
                    <SPLIT distance="200" swimtime="00:03:43.62" />
                    <SPLIT distance="250" swimtime="00:04:42.56" />
                    <SPLIT distance="300" swimtime="00:05:41.74" />
                    <SPLIT distance="350" swimtime="00:06:40.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1088" points="455" swimtime="00:05:16.29" resultid="3662" heatid="4735" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                    <SPLIT distance="100" swimtime="00:01:14.81" />
                    <SPLIT distance="150" swimtime="00:01:55.79" />
                    <SPLIT distance="200" swimtime="00:02:37.57" />
                    <SPLIT distance="250" swimtime="00:03:18.35" />
                    <SPLIT distance="300" swimtime="00:04:05.68" />
                    <SPLIT distance="350" swimtime="00:04:38.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3590" number="1" />
                    <RELAYPOSITION athleteid="3591" number="2" />
                    <RELAYPOSITION athleteid="3593" number="3" />
                    <RELAYPOSITION athleteid="3594" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1329" points="373" swimtime="00:02:42.08" resultid="3663" heatid="4738" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.29" />
                    <SPLIT distance="100" swimtime="00:01:29.77" />
                    <SPLIT distance="150" swimtime="00:02:09.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3590" number="1" />
                    <RELAYPOSITION athleteid="3591" number="2" />
                    <RELAYPOSITION athleteid="3592" number="3" />
                    <RELAYPOSITION athleteid="3594" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="NIEGLO" nation="POL" region="01" clubid="2161" name="Zawodnik Niezrzeszony Głogów">
          <ATHLETES>
            <ATHLETE firstname="Rafał" lastname="Szklarzewski" birthdate="1985-05-06" gender="M" nation="POL" athleteid="2160">
              <RESULTS>
                <RESULT eventid="1102" status="DNS" swimtime="00:00:00.00" resultid="2162" heatid="4680" lane="5" entrytime="00:00:26.00" />
                <RESULT eventid="1407" status="DNS" swimtime="00:00:00.00" resultid="2163" heatid="4763" lane="5" entrytime="00:00:59.00" />
                <RESULT eventid="1199" status="DNS" swimtime="00:00:00.00" resultid="2164" heatid="4712" lane="1" entrytime="00:02:30.00" />
                <RESULT eventid="1379" status="DNS" swimtime="00:00:00.00" resultid="2165" heatid="4749" lane="5" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02607" nation="POL" region="06" clubid="2799" name="UKS JASIEŃ Sucha Beskidzka">
          <CONTACT city="Sucha Beskidzka" name="Miklusiak" phone="668803392" state="MAŁOP" />
          <ATHLETES>
            <ATHLETE firstname="Sabina" lastname="Sikora" birthdate="1984-10-03" gender="F" nation="POL" license="102706600159" athleteid="2800">
              <RESULTS>
                <RESULT eventid="1157" points="637" swimtime="00:00:36.80" resultid="2801" heatid="4694" lane="2" entrytime="00:00:36.40" />
                <RESULT eventid="1269" points="523" swimtime="00:03:07.00" resultid="2802" heatid="4728" lane="3" entrytime="00:03:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.66" />
                    <SPLIT distance="100" swimtime="00:01:30.23" />
                    <SPLIT distance="150" swimtime="00:02:19.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1575" points="512" swimtime="00:01:26.35" resultid="2803" heatid="4768" lane="2" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1477" points="540" swimtime="00:01:17.57" resultid="2804" heatid="4783" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIEPAW" nation="POL" region="11" clubid="2318" name="Zawodnik Niezrzeszony Pawłowice" shortname="Zawodnik Niezrzeszony Pawłowic">
          <ATHLETES>
            <ATHLETE firstname="Alicja" lastname="Gruca" birthdate="2000-12-14" gender="F" nation="POL" athleteid="2319">
              <RESULTS>
                <RESULT eventid="1269" swimtime="00:02:58.99" resultid="2320" heatid="4728" lane="1" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.91" />
                    <SPLIT distance="100" swimtime="00:01:24.93" />
                    <SPLIT distance="150" swimtime="00:02:11.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1575" swimtime="00:01:23.28" resultid="2322" heatid="4768" lane="1" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1477" swimtime="00:01:16.33" resultid="2323" heatid="4785" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" swimtime="00:00:38.66" resultid="2341" heatid="4693" lane="5" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAKWAR" nation="POL" region="14" clubid="3030" name="Klub Sportowy MAKO Warszawa">
          <CONTACT city="Warszawa" email="ania.plywanie@gmail.com" name="Anna Dąbrowska" phone="601 480 280" state="MAZOW" />
          <ATHLETES>
            <ATHLETE firstname="Timea" lastname="Balajcza" birthdate="1971-09-22" gender="F" nation="POL" athleteid="3031">
              <RESULTS>
                <RESULT eventid="1157" points="691" swimtime="00:00:38.42" resultid="3032" heatid="4694" lane="6" entrytime="00:00:38.11" />
                <RESULT eventid="1269" points="713" swimtime="00:03:06.04" resultid="3033" heatid="4729" lane="5" entrytime="00:03:04.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.73" />
                    <SPLIT distance="100" swimtime="00:01:28.19" />
                    <SPLIT distance="150" swimtime="00:02:16.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1575" points="665" swimtime="00:01:25.95" resultid="3034" heatid="4768" lane="5" entrytime="00:01:23.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1533" points="531" swimtime="00:05:38.19" resultid="3035" heatid="4805" lane="3" entrytime="00:05:38.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.09" />
                    <SPLIT distance="100" swimtime="00:01:20.01" />
                    <SPLIT distance="150" swimtime="00:02:03.10" />
                    <SPLIT distance="200" swimtime="00:02:46.27" />
                    <SPLIT distance="250" swimtime="00:03:29.15" />
                    <SPLIT distance="300" swimtime="00:04:12.62" />
                    <SPLIT distance="350" swimtime="00:04:55.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Rudziński" birthdate="1966-05-10" gender="M" nation="POL" athleteid="3036">
              <RESULTS>
                <RESULT eventid="1171" points="290" swimtime="00:00:44.17" resultid="3037" heatid="4697" lane="2" entrytime="00:00:43.87" />
                <RESULT eventid="1283" points="300" swimtime="00:03:33.42" resultid="3038" heatid="4732" lane="6" entrytime="00:03:27.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.54" />
                    <SPLIT distance="100" swimtime="00:01:39.67" />
                    <SPLIT distance="150" swimtime="00:02:36.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="190" swimtime="00:03:56.69" resultid="3039" heatid="4781" lane="5" entrytime="00:03:47.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.15" />
                    <SPLIT distance="100" swimtime="00:01:48.55" />
                    <SPLIT distance="150" swimtime="00:02:54.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Piórkowski" birthdate="1965-07-28" gender="M" nation="POL" athleteid="3045">
              <RESULTS>
                <RESULT eventid="1143" points="188" swimtime="00:01:46.19" resultid="3046" heatid="4687" lane="1" entrytime="00:01:50.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1199" points="155" swimtime="00:03:41.68" resultid="3047" heatid="4710" lane="6" entrytime="00:03:37.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.16" />
                    <SPLIT distance="100" swimtime="00:01:38.40" />
                    <SPLIT distance="150" swimtime="00:02:39.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1435" points="194" swimtime="00:03:54.01" resultid="3048" heatid="4778" lane="6" entrytime="00:03:53.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.13" />
                    <SPLIT distance="100" swimtime="00:01:54.38" />
                    <SPLIT distance="150" swimtime="00:02:53.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1519" points="160" swimtime="00:00:51.29" resultid="3049" heatid="4800" lane="6" entrytime="00:00:48.22" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Adamowicz" birthdate="1967-07-11" gender="M" nation="POL" athleteid="3040">
              <RESULTS>
                <RESULT eventid="1102" points="286" swimtime="00:00:37.00" resultid="3041" heatid="4672" lane="6" entrytime="00:00:37.06" />
                <RESULT eventid="1171" points="294" swimtime="00:00:43.94" resultid="3042" heatid="4698" lane="1" entrytime="00:00:42.88" />
                <RESULT eventid="1589" points="247" swimtime="00:01:42.42" resultid="3043" heatid="4770" lane="4" entrytime="00:01:41.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="178" swimtime="00:01:48.86" resultid="3044" heatid="4788" lane="1" entrytime="00:01:50.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00115" nation="POL" region="15" clubid="3307" name="KS Warta Poznań">
          <CONTACT city="Poznań" email="marcin@infopomoc.pl" name="Szymkowiak, Marcin" phone="691470291" state="WIELK" street="Droga Dębińska 12" zip="61-555" />
          <ATHLETES>
            <ATHLETE firstname="Przemysław" lastname="Waraczewski" birthdate="1962-04-19" gender="M" nation="POL" license="100115700344" athleteid="3323">
              <RESULTS>
                <RESULT eventid="1171" points="483" swimtime="00:00:40.17" resultid="3324" heatid="4698" lane="4" entrytime="00:00:41.00" entrycourse="SCM" />
                <RESULT eventid="1283" points="493" swimtime="00:03:12.86" resultid="3325" heatid="4732" lane="5" entrytime="00:03:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.90" />
                    <SPLIT distance="100" swimtime="00:01:30.80" />
                    <SPLIT distance="150" swimtime="00:02:21.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1589" points="485" swimtime="00:01:28.51" resultid="3326" heatid="4772" lane="6" entrytime="00:01:28.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="430" swimtime="00:01:25.07" resultid="3327" heatid="4790" lane="6" entrytime="00:01:24.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Osik" birthdate="1976-01-02" gender="M" nation="POL" license="500115700521" athleteid="3337">
              <RESULTS>
                <RESULT eventid="1143" points="539" swimtime="00:01:10.03" resultid="3338" heatid="4689" lane="4" entrytime="00:01:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1199" points="558" swimtime="00:02:17.11" resultid="3339" heatid="4713" lane="6" entrytime="00:02:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.07" />
                    <SPLIT distance="100" swimtime="00:01:05.32" />
                    <SPLIT distance="150" swimtime="00:01:41.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1435" points="452" swimtime="00:02:43.55" resultid="3340" heatid="4779" lane="6" entrytime="00:02:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                    <SPLIT distance="100" swimtime="00:01:16.11" />
                    <SPLIT distance="150" swimtime="00:01:59.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1519" points="495" swimtime="00:00:33.15" resultid="3341" heatid="4802" lane="2" entrytime="00:00:32.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Witt" birthdate="1991-08-11" gender="M" nation="POL" license="500115700645" athleteid="3318">
              <RESULTS>
                <RESULT eventid="1102" points="612" swimtime="00:00:25.36" resultid="3319" heatid="4682" lane="6" entrytime="00:00:24.34" entrycourse="SCM" />
                <RESULT eventid="1199" points="562" swimtime="00:02:08.57" resultid="3320" heatid="4713" lane="5" entrytime="00:02:05.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.39" />
                    <SPLIT distance="100" swimtime="00:01:02.50" />
                    <SPLIT distance="150" swimtime="00:01:35.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="584" swimtime="00:00:56.59" resultid="3321" heatid="4764" lane="5" entrytime="00:00:53.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="503" swimtime="00:01:06.98" resultid="3322" heatid="4793" lane="3" entrytime="00:01:04.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sylwia" lastname="Gorockiewicz" birthdate="1975-03-29" gender="F" nation="POL" license="500115600525" athleteid="3333">
              <RESULTS>
                <RESULT eventid="1059" points="97" swimtime="00:00:57.20" resultid="3334" heatid="4665" lane="5" entrytime="00:01:00.90" entrycourse="SCM" />
                <RESULT eventid="1269" points="180" swimtime="00:04:40.06" resultid="3335" heatid="4726" lane="3" entrytime="00:04:58.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.34" />
                    <SPLIT distance="100" swimtime="00:02:12.89" />
                    <SPLIT distance="150" swimtime="00:03:26.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1575" points="131" swimtime="00:02:19.07" resultid="3336" heatid="4765" lane="3" entrytime="00:02:21.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Błażej" lastname="Wachowski" birthdate="1980-10-08" gender="M" nation="POL" license="100115700545" athleteid="3313">
              <RESULTS>
                <RESULT eventid="1199" points="490" swimtime="00:02:19.63" resultid="3314" heatid="4712" lane="3" entrytime="00:02:16.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.91" />
                    <SPLIT distance="100" swimtime="00:01:07.47" />
                    <SPLIT distance="150" swimtime="00:01:43.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1255" points="449" swimtime="00:01:10.27" resultid="3315" heatid="4722" lane="4" entrytime="00:01:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="414" swimtime="00:02:45.00" resultid="3316" heatid="4782" lane="6" entrytime="00:02:41.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                    <SPLIT distance="100" swimtime="00:01:18.01" />
                    <SPLIT distance="150" swimtime="00:02:01.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="503" swimtime="00:05:02.63" resultid="3317" heatid="4810" lane="5" entrytime="00:04:57.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.80" />
                    <SPLIT distance="100" swimtime="00:01:13.87" />
                    <SPLIT distance="150" swimtime="00:01:53.00" />
                    <SPLIT distance="200" swimtime="00:02:31.93" />
                    <SPLIT distance="250" swimtime="00:03:10.55" />
                    <SPLIT distance="300" swimtime="00:03:48.83" />
                    <SPLIT distance="350" swimtime="00:04:27.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Szymkowiak" birthdate="1980-04-12" gender="M" nation="POL" license="500115700523" athleteid="3308">
              <RESULTS>
                <RESULT eventid="1102" points="647" swimtime="00:00:26.31" resultid="3309" heatid="4680" lane="4" entrytime="00:00:25.63" entrycourse="SCM" />
                <RESULT eventid="1171" points="730" swimtime="00:00:31.17" resultid="3310" heatid="4703" lane="4" entrytime="00:00:31.33" entrycourse="SCM" />
                <RESULT eventid="1589" points="647" swimtime="00:01:11.01" resultid="3311" heatid="4774" lane="5" entrytime="00:01:10.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="3312" heatid="4793" lane="6" entrytime="00:01:08.72" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Kotecka" birthdate="1965-05-08" gender="F" nation="POL" license="100115600357" athleteid="3328">
              <RESULTS>
                <RESULT eventid="1129" points="300" swimtime="00:01:40.29" resultid="3329" heatid="4684" lane="2" entrytime="00:01:37.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1185" points="366" swimtime="00:03:06.78" resultid="3330" heatid="4707" lane="6" entrytime="00:03:00.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.88" />
                    <SPLIT distance="100" swimtime="00:01:29.99" />
                    <SPLIT distance="150" swimtime="00:02:18.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="353" swimtime="00:01:25.74" resultid="3331" heatid="4753" lane="2" entrytime="00:01:23.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1421" points="312" swimtime="00:03:34.14" resultid="3332" heatid="4776" lane="1" entrytime="00:03:28.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.67" />
                    <SPLIT distance="100" swimtime="00:01:44.15" />
                    <SPLIT distance="150" swimtime="00:02:40.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1325" points="679" swimtime="00:03:55.97" resultid="3342" heatid="4737" lane="4" entrytime="00:03:58.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.15" />
                    <SPLIT distance="100" swimtime="00:01:01.32" />
                    <SPLIT distance="150" swimtime="00:01:29.33" />
                    <SPLIT distance="200" swimtime="00:01:59.77" />
                    <SPLIT distance="250" swimtime="00:02:29.36" />
                    <SPLIT distance="300" swimtime="00:03:01.10" />
                    <SPLIT distance="350" swimtime="00:03:26.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3337" number="1" />
                    <RELAYPOSITION athleteid="3313" number="2" />
                    <RELAYPOSITION athleteid="3308" number="3" />
                    <RELAYPOSITION athleteid="3318" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1350" points="636" swimtime="00:01:59.68" resultid="3343" heatid="4740" lane="2" entrytime="00:01:58.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                    <SPLIT distance="100" swimtime="00:01:01.82" />
                    <SPLIT distance="150" swimtime="00:01:31.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3318" number="1" />
                    <RELAYPOSITION athleteid="3308" number="2" />
                    <RELAYPOSITION athleteid="3337" number="3" />
                    <RELAYPOSITION athleteid="3313" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="IKSKRA" nation="POL" region="06" clubid="2308" name="IKS DSS Kraków">
          <CONTACT city="Kraków" name="Bochenek" state="MAŁOP" street="Anna" />
          <ATHLETES>
            <ATHLETE firstname="Ewa" lastname="Rupp" birthdate="1956-03-06" gender="F" nation="POL" athleteid="2309">
              <RESULTS>
                <RESULT eventid="1129" points="168" swimtime="00:02:12.52" resultid="2310" heatid="4683" lane="5" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="173" swimtime="00:04:57.91" resultid="2311" heatid="4714" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.52" />
                    <SPLIT distance="100" swimtime="00:02:22.64" />
                    <SPLIT distance="150" swimtime="00:03:51.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="150" swimtime="00:02:01.24" resultid="2312" heatid="4752" lane="2" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1533" points="177" swimtime="00:08:57.57" resultid="2313" heatid="4804" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.53" />
                    <SPLIT distance="100" swimtime="00:02:06.66" />
                    <SPLIT distance="150" swimtime="00:03:15.98" />
                    <SPLIT distance="200" swimtime="00:04:25.88" />
                    <SPLIT distance="250" swimtime="00:05:35.06" />
                    <SPLIT distance="300" swimtime="00:06:43.27" />
                    <SPLIT distance="350" swimtime="00:07:50.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIEPOZ" nation="POL" region="15" clubid="3287" name="Zawodnik Niezrzeszony Poznań">
          <ATHLETES>
            <ATHLETE firstname="Krzysztof" lastname="Kubiak" birthdate="1989-07-05" gender="M" nation="POL" athleteid="3289">
              <RESULTS>
                <RESULT eventid="1143" points="129" swimtime="00:01:44.00" resultid="3290" heatid="4687" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1255" points="175" swimtime="00:01:33.84" resultid="3291" heatid="4721" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="281" swimtime="00:05:54.22" resultid="3293" heatid="4809" lane="2" entrytime="00:05:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.56" />
                    <SPLIT distance="100" swimtime="00:01:23.05" />
                    <SPLIT distance="150" swimtime="00:02:07.79" />
                    <SPLIT distance="200" swimtime="00:02:52.46" />
                    <SPLIT distance="250" swimtime="00:03:38.67" />
                    <SPLIT distance="300" swimtime="00:04:23.63" />
                    <SPLIT distance="350" swimtime="00:05:09.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="177" swimtime="00:03:22.26" resultid="4824" heatid="4782" lane="1" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.20" />
                    <SPLIT distance="100" swimtime="00:01:39.65" />
                    <SPLIT distance="150" swimtime="00:02:31.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Kędzior" birthdate="1973-12-08" gender="M" nation="POL" athleteid="3288">
              <RESULTS>
                <RESULT eventid="1102" points="342" swimtime="00:00:32.66" resultid="3294" heatid="4674" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1227" points="229" swimtime="00:03:23.60" resultid="3295" heatid="4716" lane="4" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.12" />
                    <SPLIT distance="100" swimtime="00:01:35.18" />
                    <SPLIT distance="150" swimtime="00:02:41.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="322" swimtime="00:01:12.90" resultid="3296" heatid="4760" lane="4" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="323" swimtime="00:05:54.29" resultid="3297" heatid="4809" lane="6" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.31" />
                    <SPLIT distance="100" swimtime="00:01:21.98" />
                    <SPLIT distance="150" swimtime="00:02:06.79" />
                    <SPLIT distance="200" swimtime="00:02:53.24" />
                    <SPLIT distance="250" swimtime="00:03:38.51" />
                    <SPLIT distance="300" swimtime="00:04:24.57" />
                    <SPLIT distance="350" swimtime="00:05:10.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIECZE" nation="POL" region="11" clubid="1607" name="Zawodnik Niezrzeszony Częstochowa" shortname="Zawodnik Niezrzeszony Częstoch">
          <ATHLETES>
            <ATHLETE firstname="Izabela" lastname="Wypych-Staszewska" birthdate="1970-08-16" gender="F" nation="POL" athleteid="2156">
              <RESULTS>
                <RESULT eventid="1059" points="363" swimtime="00:00:36.81" resultid="2157" heatid="4666" lane="3" entrytime="00:00:37.00" />
                <RESULT eventid="1358" points="347" swimtime="00:00:41.62" resultid="2158" heatid="4741" lane="4" entrytime="00:00:41.00" />
                <RESULT eventid="1393" points="399" swimtime="00:01:19.63" resultid="2159" heatid="4753" lane="4" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SWIRZE" nation="POL" region="08" clubid="3496" name="SWIM TRI Rzeszów">
          <CONTACT city="Rzeszów" name="SWIM TRI RZESZÓW" state="PODKA" />
          <ATHLETES>
            <ATHLETE firstname="Mariusz" lastname="Faff" birthdate="1963-11-15" gender="M" nation="POL" athleteid="3501">
              <RESULTS>
                <RESULT eventid="1102" points="602" swimtime="00:00:28.86" resultid="3502" heatid="4677" lane="3" entrytime="00:00:28.28" />
                <RESULT eventid="1199" points="516" swimtime="00:02:28.46" resultid="3503" heatid="4712" lane="6" entrytime="00:02:38.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                    <SPLIT distance="100" swimtime="00:01:09.67" />
                    <SPLIT distance="150" swimtime="00:01:49.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="556" swimtime="00:00:32.14" resultid="3504" heatid="4747" lane="2" entrytime="00:00:32.87" />
                <RESULT eventid="1407" points="572" swimtime="00:01:05.42" resultid="3505" heatid="4762" lane="6" entrytime="00:01:05.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Sarna" birthdate="1975-10-31" gender="M" nation="POL" athleteid="3497">
              <RESULTS>
                <RESULT eventid="1102" points="595" swimtime="00:00:27.16" resultid="3498" heatid="4679" lane="4" entrytime="00:00:26.44" />
                <RESULT eventid="1199" points="570" swimtime="00:02:16.13" resultid="3499" heatid="4713" lane="1" entrytime="00:02:11.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.06" />
                    <SPLIT distance="100" swimtime="00:01:02.16" />
                    <SPLIT distance="150" swimtime="00:01:38.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="581" swimtime="00:00:59.91" resultid="3500" heatid="4763" lane="1" entrytime="00:00:59.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="BAZMYS" nation="POL" region="11" clubid="3243" name="Baza pływania Mysłowice">
          <CONTACT city="41-200" email="adrian.kisiel93@gmail.com" name="Kisiel" phone="502593038" state="ŚLĄSK" street="Czarna" zip="8" />
          <ATHLETES>
            <ATHLETE firstname="Adrian" lastname="Kisiel" birthdate="1993-03-26" gender="M" nation="POL" athleteid="3244">
              <RESULTS>
                <RESULT eventid="1143" points="658" swimtime="00:01:00.86" resultid="3245" heatid="4690" lane="2" entrytime="00:00:59.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1255" status="DNS" swimtime="00:00:00.00" resultid="3246" heatid="4725" lane="1" entrytime="00:00:59.00" entrycourse="SCM" />
                <RESULT eventid="1379" points="680" swimtime="00:00:26.33" resultid="3247" heatid="4751" lane="1" entrytime="00:00:25.50" entrycourse="SCM" />
                <RESULT eventid="1435" points="589" swimtime="00:02:18.62" resultid="3248" heatid="4779" lane="4" entrytime="00:02:12.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                    <SPLIT distance="100" swimtime="00:01:05.72" />
                    <SPLIT distance="150" swimtime="00:01:42.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Kisiel" birthdate="1996-05-27" gender="F" nation="POL" athleteid="3259">
              <RESULTS>
                <RESULT eventid="1129" points="624" swimtime="00:01:10.96" resultid="3260" heatid="4685" lane="4" entrytime="00:01:11.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1505" points="606" swimtime="00:00:32.94" resultid="3261" heatid="4798" lane="5" entrytime="00:00:33.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewa" lastname="Dymarek" birthdate="1995-01-21" gender="F" nation="POL" athleteid="3254">
              <RESULTS>
                <RESULT eventid="1157" points="634" swimtime="00:00:35.50" resultid="3255" heatid="4694" lane="5" entrytime="00:00:36.73" entrycourse="SCM" />
                <RESULT eventid="1269" points="695" swimtime="00:02:47.49" resultid="3256" heatid="4729" lane="4" entrytime="00:02:50.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.20" />
                    <SPLIT distance="100" swimtime="00:01:20.12" />
                    <SPLIT distance="150" swimtime="00:02:03.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1575" points="656" swimtime="00:01:16.91" resultid="3257" heatid="4768" lane="4" entrytime="00:01:17.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1533" status="DNS" swimtime="00:00:00.00" resultid="3258" heatid="4806" lane="3" entrytime="00:04:55.55" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Czwartosz" birthdate="1993-04-08" gender="M" nation="POL" athleteid="3249">
              <RESULTS>
                <RESULT eventid="1102" points="560" swimtime="00:00:25.81" resultid="3250" heatid="4681" lane="5" entrytime="00:00:25.00" entrycourse="SCM" />
                <RESULT eventid="1227" points="502" swimtime="00:02:29.60" resultid="3251" heatid="4717" lane="3" entrytime="00:02:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:12.15" />
                    <SPLIT distance="150" swimtime="00:01:55.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="589" swimtime="00:00:27.62" resultid="3252" heatid="4750" lane="2" entrytime="00:00:27.00" entrycourse="SCM" />
                <RESULT eventid="1491" points="517" swimtime="00:01:05.78" resultid="3253" heatid="4794" lane="1" entrytime="00:01:04.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIEWOD" nation="POL" region="11" clubid="2184" name="Zawodnik Niezrzeszony Wodzisław Śląski" shortname="Zawodnik Niezrzeszony Wodzisła">
          <ATHLETES>
            <ATHLETE firstname="Michał" lastname="Brochocki" birthdate="2000-04-27" gender="M" nation="POL" athleteid="2185">
              <RESULTS>
                <RESULT eventid="1102" swimtime="00:00:26.46" resultid="2186" heatid="4679" lane="5" entrytime="00:00:27.00" />
                <RESULT eventid="1171" swimtime="00:00:34.87" resultid="2187" heatid="4701" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1379" swimtime="00:00:28.95" resultid="2188" heatid="4749" lane="2" entrytime="00:00:28.84" />
                <RESULT eventid="1491" swimtime="00:01:09.18" resultid="2189" heatid="4792" lane="2" entrytime="00:01:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06611" nation="POL" region="11" clubid="3605" name="MKP Wodnik 29 Tychy">
          <CONTACT city="Tychy" email="marekmrozw29@gmail.com" name="Mróz Marek" phone="782-985-239" state="ŚLĄSK" street="Damrota 170" zip="43-100" />
          <ATHLETES>
            <ATHLETE firstname="Anna" lastname="Zawadzka" birthdate="2000-06-22" gender="F" nation="POL" athleteid="3606">
              <RESULTS>
                <RESULT eventid="1059" swimtime="00:00:29.22" resultid="3607" heatid="4669" lane="6" entrytime="00:00:28.50" />
                <RESULT eventid="1393" swimtime="00:01:03.85" resultid="3608" heatid="4756" lane="1" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Poprawa - Jakubas" birthdate="2002-10-01" gender="M" nation="POL" athleteid="3609">
              <RESULTS>
                <RESULT eventid="1171" swimtime="00:00:30.01" resultid="3610" heatid="4704" lane="2" entrytime="00:00:30.00" />
                <RESULT eventid="1283" swimtime="00:02:23.57" resultid="3611" heatid="4734" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                    <SPLIT distance="100" swimtime="00:01:10.12" />
                    <SPLIT distance="150" swimtime="00:01:47.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1589" swimtime="00:01:05.28" resultid="3612" heatid="4775" lane="4" entrytime="00:01:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" swimtime="00:02:15.53" resultid="3613" heatid="4782" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.42" />
                    <SPLIT distance="100" swimtime="00:01:04.75" />
                    <SPLIT distance="150" swimtime="00:01:40.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIEUKR" nation="UKR" clubid="3823" name="Zawodnik Niezrzeszony Kijów">
          <ATHLETES>
            <ATHLETE firstname="Tetiana" lastname="Sytnyak" birthdate="1985-06-15" gender="F" nation="UKR" athleteid="3824">
              <RESULTS>
                <RESULT eventid="1129" points="146" swimtime="00:01:54.75" resultid="3825" heatid="4684" lane="6" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1185" points="191" swimtime="00:03:33.86" resultid="3826" heatid="4706" lane="6" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.63" />
                    <SPLIT distance="100" swimtime="00:01:42.03" />
                    <SPLIT distance="150" swimtime="00:02:38.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1505" points="157" swimtime="00:00:51.22" resultid="3827" heatid="4796" lane="5" entrytime="00:00:50.10" />
                <RESULT eventid="1393" points="193" swimtime="00:01:35.07" resultid="3828" heatid="4752" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIEMYS" nation="POL" region="11" clubid="3304" name="Zawodnik Niezrzeszony Mysłowice">
          <CONTACT name="Zawodnik Niezrzeszony Mysłowice" />
        </CLUB>
        <CLUB type="CLUB" code="UNIWAR" nation="POL" region="14" clubid="3595" name="KU AZS Uniwersytetu Warszawskiego" shortname="KU AZS Uniwersytetu Warszawski">
          <CONTACT city="Warszawa" name="Rębas" state="MAZOW" />
          <ATHLETES>
            <ATHLETE firstname="Igor" lastname="Rębas" birthdate="1989-01-01" gender="M" nation="POL" athleteid="3596">
              <RESULTS>
                <RESULT eventid="1255" status="DNS" swimtime="00:00:00.00" resultid="3597" heatid="4725" lane="5" entrytime="00:00:58.66" />
                <RESULT eventid="1407" status="DNS" swimtime="00:00:00.00" resultid="3598" heatid="4764" lane="4" entrytime="00:00:53.17" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MASOPO" nation="POL" region="07" clubid="3266" name="T.P. MASTERS Opole">
          <CONTACT city="Opole" name="KRASNODĘBSKI" state="OPOLS" />
          <ATHLETES>
            <ATHLETE firstname="Agnieszka" lastname="Bartnikowska" birthdate="1990-01-01" gender="F" nation="POL" athleteid="3267">
              <RESULTS>
                <RESULT eventid="1129" points="589" swimtime="00:01:12.65" resultid="3268" heatid="4685" lane="2" entrytime="00:01:11.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="523" swimtime="00:00:33.62" resultid="3269" heatid="4742" lane="5" entrytime="00:00:34.25" />
                <RESULT eventid="1505" points="536" swimtime="00:00:33.77" resultid="3270" heatid="4798" lane="1" entrytime="00:00:33.09" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zbigniew" lastname="Januszkiewicz" birthdate="1962-01-01" gender="M" nation="POL" athleteid="3271">
              <RESULTS>
                <RESULT eventid="1143" points="846" swimtime="00:01:06.77" resultid="3272" heatid="4690" lane="1" entrytime="00:01:06.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1255" points="665" swimtime="00:01:08.97" resultid="3273" heatid="4722" lane="1" entrytime="00:01:12.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1435" points="820" swimtime="00:02:26.55" resultid="3274" heatid="4779" lane="2" entrytime="00:02:24.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                    <SPLIT distance="100" swimtime="00:01:12.93" />
                    <SPLIT distance="150" swimtime="00:01:50.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1519" points="870" swimtime="00:00:30.84" resultid="3275" heatid="4803" lane="1" entrytime="00:00:30.87" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="REKMIK" nation="POL" region="11" clubid="3664" name="KS REKIN Kamionka Mikołów">
          <ATHLETES>
            <ATHLETE firstname="Przemysław" lastname="Wańha" birthdate="1983-04-19" gender="M" nation="POL" athleteid="3665">
              <RESULTS>
                <RESULT eventid="1102" points="391" swimtime="00:00:29.44" resultid="3666" heatid="4676" lane="2" entrytime="00:00:29.72" />
                <RESULT eventid="1199" points="382" swimtime="00:02:29.38" resultid="3667" heatid="4711" lane="3" entrytime="00:02:39.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                    <SPLIT distance="100" swimtime="00:01:12.63" />
                    <SPLIT distance="150" swimtime="00:01:51.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" status="DNS" swimtime="00:00:00.00" resultid="3668" heatid="4746" lane="3" entrytime="00:00:33.15" />
                <RESULT eventid="1407" points="388" swimtime="00:01:05.40" resultid="3669" heatid="4761" lane="1" entrytime="00:01:09.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ACAOLA" nation="POL" region="01" clubid="3599" name="MKS Swim Academy Termy Jakuba Oława" shortname="MKS Swim Academy Termy Jakuba ">
          <CONTACT city="Oława" email="biuro@swim-academy.pl" internet="www.swim-academy.pl" name="Grzegorz Fidala / Jacek Bereżnicki" phone="601316031 / 69643365" state="DOLNO" street="1 Maja 33a" zip="55-200" />
          <ATHLETES>
            <ATHLETE firstname="Magdalena" lastname="Chorąży" birthdate="1978-09-27" gender="F" nation="POL" license="104501600044" athleteid="3600">
              <RESULTS>
                <RESULT eventid="1157" points="623" swimtime="00:00:37.66" resultid="3601" heatid="4693" lane="4" entrytime="00:00:38.90" />
                <RESULT eventid="1269" points="539" swimtime="00:03:07.19" resultid="3602" heatid="4728" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.78" />
                    <SPLIT distance="100" swimtime="00:01:30.85" />
                    <SPLIT distance="150" swimtime="00:02:20.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="634" swimtime="00:00:32.81" resultid="3603" heatid="4742" lane="4" entrytime="00:00:33.90" />
                <RESULT eventid="1575" status="DNS" swimtime="00:00:00.00" resultid="3604" heatid="4767" lane="4" entrytime="00:01:26.80" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03311" nation="POL" region="11" clubid="3154" name="UKS WODNIK 29 Katowice">
          <CONTACT city="Katowice" email="biuro.wodnik29@gmail.com" name="Spławiński" phone="603646226" state="ŚLĄSK" />
          <ATHLETES>
            <ATHLETE firstname="Julia" lastname="Koral" birthdate="1998-01-01" gender="F" nation="POL" athleteid="3214">
              <RESULTS>
                <RESULT eventid="1129" swimtime="00:01:21.66" resultid="3215" heatid="4685" lane="6" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1477" swimtime="00:01:23.56" resultid="3216" heatid="4785" lane="4" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1505" swimtime="00:00:38.47" resultid="3217" heatid="4798" lane="2" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Oracz" birthdate="1971-01-01" gender="F" nation="POL" athleteid="3189">
              <RESULTS>
                <RESULT eventid="1185" status="DNS" swimtime="00:00:00.00" resultid="3190" heatid="4706" lane="2" entrytime="00:03:15.00" />
                <RESULT eventid="1269" status="DNS" swimtime="00:00:00.00" resultid="3191" heatid="4728" lane="6" entrytime="00:03:40.00" />
                <RESULT eventid="1533" status="DNS" swimtime="00:00:00.00" resultid="3192" heatid="4805" lane="1" entrytime="00:06:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dominik" lastname="Sieroń" birthdate="1981-08-22" gender="M" nation="POL" athleteid="4006">
              <RESULTS>
                <RESULT eventid="1171" points="359" swimtime="00:00:39.47" resultid="4007" heatid="4697" lane="5" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Sikora" birthdate="1996-11-14" gender="F" nation="POL" athleteid="3179">
              <RESULTS>
                <RESULT eventid="1505" points="610" swimtime="00:00:32.87" resultid="3180" heatid="4798" lane="6" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Mroziński" birthdate="1959-01-01" gender="M" nation="POL" athleteid="3166">
              <RESULTS>
                <RESULT eventid="1171" points="670" swimtime="00:00:36.01" resultid="3167" heatid="4701" lane="6" entrytime="00:00:35.50" />
                <RESULT eventid="1283" points="544" swimtime="00:03:06.56" resultid="3168" heatid="4732" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.15" />
                    <SPLIT distance="100" swimtime="00:01:29.91" />
                    <SPLIT distance="150" swimtime="00:02:17.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1589" points="588" swimtime="00:01:23.01" resultid="3169" heatid="4772" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agata" lastname="Kowalczyk" birthdate="2001-01-01" gender="F" nation="POL" athleteid="3174">
              <RESULTS>
                <RESULT eventid="1157" swimtime="00:00:37.45" resultid="3175" heatid="4694" lane="4" entrytime="00:00:35.50" />
                <RESULT eventid="1269" swimtime="00:02:59.83" resultid="3176" heatid="4729" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.16" />
                    <SPLIT distance="100" swimtime="00:01:26.00" />
                    <SPLIT distance="150" swimtime="00:02:12.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1575" swimtime="00:01:23.89" resultid="3177" heatid="4767" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1477" swimtime="00:01:16.22" resultid="3178" heatid="4785" lane="2" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Ferdek" birthdate="1988-07-12" gender="F" nation="POL" athleteid="3197">
              <RESULTS>
                <RESULT eventid="1393" points="453" swimtime="00:01:11.31" resultid="3198" heatid="4755" lane="1" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1505" status="DNS" swimtime="00:00:00.00" resultid="3199" heatid="4797" lane="1" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jarosław" lastname="Silwonik" birthdate="1966-11-14" gender="M" nation="POL" athleteid="3204">
              <RESULTS>
                <RESULT eventid="1102" points="640" swimtime="00:00:28.28" resultid="3205" heatid="4677" lane="5" entrytime="00:00:29.00" />
                <RESULT eventid="1379" points="556" swimtime="00:00:32.14" resultid="3206" heatid="4748" lane="6" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Weronika" lastname="Grychtoł" birthdate="2001-02-10" gender="F" nation="POL" athleteid="3207">
              <RESULTS>
                <RESULT eventid="1421" swimtime="00:02:47.44" resultid="3208" heatid="4776" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                    <SPLIT distance="100" swimtime="00:01:22.04" />
                    <SPLIT distance="150" swimtime="00:02:04.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1533" swimtime="00:05:21.44" resultid="3209" heatid="4806" lane="6" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                    <SPLIT distance="100" swimtime="00:01:17.00" />
                    <SPLIT distance="150" swimtime="00:01:57.32" />
                    <SPLIT distance="200" swimtime="00:02:37.80" />
                    <SPLIT distance="250" swimtime="00:03:18.74" />
                    <SPLIT distance="300" swimtime="00:03:59.91" />
                    <SPLIT distance="350" swimtime="00:04:41.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Cichecka" birthdate="1983-02-05" gender="F" nation="POL" athleteid="3210">
              <RESULTS>
                <RESULT eventid="1157" points="112" swimtime="00:01:05.77" resultid="3211" heatid="4692" lane="5" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jolanta" lastname="Stefanek" birthdate="1960-03-15" gender="F" nation="POL" athleteid="3200">
              <RESULTS>
                <RESULT eventid="1157" points="466" swimtime="00:00:47.83" resultid="3201" heatid="4692" lane="1" entrytime="00:00:50.00" />
                <RESULT eventid="1269" points="455" swimtime="00:03:50.14" resultid="3202" heatid="4727" lane="2" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.43" />
                    <SPLIT distance="100" swimtime="00:01:50.71" />
                    <SPLIT distance="150" swimtime="00:02:51.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1575" points="413" swimtime="00:01:48.14" resultid="3203" heatid="4766" lane="2" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Magdalena" lastname="Madejska" birthdate="1982-01-01" gender="F" nation="POL" athleteid="3181">
              <RESULTS>
                <RESULT eventid="1358" points="252" swimtime="00:00:44.64" resultid="3182" heatid="4741" lane="5" entrytime="00:00:45.00" />
                <RESULT eventid="1393" points="215" swimtime="00:01:35.32" resultid="3183" heatid="4753" lane="5" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Ilnicki" birthdate="1956-01-01" gender="M" nation="POL" athleteid="4815">
              <RESULTS>
                <RESULT eventid="1171" status="DNS" swimtime="00:00:00.00" resultid="4816" heatid="4695" lane="5" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Koenig" birthdate="1987-01-01" gender="F" nation="POL" athleteid="3184">
              <RESULTS>
                <RESULT eventid="1157" points="163" swimtime="00:00:57.95" resultid="3185" heatid="4691" lane="3" entrytime="00:01:00.00" />
                <RESULT eventid="1269" points="160" swimtime="00:04:37.35" resultid="3186" heatid="4727" lane="1" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.81" />
                    <SPLIT distance="100" swimtime="00:02:07.12" />
                    <SPLIT distance="150" swimtime="00:03:21.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1575" points="174" swimtime="00:02:03.75" resultid="3187" heatid="4766" lane="6" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1505" points="79" swimtime="00:01:04.37" resultid="3188" heatid="4795" lane="3" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Kołodziej" birthdate="2002-01-01" gender="M" nation="POL" athleteid="3162">
              <RESULTS>
                <RESULT eventid="1102" swimtime="00:00:26.15" resultid="3163" heatid="4679" lane="1" entrytime="00:00:27.00" />
                <RESULT eventid="1171" swimtime="00:00:33.62" resultid="3164" heatid="4703" lane="6" entrytime="00:00:32.00" />
                <RESULT eventid="1407" swimtime="00:00:57.33" resultid="3165" heatid="4763" lane="2" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Dąbrowski" birthdate="1988-02-20" gender="M" nation="POL" athleteid="3155">
              <RESULTS>
                <RESULT eventid="1102" points="666" swimtime="00:00:24.66" resultid="3156" heatid="4681" lane="4" entrytime="00:00:24.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Radosław" lastname="Łapot" birthdate="1999-05-25" gender="M" nation="POL" athleteid="3849">
              <RESULTS>
                <RESULT eventid="1283" swimtime="00:02:38.92" resultid="3850" heatid="4734" lane="4" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                    <SPLIT distance="100" swimtime="00:01:14.08" />
                    <SPLIT distance="150" swimtime="00:01:54.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Bajura" birthdate="1998-10-22" gender="F" nation="POL" athleteid="3212">
              <RESULTS>
                <RESULT eventid="1505" swimtime="00:00:33.20" resultid="3213" heatid="4797" lane="3" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Wiśniewski" birthdate="1987-11-13" gender="M" nation="POL" athleteid="3829">
              <RESULTS>
                <RESULT eventid="1379" points="657" swimtime="00:00:26.59" resultid="3830" heatid="4751" lane="4" entrytime="00:00:25.10" />
                <RESULT eventid="1519" points="703" swimtime="00:00:27.53" resultid="3831" heatid="4803" lane="2" entrytime="00:00:27.40" />
                <RESULT eventid="1255" points="686" swimtime="00:00:59.84" resultid="3832" heatid="4725" lane="4" entrytime="00:00:56.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Niedziela- Sołtysiak" birthdate="1972-01-27" gender="F" nation="POL" athleteid="3851">
              <RESULTS>
                <RESULT eventid="1129" points="413" swimtime="00:01:28.45" resultid="3852" heatid="4684" lane="1" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1505" status="DNS" swimtime="00:00:00.00" resultid="3853" heatid="4796" lane="2" entrytime="00:00:50.00" />
                <RESULT eventid="1575" points="408" swimtime="00:01:41.13" resultid="3854" heatid="4766" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krystyna" lastname="Nicpoń" birthdate="1940-01-01" gender="F" nation="POL" athleteid="3193">
              <RESULTS>
                <RESULT eventid="1059" points="117" swimtime="00:01:13.72" resultid="3194" heatid="4665" lane="1" entrytime="00:01:20.00" />
                <RESULT eventid="1393" points="122" swimtime="00:02:43.77" resultid="3195" heatid="4752" lane="1" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1505" points="184" swimtime="00:01:18.75" resultid="3196" heatid="4795" lane="4" entrytime="00:01:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kamil" lastname="Ogorzałek" birthdate="1999-01-01" gender="M" nation="POL" athleteid="3157">
              <RESULTS>
                <RESULT eventid="1102" swimtime="00:00:24.52" resultid="3158" heatid="4682" lane="1" entrytime="00:00:24.30" />
                <RESULT eventid="1199" swimtime="00:01:57.33" resultid="3159" heatid="4713" lane="3" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.22" />
                    <SPLIT distance="100" swimtime="00:00:58.65" />
                    <SPLIT distance="150" swimtime="00:01:29.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" swimtime="00:00:26.38" resultid="3160" heatid="4750" lane="4" entrytime="00:00:26.30" />
                <RESULT eventid="1407" swimtime="00:00:52.80" resultid="3161" heatid="4764" lane="2" entrytime="00:00:53.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Urszula" lastname="Walkowicz" birthdate="1932-05-18" gender="F" nation="POL" athleteid="3836">
              <RESULTS>
                <RESULT eventid="1059" points="121" swimtime="00:01:31.89" resultid="3837" heatid="4665" lane="6" entrytime="00:01:30.00" />
                <RESULT eventid="1505" points="335" swimtime="00:01:20.03" resultid="3838" heatid="4795" lane="2" entrytime="00:01:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edyta" lastname="Mróz" birthdate="1979-06-09" gender="F" nation="POL" athleteid="3835">
              <RESULTS>
                <RESULT eventid="1129" status="DNS" swimtime="00:00:00.00" resultid="3839" heatid="4684" lane="5" entrytime="00:01:40.00" />
                <RESULT eventid="1185" status="DNS" swimtime="00:00:00.00" resultid="3840" heatid="4706" lane="4" entrytime="00:03:15.00" />
                <RESULT eventid="1421" status="DNS" swimtime="00:00:00.00" resultid="3841" heatid="4776" lane="5" entrytime="00:03:15.00" />
                <RESULT eventid="1505" status="DNS" swimtime="00:00:00.00" resultid="3842" heatid="4797" lane="4" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Wilczek" birthdate="1958-03-01" gender="M" nation="POL" athleteid="3170">
              <RESULTS>
                <RESULT eventid="1102" points="544" swimtime="00:00:30.51" resultid="3171" heatid="4676" lane="4" entrytime="00:00:29.50" />
                <RESULT eventid="1255" points="362" swimtime="00:01:24.43" resultid="3172" heatid="4721" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="471" swimtime="00:00:34.43" resultid="3173" heatid="4746" lane="2" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1350" status="DNS" swimtime="00:00:00.00" resultid="3223" heatid="4739" lane="5">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3166" number="1" />
                    <RELAYPOSITION athleteid="3170" number="2" />
                    <RELAYPOSITION athleteid="3155" number="3" />
                    <RELAYPOSITION athleteid="3829" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1329" points="140" swimtime="00:04:28.78" resultid="3224" heatid="4738" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.09" />
                    <SPLIT distance="100" swimtime="00:02:13.33" />
                    <SPLIT distance="150" swimtime="00:03:07.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3193" number="1" />
                    <RELAYPOSITION athleteid="3184" number="2" />
                    <RELAYPOSITION athleteid="3200" number="3" />
                    <RELAYPOSITION athleteid="3836" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="ASBYD" nation="POL" region="02" clubid="2178" name="MKS ASTORIA Bydgoszcz" shortname="MKS ASTORIA Bydgoszcz	">
          <ATHLETES>
            <ATHLETE firstname="Dariusz" lastname="Kostkowski" birthdate="1970-01-13" gender="M" nation="POL" athleteid="2179">
              <RESULTS>
                <RESULT eventid="1143" points="119" swimtime="00:01:57.89" resultid="2180" heatid="4687" lane="6" entrytime="00:01:55.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="256" swimtime="00:00:46.80" resultid="2181" heatid="4697" lane="6" entrytime="00:00:45.57" />
                <RESULT eventid="1435" points="127" swimtime="00:04:12.69" resultid="2182" heatid="4777" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.48" />
                    <SPLIT distance="100" swimtime="00:02:01.90" />
                    <SPLIT distance="150" swimtime="00:03:07.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1519" points="144" swimtime="00:00:50.97" resultid="2183" heatid="4799" lane="3" entrytime="00:00:49.92" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MASWAR" nation="POL" region="14" clubid="2354" name="Warsaw Masters Team">
          <CONTACT city="Warszawa" email="marlena@masters.waw.pl" name="Dobrasiewicz" state="MAZOW" />
          <ATHLETES>
            <ATHLETE firstname="Rafał" lastname="Skośkiewicz" birthdate="1966-05-05" gender="M" nation="POL" athleteid="3455">
              <RESULTS>
                <RESULT eventid="1143" status="DNS" swimtime="00:00:00.00" resultid="3456" heatid="4689" lane="2" entrytime="00:01:09.00" />
                <RESULT eventid="1255" status="DNS" swimtime="00:00:00.00" resultid="3457" heatid="4723" lane="1" entrytime="00:01:08.00" />
                <RESULT eventid="1379" points="657" swimtime="00:00:30.40" resultid="3458" heatid="4747" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1491" points="677" swimtime="00:01:09.79" resultid="3459" heatid="4792" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mirosław" lastname="Warchoł" birthdate="1953-08-30" gender="M" nation="POL" athleteid="3483">
              <RESULTS>
                <RESULT eventid="1143" points="600" swimtime="00:01:20.26" resultid="3484" heatid="4688" lane="5" entrytime="00:01:18.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="423" swimtime="00:03:07.04" resultid="3485" heatid="4717" lane="1" entrytime="00:02:47.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.90" />
                    <SPLIT distance="100" swimtime="00:01:27.08" />
                    <SPLIT distance="150" swimtime="00:02:26.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1435" points="653" swimtime="00:02:53.99" resultid="3486" heatid="4778" lane="2" entrytime="00:02:48.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.29" />
                    <SPLIT distance="100" swimtime="00:01:25.33" />
                    <SPLIT distance="150" swimtime="00:02:09.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leszek" lastname="Madej" birthdate="1960-06-17" gender="M" nation="POL" athleteid="3465">
              <RESULTS>
                <RESULT eventid="1102" points="674" swimtime="00:00:28.40" resultid="3466" heatid="4678" lane="2" entrytime="00:00:27.70" />
                <RESULT eventid="1199" points="707" swimtime="00:02:16.57" resultid="3467" heatid="4712" lane="4" entrytime="00:02:18.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                    <SPLIT distance="100" swimtime="00:01:06.88" />
                    <SPLIT distance="150" swimtime="00:01:41.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="736" swimtime="00:01:01.87" resultid="3468" heatid="4762" lane="5" entrytime="00:01:02.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="3469" heatid="4792" lane="1" entrytime="00:01:11.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dymitr" lastname="Bielski" birthdate="1977-08-13" gender="M" nation="POL" athleteid="3460">
              <RESULTS>
                <RESULT eventid="1171" status="DNS" swimtime="00:00:00.00" resultid="3461" heatid="4700" lane="2" entrytime="00:00:37.00" />
                <RESULT eventid="1199" status="DNS" swimtime="00:00:00.00" resultid="3462" heatid="4711" lane="4" entrytime="00:02:40.00" />
                <RESULT eventid="1589" status="DNS" swimtime="00:00:00.00" resultid="3463" heatid="4773" lane="6" entrytime="00:01:20.00" />
                <RESULT eventid="1547" status="DNS" swimtime="00:00:00.00" resultid="3464" heatid="4809" lane="5" entrytime="00:05:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Witkowski" birthdate="1981-06-16" gender="M" nation="POL" athleteid="3470">
              <RESULTS>
                <RESULT eventid="1171" points="553" swimtime="00:00:34.18" resultid="3471" heatid="4701" lane="2" entrytime="00:00:34.50" />
                <RESULT eventid="1589" points="493" swimtime="00:01:17.77" resultid="3472" heatid="4773" lane="3" entrytime="00:01:16.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Ostrowski" birthdate="1977-05-14" gender="M" nation="POL" athleteid="3487">
              <RESULTS>
                <RESULT eventid="1171" points="698" swimtime="00:00:32.30" resultid="3488" heatid="4703" lane="2" entrytime="00:00:31.50" />
                <RESULT eventid="1589" points="656" swimtime="00:01:11.60" resultid="3489" heatid="4774" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" status="DNS" swimtime="00:00:00.00" resultid="3490" heatid="4809" lane="3" entrytime="00:05:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tomasz" lastname="Porada" birthdate="1983-06-10" gender="M" nation="POL" athleteid="3473">
              <RESULTS>
                <RESULT eventid="1171" points="503" swimtime="00:00:33.53" resultid="3474" heatid="4702" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="1283" points="596" swimtime="00:02:40.95" resultid="3475" heatid="4734" lane="6" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                    <SPLIT distance="100" swimtime="00:01:16.94" />
                    <SPLIT distance="150" swimtime="00:01:58.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" status="DNS" swimtime="00:00:00.00" resultid="3476" heatid="4762" lane="3" entrytime="00:00:59.97" />
                <RESULT eventid="1463" points="471" swimtime="00:02:38.11" resultid="3477" heatid="4782" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                    <SPLIT distance="100" swimtime="00:01:12.30" />
                    <SPLIT distance="150" swimtime="00:01:54.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Rogosz" birthdate="1976-04-28" gender="M" nation="POL" athleteid="3478">
              <RESULTS>
                <RESULT eventid="1143" points="395" swimtime="00:01:17.66" resultid="3479" heatid="4688" lane="1" entrytime="00:01:21.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1283" points="504" swimtime="00:02:50.22" resultid="3480" heatid="4733" lane="1" entrytime="00:02:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.21" />
                    <SPLIT distance="100" swimtime="00:01:22.96" />
                    <SPLIT distance="150" swimtime="00:02:06.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1589" points="505" swimtime="00:01:18.13" resultid="3481" heatid="4773" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" status="DNS" swimtime="00:00:00.00" resultid="3482" heatid="4781" lane="3" entrytime="00:02:50.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1350" status="DNS" swimtime="00:00:00.00" resultid="3491" heatid="4740" lane="5" entrytime="00:02:00.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3455" number="1" />
                    <RELAYPOSITION athleteid="3470" number="2" />
                    <RELAYPOSITION athleteid="3487" number="3" />
                    <RELAYPOSITION athleteid="3465" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="02211" nation="POL" region="11" clubid="2360" name="MUKS GILUS Gilowice">
          <CONTACT city="Miedźna" email="js.formasy@interia.pl" name="Gilus Gilowice" phone="793691105" state="ŚLĄSK" street="Korfantego 38" zip="43-227" />
          <ATHLETES>
            <ATHLETE firstname="Sławomir" lastname="Formas" birthdate="1969-11-05" gender="M" nation="POL" license="502211700187" athleteid="2361">
              <RESULTS>
                <RESULT eventid="1171" points="808" swimtime="00:00:31.90" resultid="2362" heatid="4703" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="1283" points="718" swimtime="00:02:35.66" resultid="2363" heatid="4733" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                    <SPLIT distance="100" swimtime="00:01:14.58" />
                    <SPLIT distance="150" swimtime="00:01:55.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1589" points="751" swimtime="00:01:10.72" resultid="2364" heatid="4774" lane="1" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="634" swimtime="00:01:07.17" resultid="2365" heatid="4793" lane="5" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Siedmina" birthdate="1980-06-26" gender="M" nation="POL" license="502211700190" athleteid="2371">
              <RESULTS>
                <RESULT eventid="1102" points="256" swimtime="00:00:35.83" resultid="2372" heatid="4674" lane="6" entrytime="00:00:33.50" />
                <RESULT eventid="1199" points="174" swimtime="00:03:17.35" resultid="2373" heatid="4709" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.37" />
                    <SPLIT distance="100" swimtime="00:01:30.51" />
                    <SPLIT distance="150" swimtime="00:02:21.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="231" swimtime="00:01:20.91" resultid="2374" heatid="4757" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Michalski" birthdate="2001-03-15" gender="M" nation="POL" license="102211700163" athleteid="2375">
              <RESULTS>
                <RESULT eventid="1102" swimtime="00:00:25.31" resultid="2376" heatid="4681" lane="6" entrytime="00:00:25.40" />
                <RESULT eventid="1199" swimtime="00:01:57.98" resultid="2377" heatid="4713" lane="4" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.79" />
                    <SPLIT distance="100" swimtime="00:00:58.55" />
                    <SPLIT distance="150" swimtime="00:01:28.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" swimtime="00:00:54.38" resultid="2378" heatid="4763" lane="4" entrytime="00:00:55.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" swimtime="00:04:18.43" resultid="2379" heatid="4810" lane="4" entrytime="00:04:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.92" />
                    <SPLIT distance="100" swimtime="00:01:01.55" />
                    <SPLIT distance="150" swimtime="00:01:34.20" />
                    <SPLIT distance="200" swimtime="00:02:07.59" />
                    <SPLIT distance="250" swimtime="00:02:40.73" />
                    <SPLIT distance="300" swimtime="00:03:13.92" />
                    <SPLIT distance="350" swimtime="00:03:47.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karol" lastname="Trela" birthdate="1998-03-16" gender="M" nation="POL" license="102211700189" athleteid="2366">
              <RESULTS>
                <RESULT eventid="1102" swimtime="00:00:25.94" resultid="2367" heatid="4680" lane="2" entrytime="00:00:25.80" />
                <RESULT eventid="1171" swimtime="00:00:30.22" resultid="2368" heatid="4703" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="1589" swimtime="00:01:07.75" resultid="2369" heatid="4775" lane="2" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" swimtime="00:01:03.86" resultid="2370" heatid="4793" lane="4" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MASLOD" nation="POL" region="05" clubid="2469" name="MASTERS Łódź">
          <CONTACT city="Łodź" email="sport@masterslodz.pl" internet="http://masterslodz.pl" name="Trudnos" phone="604184311" state="ŁÓDZK" />
          <ATHLETES>
            <ATHLETE firstname="Michał" lastname="Woźniak" birthdate="1981-08-25" gender="M" nation="POL" license="503605700034" athleteid="2470">
              <RESULTS>
                <RESULT eventid="1143" points="561" swimtime="00:01:06.50" resultid="2471" heatid="4690" lane="5" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1255" points="523" swimtime="00:01:06.80" resultid="2472" heatid="4723" lane="3" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1435" points="601" swimtime="00:02:26.75" resultid="2473" heatid="4779" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                    <SPLIT distance="100" swimtime="00:01:11.18" />
                    <SPLIT distance="150" swimtime="00:01:49.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1519" points="593" swimtime="00:00:30.33" resultid="2474" heatid="4803" lane="5" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAXSZA" nation="POL" region="15" clubid="2876" name="Max Masters Swimm Club Szamotuły" shortname="Max Masters Swimm Club Szamotu">
          <CONTACT city="Szamotuły" email="karolbartkowiak88@gmail.com" name="Bartkowiak" phone="721573722" />
          <ATHLETES>
            <ATHLETE firstname="Karol" lastname="Bartkowiak" birthdate="1988-01-25" gender="M" nation="POL" athleteid="2877">
              <RESULTS>
                <RESULT eventid="1102" points="457" swimtime="00:00:27.96" resultid="2878" heatid="4679" lane="6" entrytime="00:00:27.14" />
                <RESULT eventid="1255" points="399" swimtime="00:01:11.23" resultid="2879" heatid="4722" lane="3" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="426" swimtime="00:00:30.40" resultid="2880" heatid="4749" lane="1" entrytime="00:00:29.17" />
                <RESULT eventid="1407" status="DNS" swimtime="00:00:00.00" resultid="2881" heatid="4763" lane="6" entrytime="00:00:59.82" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Przemysław" lastname="Pernak" birthdate="1990-11-06" gender="M" nation="POL" athleteid="2882">
              <RESULTS>
                <RESULT eventid="1102" points="222" swimtime="00:00:35.55" resultid="2883" heatid="4671" lane="1" entrytime="00:00:39.00" />
                <RESULT eventid="1171" points="207" swimtime="00:00:45.20" resultid="2884" heatid="4697" lane="4" entrytime="00:00:43.50" />
                <RESULT eventid="1379" points="189" swimtime="00:00:39.82" resultid="2885" heatid="4744" lane="5" entrytime="00:00:42.00" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="2886" heatid="4787" lane="3" entrytime="00:03:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Sędrowicz" birthdate="1997-04-17" gender="M" nation="POL" athleteid="2892">
              <RESULTS>
                <RESULT eventid="1171" points="443" swimtime="00:00:35.41" resultid="2893" heatid="4702" lane="1" entrytime="00:00:34.00" />
                <RESULT eventid="1283" points="361" swimtime="00:02:59.11" resultid="2894" heatid="4733" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.82" />
                    <SPLIT distance="100" swimtime="00:01:24.58" />
                    <SPLIT distance="150" swimtime="00:02:12.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1589" points="405" swimtime="00:01:18.58" resultid="2895" heatid="4773" lane="4" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="347" swimtime="00:01:15.10" resultid="2896" heatid="4791" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Konrad" lastname="Zajas" birthdate="1999-06-16" gender="M" nation="POL" athleteid="2897">
              <RESULTS>
                <RESULT eventid="1102" swimtime="00:00:26.53" resultid="2898" heatid="4680" lane="6" entrytime="00:00:26.35" />
                <RESULT eventid="1255" swimtime="00:01:10.44" resultid="2899" heatid="4723" lane="6" entrytime="00:01:08.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" swimtime="00:00:30.53" resultid="2900" heatid="4749" lane="6" entrytime="00:00:29.19" />
                <RESULT eventid="1407" swimtime="00:01:00.26" resultid="2901" heatid="4762" lane="4" entrytime="00:01:00.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Szmania" birthdate="1984-12-17" gender="M" nation="POL" athleteid="2887">
              <RESULTS>
                <RESULT eventid="1102" points="241" swimtime="00:00:34.59" resultid="2888" heatid="4673" lane="5" entrytime="00:00:34.00" />
                <RESULT eventid="1171" points="262" swimtime="00:00:41.68" resultid="2889" heatid="4700" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1379" points="216" swimtime="00:00:38.55" resultid="2890" heatid="4745" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1491" points="202" swimtime="00:01:33.61" resultid="2891" heatid="4788" lane="4" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1325" points="333" swimtime="00:04:53.56" resultid="2902" heatid="4736" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.95" />
                    <SPLIT distance="100" swimtime="00:01:02.00" />
                    <SPLIT distance="150" swimtime="00:01:39.88" />
                    <SPLIT distance="200" swimtime="00:02:22.05" />
                    <SPLIT distance="250" swimtime="00:03:01.71" />
                    <SPLIT distance="300" swimtime="00:03:42.80" />
                    <SPLIT distance="350" swimtime="00:04:15.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2877" number="1" />
                    <RELAYPOSITION athleteid="2887" number="2" />
                    <RELAYPOSITION athleteid="2882" number="3" />
                    <RELAYPOSITION athleteid="2892" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1350" points="279" swimtime="00:02:30.63" resultid="2903" heatid="4739" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.39" />
                    <SPLIT distance="100" swimtime="00:01:26.14" />
                    <SPLIT distance="150" swimtime="00:01:56.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2882" number="1" />
                    <RELAYPOSITION athleteid="2892" number="2" />
                    <RELAYPOSITION athleteid="2877" number="3" />
                    <RELAYPOSITION athleteid="2887" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="NIESWI" nation="POL" region="01" clubid="2916" name="Zawodnik Niezrzeszony Świebodzice" shortname="Zawodnik Niezrzeszony Świebodz">
          <ATHLETES>
            <ATHLETE firstname="Agnieszka" lastname="Gajdowska" birthdate="1995-07-17" gender="F" nation="POL" athleteid="2918">
              <RESULTS>
                <RESULT eventid="1059" points="753" swimtime="00:00:27.48" resultid="2919" heatid="4669" lane="2" entrytime="00:00:27.00" />
                <RESULT eventid="1157" points="558" swimtime="00:00:37.04" resultid="2920" heatid="4694" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="1393" points="765" swimtime="00:00:59.53" resultid="2921" heatid="4756" lane="4" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1477" points="697" swimtime="00:01:09.70" resultid="2922" heatid="4786" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SWISLE" nation="POL" region="01" clubid="3276" name="Swim Club Masters Ślęza">
          <CONTACT city="Wrocław" email="pawel-chudoba@poczta.fm" name="Chudoba" phone="608623685" state="DOLNO" street="Sowia" zip="53-024" />
          <ATHLETES>
            <ATHLETE firstname="Radosław" lastname="Stefurak" birthdate="1974-09-07" gender="M" nation="POL" athleteid="3277">
              <RESULTS>
                <RESULT eventid="1171" points="450" swimtime="00:00:37.40" resultid="3278" heatid="4700" lane="1" entrytime="00:00:37.87" entrycourse="SCM" />
                <RESULT eventid="1283" points="410" swimtime="00:03:02.26" resultid="3279" heatid="4732" lane="4" entrytime="00:03:01.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                    <SPLIT distance="100" swimtime="00:01:25.23" />
                    <SPLIT distance="150" swimtime="00:02:13.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1589" points="396" swimtime="00:01:24.70" resultid="3280" heatid="4772" lane="1" entrytime="00:01:23.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="357" swimtime="00:01:21.31" resultid="3281" heatid="4790" lane="5" entrytime="00:01:23.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Dusza" birthdate="1983-10-11" gender="F" nation="POL" athleteid="3282">
              <RESULTS>
                <RESULT eventid="1059" points="312" swimtime="00:00:37.02" resultid="3283" heatid="4667" lane="1" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1185" points="334" swimtime="00:02:57.37" resultid="3284" heatid="4707" lane="3" entrytime="00:02:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.53" />
                    <SPLIT distance="100" swimtime="00:01:24.15" />
                    <SPLIT distance="150" swimtime="00:02:10.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="294" swimtime="00:01:22.66" resultid="3285" heatid="4754" lane="2" entrytime="00:01:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1533" points="354" swimtime="00:06:11.06" resultid="3286" heatid="4805" lane="5" entrytime="00:06:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.46" />
                    <SPLIT distance="100" swimtime="00:01:25.17" />
                    <SPLIT distance="150" swimtime="00:02:12.95" />
                    <SPLIT distance="200" swimtime="00:03:01.22" />
                    <SPLIT distance="250" swimtime="00:03:49.02" />
                    <SPLIT distance="300" swimtime="00:04:36.69" />
                    <SPLIT distance="350" swimtime="00:05:24.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03415" nation="POL" region="15" clubid="3549" name="UKS Cityzen Poznań">
          <CONTACT city="Poznań" name="Pietraszewski" phone="501648415" state="WIELK" />
          <ATHLETES>
            <ATHLETE firstname="Jacek" lastname="Matyszczak" birthdate="1970-01-01" gender="M" nation="POL" athleteid="3560">
              <RESULTS>
                <RESULT eventid="1102" points="440" swimtime="00:00:30.74" resultid="3561" heatid="4675" lane="2" entrytime="00:00:30.50" />
                <RESULT eventid="1199" points="319" swimtime="00:02:47.72" resultid="3562" heatid="4711" lane="1" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                    <SPLIT distance="100" swimtime="00:01:19.19" />
                    <SPLIT distance="150" swimtime="00:02:03.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="395" swimtime="00:01:10.15" resultid="3563" heatid="4760" lane="3" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1491" points="338" swimtime="00:01:22.81" resultid="3564" heatid="4789" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zbigniew" lastname="Pietraszewski" birthdate="1955-01-01" gender="M" nation="POL" athleteid="3555">
              <RESULTS>
                <RESULT eventid="1143" points="382" swimtime="00:01:33.27" resultid="3556" heatid="4688" lane="6" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="312" swimtime="00:03:27.02" resultid="3557" heatid="4716" lane="5" entrytime="00:03:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.68" />
                    <SPLIT distance="100" swimtime="00:01:42.17" />
                    <SPLIT distance="150" swimtime="00:02:39.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1435" points="411" swimtime="00:03:22.95" resultid="3558" heatid="4778" lane="1" entrytime="00:03:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.38" />
                    <SPLIT distance="100" swimtime="00:01:38.70" />
                    <SPLIT distance="150" swimtime="00:02:31.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="357" swimtime="00:06:17.59" resultid="3559" heatid="4808" lane="4" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.60" />
                    <SPLIT distance="100" swimtime="00:01:29.51" />
                    <SPLIT distance="150" swimtime="00:02:17.83" />
                    <SPLIT distance="200" swimtime="00:03:05.85" />
                    <SPLIT distance="250" swimtime="00:03:54.15" />
                    <SPLIT distance="300" swimtime="00:04:42.68" />
                    <SPLIT distance="350" swimtime="00:05:31.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Rolewski" birthdate="1967-01-01" gender="M" nation="POL" athleteid="3565">
              <RESULTS>
                <RESULT eventid="1102" points="34" swimtime="00:01:15.13" resultid="3566" heatid="4670" lane="5" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Łutowicz" birthdate="1950-01-01" gender="F" nation="POL" athleteid="3550">
              <RESULTS>
                <RESULT eventid="1059" points="290" swimtime="00:00:48.92" resultid="3551" heatid="4665" lane="3" entrytime="00:00:52.00" />
                <RESULT eventid="1129" points="238" swimtime="00:02:03.53" resultid="3552" heatid="4683" lane="4" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1393" points="261" swimtime="00:01:49.95" resultid="3553" heatid="4752" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1505" points="209" swimtime="00:00:59.25" resultid="3554" heatid="4796" lane="1" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MASZDZ" nation="POL" region="07" clubid="3571" name="MASTERS Zdzieszowice">
          <CONTACT city="Zdzieszowice" email="masters.zdzieszowice@gmail.com" name="Jajuga" phone="505127695" state="OPOLS" street="Fabryczna" zip="47-330" />
          <ATHLETES>
            <ATHLETE firstname="Szymon" lastname="Paciej" birthdate="1988-07-05" gender="M" nation="POL" athleteid="3572">
              <RESULTS>
                <RESULT eventid="1143" status="DNS" swimtime="00:00:00.00" resultid="3573" heatid="4689" lane="6" entrytime="00:01:14.54" />
                <RESULT eventid="1227" status="DNS" swimtime="00:00:00.00" resultid="3574" heatid="4717" lane="6" entrytime="00:02:48.76" />
                <RESULT eventid="1435" status="DNS" swimtime="00:00:00.00" resultid="3575" heatid="4778" lane="4" entrytime="00:02:45.66" />
                <RESULT eventid="1491" status="DNS" swimtime="00:00:00.00" resultid="3576" heatid="4791" lane="2" entrytime="00:01:13.32" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Jajuga" birthdate="1986-02-15" gender="M" nation="POL" athleteid="3577">
              <RESULTS>
                <RESULT eventid="1143" status="DNS" swimtime="00:00:00.00" resultid="3578" heatid="4688" lane="3" entrytime="00:01:15.11" />
                <RESULT eventid="1255" status="DNS" swimtime="00:00:00.00" resultid="3579" heatid="4723" lane="4" entrytime="00:01:06.12" />
                <RESULT eventid="1379" status="DNS" swimtime="00:00:00.00" resultid="3580" heatid="4749" lane="4" entrytime="00:00:28.23" />
                <RESULT eventid="1463" swimtime="00:00:00.00" resultid="3581" entrytime="00:02:40.22" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIERAC" nation="POL" region="11" clubid="2231" name="Zawodnik Niezrzeszony Racibórz" />
        <CLUB type="CLUB" code="5STWAR" nation="POL" region="14" clubid="3614" name="5 Styl Warszawa">
          <CONTACT city="Warszawa" name="Korzeniowski" state="MAZOW" />
          <ATHLETES>
            <ATHLETE firstname="Kuba" lastname="Niedźwiadek" birthdate="1993-10-18" gender="M" nation="POL" athleteid="3619">
              <RESULTS>
                <RESULT eventid="1102" points="375" swimtime="00:00:29.52" resultid="3620" heatid="4677" lane="6" entrytime="00:00:29.00" />
                <RESULT eventid="1199" points="447" swimtime="00:02:17.16" resultid="3621" heatid="4712" lane="2" entrytime="00:02:19.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                    <SPLIT distance="100" swimtime="00:01:06.70" />
                    <SPLIT distance="150" swimtime="00:01:41.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="423" swimtime="00:01:03.20" resultid="3622" heatid="4762" lane="1" entrytime="00:01:04.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="512" swimtime="00:04:51.11" resultid="3623" heatid="4810" lane="1" entrytime="00:05:07.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.14" />
                    <SPLIT distance="100" swimtime="00:01:08.63" />
                    <SPLIT distance="150" swimtime="00:01:45.51" />
                    <SPLIT distance="200" swimtime="00:02:22.55" />
                    <SPLIT distance="250" swimtime="00:02:59.96" />
                    <SPLIT distance="300" swimtime="00:03:37.54" />
                    <SPLIT distance="350" swimtime="00:04:14.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kuba" lastname="Broniszewski" birthdate="1980-09-26" gender="M" nation="POL" athleteid="3615">
              <RESULTS>
                <RESULT eventid="1102" points="275" swimtime="00:00:34.99" resultid="3616" heatid="4671" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="1199" points="253" swimtime="00:02:53.97" resultid="3617" heatid="4710" lane="3" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.10" />
                    <SPLIT distance="100" swimtime="00:01:21.36" />
                    <SPLIT distance="150" swimtime="00:02:07.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="253" swimtime="00:01:18.50" resultid="3618" heatid="4759" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Wziątek" birthdate="1988-01-18" gender="M" nation="POL" athleteid="3629">
              <RESULTS>
                <RESULT eventid="1102" points="311" swimtime="00:00:31.78" resultid="3630" heatid="4674" lane="3" entrytime="00:00:31.11" />
                <RESULT eventid="1491" points="266" swimtime="00:01:22.88" resultid="3631" heatid="4790" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Barnasiuk" birthdate="1992-02-04" gender="M" nation="POL" athleteid="3624">
              <RESULTS>
                <RESULT eventid="1255" points="526" swimtime="00:01:04.98" resultid="3626" heatid="4723" lane="5" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1589" points="572" swimtime="00:01:11.20" resultid="3627" heatid="4774" lane="6" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1463" points="469" swimtime="00:02:26.17" resultid="3628" heatid="4782" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                    <SPLIT distance="100" swimtime="00:01:08.65" />
                    <SPLIT distance="150" swimtime="00:01:47.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="558" swimtime="00:00:32.45" resultid="3833" heatid="4695" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1325" points="415" swimtime="00:04:32.83" resultid="4811" heatid="4736" lane="5" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.71" />
                    <SPLIT distance="100" swimtime="00:00:59.57" />
                    <SPLIT distance="150" swimtime="00:01:32.74" />
                    <SPLIT distance="200" swimtime="00:02:11.94" />
                    <SPLIT distance="250" swimtime="00:02:48.32" />
                    <SPLIT distance="300" swimtime="00:03:28.58" />
                    <SPLIT distance="350" swimtime="00:03:59.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3624" number="1" />
                    <RELAYPOSITION athleteid="3629" number="2" />
                    <RELAYPOSITION athleteid="3615" number="3" />
                    <RELAYPOSITION athleteid="3619" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1350" points="328" swimtime="00:02:22.78" resultid="4812" heatid="4739" lane="6" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.34" />
                    <SPLIT distance="100" swimtime="00:01:24.13" />
                    <SPLIT distance="150" swimtime="00:01:53.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3629" number="1" />
                    <RELAYPOSITION athleteid="3615" number="2" />
                    <RELAYPOSITION athleteid="3624" number="3" />
                    <RELAYPOSITION athleteid="3619" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="COLKRA" nation="POL" region="06" clubid="2324" name="AZS Collegium Medicum UJ Kraków" shortname="AZS Collegium Medicum UJ Krakó">
          <CONTACT city="Kraków" email="karolinaszkudlarek555@gmail.com" name="Szkudlarek Karolina" phone="889018457" state="MAŁOP" />
          <ATHLETES>
            <ATHLETE firstname="Karolina" lastname="Szkudlarek" birthdate="1996-04-04" gender="F" nation="POL" athleteid="2325">
              <RESULTS>
                <RESULT eventid="1185" points="582" swimtime="00:02:22.99" resultid="2326" heatid="4705" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                    <SPLIT distance="100" swimtime="00:01:06.43" />
                    <SPLIT distance="150" swimtime="00:01:44.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1241" points="458" swimtime="00:01:15.36" resultid="2327" heatid="4718" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="534" swimtime="00:00:32.21" resultid="2328" heatid="4743" lane="1" entrytime="00:00:31.55" />
                <RESULT eventid="1393" points="607" swimtime="00:01:04.30" resultid="2329" heatid="4756" lane="5" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIEWRO" nation="POL" region="01" clubid="3016" name="Zawodnik Niezrzeszony Wrocław">
          <ATHLETES>
            <ATHLETE firstname="Łukasz" lastname="Ptak" birthdate="1983-06-07" gender="M" nation="POL" athleteid="3567">
              <RESULTS>
                <RESULT eventid="1171" points="585" swimtime="00:00:31.88" resultid="3568" heatid="4703" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1283" points="645" swimtime="00:02:36.70" resultid="3569" heatid="4733" lane="2" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                    <SPLIT distance="100" swimtime="00:01:15.74" />
                    <SPLIT distance="150" swimtime="00:01:57.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1589" points="621" swimtime="00:01:10.58" resultid="3570" heatid="4774" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Sokulski" birthdate="1991-02-10" gender="M" nation="POL" athleteid="3067">
              <RESULTS>
                <RESULT eventid="1102" points="719" swimtime="00:00:24.03" resultid="3068" heatid="4681" lane="2" entrytime="00:00:24.50" />
                <RESULT eventid="1255" points="744" swimtime="00:00:57.86" resultid="3069" heatid="4724" lane="4" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="778" swimtime="00:00:24.87" resultid="3070" heatid="4751" lane="6" entrytime="00:00:25.50" />
                <RESULT eventid="1407" points="784" swimtime="00:00:51.29" resultid="3071" heatid="4763" lane="3" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Kopacki" birthdate="1998-02-25" gender="M" nation="POL" athleteid="3078">
              <RESULTS>
                <RESULT eventid="1102" swimtime="00:00:23.43" resultid="3079" heatid="4682" lane="3" entrytime="00:00:23.00" />
                <RESULT eventid="1379" swimtime="00:00:26.34" resultid="3080" heatid="4751" lane="5" entrytime="00:00:25.50" />
                <RESULT eventid="1407" swimtime="00:00:51.47" resultid="3081" heatid="4764" lane="3" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Picher" birthdate="1983-02-05" gender="M" nation="POL" athleteid="3075">
              <RESULTS>
                <RESULT eventid="1102" points="289" swimtime="00:00:32.57" resultid="3076" heatid="4674" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="1379" points="289" swimtime="00:00:34.96" resultid="3077" heatid="4745" lane="4" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Bołtuć" birthdate="1983-06-13" gender="F" nation="POL" athleteid="3017">
              <RESULTS>
                <RESULT eventid="1185" points="424" swimtime="00:02:43.86" resultid="3018" heatid="4707" lane="4" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                    <SPLIT distance="100" swimtime="00:01:21.92" />
                    <SPLIT distance="150" swimtime="00:02:03.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="325" swimtime="00:03:20.22" resultid="3019" heatid="4715" lane="6" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.06" />
                    <SPLIT distance="100" swimtime="00:01:37.89" />
                    <SPLIT distance="150" swimtime="00:02:35.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1477" points="276" swimtime="00:01:37.08" resultid="3020" heatid="4784" lane="1" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1533" points="444" swimtime="00:05:44.15" resultid="3021" heatid="4805" lane="4" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.94" />
                    <SPLIT distance="100" swimtime="00:01:22.79" />
                    <SPLIT distance="150" swimtime="00:02:06.26" />
                    <SPLIT distance="200" swimtime="00:02:50.12" />
                    <SPLIT distance="250" swimtime="00:03:34.00" />
                    <SPLIT distance="300" swimtime="00:04:18.21" />
                    <SPLIT distance="350" swimtime="00:05:02.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIECHO" nation="POL" region="11" clubid="3236" name="Zawodnik Niezrzeszony Chorzów">
          <ATHLETES>
            <ATHLETE firstname="Dominik" lastname="Rudzki" birthdate="1992-06-21" gender="M" nation="POL" athleteid="3238">
              <RESULTS>
                <RESULT eventid="1171" points="490" swimtime="00:00:33.89" resultid="3239" heatid="4702" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="1227" points="480" swimtime="00:02:29.35" resultid="3240" heatid="4717" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.37" />
                    <SPLIT distance="100" swimtime="00:01:08.46" />
                    <SPLIT distance="150" swimtime="00:01:52.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1283" points="486" swimtime="00:02:46.89" resultid="3241" heatid="4733" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                    <SPLIT distance="100" swimtime="00:01:16.75" />
                    <SPLIT distance="150" swimtime="00:02:00.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1589" points="493" swimtime="00:01:14.83" resultid="3242" heatid="4772" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NIESOK" nation="POL" region="14" clubid="3062" name="Zawodnik Niezrzeszony Sokołów Podlaski">
          <CONTACT name="Zawodnik Niezrzeszony Sokołów Podlaski" />
          <ATHLETES>
            <ATHLETE firstname="Aneta" lastname="Dolińska" birthdate="1990-07-06" gender="F" nation="POL" athleteid="3063">
              <RESULTS>
                <RESULT eventid="1059" points="426" swimtime="00:00:33.44" resultid="3064" heatid="4667" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="1477" points="333" swimtime="00:01:30.19" resultid="3065" heatid="4784" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1505" points="264" swimtime="00:00:42.76" resultid="3066" heatid="4797" lane="6" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00701" nation="POL" region="01" clubid="2527" name="MKS Dziewiątka Dzierżoniów">
          <CONTACT city="Dzierżoniów" email="ewajuraszek99@op.pl" name="Wojtal Andrzej" phone="508509429" state="DOLNO" street="Sienkiewicza 13" zip="58-200" />
          <ATHLETES>
            <ATHLETE firstname="Zuzanna" lastname="Pisarska" birthdate="1981-06-11" gender="F" nation="POL" license="100701600113" athleteid="2533">
              <RESULTS>
                <RESULT eventid="1059" points="802" swimtime="00:00:28.01" resultid="2534" heatid="4669" lane="1" entrytime="00:00:27.92" entrycourse="SCM" />
                <RESULT eventid="1129" points="699" swimtime="00:01:11.23" resultid="2535" heatid="4685" lane="3" entrytime="00:01:09.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="847" swimtime="00:00:29.79" resultid="2536" heatid="4743" lane="2" entrytime="00:00:29.60" entrycourse="SCM" />
                <RESULT eventid="1505" points="776" swimtime="00:00:31.40" resultid="2537" heatid="4798" lane="3" entrytime="00:00:32.67" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edyta" lastname="Bejster" birthdate="1981-05-21" gender="F" nation="POL" license="100701600124" athleteid="2538">
              <RESULTS>
                <RESULT eventid="1059" points="285" swimtime="00:00:39.56" resultid="2539" heatid="4666" lane="4" entrytime="00:00:38.50" entrycourse="SCM" />
                <RESULT eventid="1157" points="251" swimtime="00:00:50.97" resultid="2540" heatid="4692" lane="2" entrytime="00:00:48.23" entrycourse="SCM" />
                <RESULT eventid="1575" points="259" swimtime="00:01:49.70" resultid="2541" heatid="4766" lane="1" entrytime="00:01:56.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1477" points="222" swimtime="00:01:46.03" resultid="2542" heatid="4784" lane="6" entrytime="00:01:46.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrianna" lastname="Falkowska" birthdate="1982-03-11" gender="F" nation="POL" license="100701600120" athleteid="2543">
              <RESULTS>
                <RESULT eventid="1059" points="176" swimtime="00:00:46.42" resultid="2544" heatid="4664" lane="2" />
                <RESULT eventid="1157" points="204" swimtime="00:00:54.64" resultid="2545" heatid="4691" lane="5" />
                <RESULT eventid="1575" points="193" swimtime="00:02:01.14" resultid="2546" heatid="4765" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1505" points="147" swimtime="00:00:54.70" resultid="2547" heatid="4795" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Kuszka" birthdate="1977-04-14" gender="M" nation="POL" license="100701700110" athleteid="2528">
              <RESULTS>
                <RESULT eventid="1171" points="322" swimtime="00:00:41.80" resultid="2529" heatid="4697" lane="1" entrytime="00:00:45.00" entrycourse="SCM" />
                <RESULT eventid="1255" points="196" swimtime="00:01:34.75" resultid="2530" heatid="4720" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="282" swimtime="00:00:37.16" resultid="2531" heatid="4744" lane="4" entrytime="00:00:40.20" entrycourse="SCM" />
                <RESULT eventid="1491" points="257" swimtime="00:01:30.75" resultid="2532" heatid="4788" lane="3" entrytime="00:01:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>

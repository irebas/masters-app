<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Dolnoslaski Okregowy Zwiazek Plywacki" version="11.74191">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Bielawa" name="XVII MISTRZOSTWA  DOLNEGO  ŚLĄSKA w PŁYWANIU  MASTERS, PUCHAR POLSKI MASTERS" course="SCM" number="1" organizer="Ośrodek Sportu i Rekreacji w Bielawie" organizer.url="http://www.osir.bielawa.pl" reservecount="2" result.url="http://www.megatiming.pl" startmethod="1" timing="AUTOMATIC" nation="POL" maxentriesathlete="99" maxentriesrelay="99">
      <AGEDATE value="2023-01-01" type="YEAR" />
      <POOL name="PŁYWALNIA AQUARIUS" lanemin="1" lanemax="6" />
      <FACILITY city="Bielawa" name="PŁYWALNIA AQUARIUS" nation="POL" />
      <POINTTABLE pointtableid="1126" name="DSV Master Performance Table" version="2022" />
      <CONTACT email="szewczyk@osir.bielawa.pl" name="Czesław Szewczyk " phone="519 331 161" />
      <FEES>
        <FEE currency="PLN" type="ATHLETE" value="8000" />
        <FEE currency="PLN" type="LATEENTRY.INDIVIDUAL" value="8000" />
      </FEES>
      <QUALIFY from="2020-01-01" until="2023-04-08" />
      <SESSIONS>
        <SESSION date="2023-04-15" daytime="15:00" endtime="17:58" name="BLOK I" number="1" officialmeeting="12:00" teamleadermeeting="12:00" warmupfrom="13:30" warmupuntil="14:30" maxentriesathlete="3" maxentriesrelay="3">
          <EVENTS>
            <EVENT eventid="1053" daytime="15:00" gender="F" number="1" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2245" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14714" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2246" agemax="34" agemin="30" name="Kategoria B" />
                <AGEGROUP agegroupid="2247" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15049" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2248" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15304" />
                    <RANKING order="2" place="2" resultid="15162" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2249" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15165" />
                    <RANKING order="2" place="2" resultid="15157" />
                    <RANKING order="3" place="3" resultid="15103" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2250" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14723" />
                    <RANKING order="2" place="2" resultid="15100" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2251" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14559" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2252" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14790" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2253" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14785" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2254" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15108" />
                    <RANKING order="2" place="2" resultid="15507" />
                    <RANKING order="3" place="3" resultid="14852" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2255" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2256" agemax="84" agemin="80" name="Kategoria L" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15549" daytime="15:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15550" daytime="15:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="15551" daytime="15:10" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1066" daytime="15:18" gender="M" number="2" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3077" agemax="29" agemin="25" name="Kategoria A" />
                <AGEGROUP agegroupid="3078" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15193" />
                    <RANKING order="2" place="2" resultid="15021" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3079" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14689" />
                    <RANKING order="2" place="2" resultid="14534" />
                    <RANKING order="3" place="3" resultid="14824" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3080" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15769" />
                    <RANKING order="2" place="2" resultid="15178" />
                    <RANKING order="3" place="3" resultid="15276" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3081" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15706" />
                    <RANKING order="2" place="2" resultid="15321" />
                    <RANKING order="3" place="3" resultid="15702" />
                    <RANKING order="4" place="4" resultid="14977" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3082" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15151" />
                    <RANKING order="2" place="2" resultid="14738" />
                    <RANKING order="3" place="3" resultid="15452" />
                    <RANKING order="4" place="-1" resultid="15054" />
                    <RANKING order="5" place="-1" resultid="15188" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3083" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15059" />
                    <RANKING order="2" place="2" resultid="15003" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3084" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15113" />
                    <RANKING order="2" place="2" resultid="15064" />
                    <RANKING order="3" place="3" resultid="15183" />
                    <RANKING order="4" place="4" resultid="15091" />
                    <RANKING order="5" place="5" resultid="14746" />
                    <RANKING order="6" place="6" resultid="15174" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3085" agemax="69" agemin="65" name="Kategoria I" />
                <AGEGROUP agegroupid="3086" agemax="74" agemin="70" name="Kategoria J" />
                <AGEGROUP agegroupid="3087" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15170" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8905" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14593" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3088" agemax="89" agemin="85" name="Kategoria M" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15552" daytime="15:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15553" daytime="15:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="15554" daytime="15:26" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="15555" daytime="15:32" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="15556" daytime="15:36" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1079" daytime="15:42" gender="F" number="3" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3089" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15037" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3090" agemax="34" agemin="30" name="Kategoria B" />
                <AGEGROUP agegroupid="3091" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15309" />
                    <RANKING order="2" place="2" resultid="14802" />
                    <RANKING order="3" place="3" resultid="14758" />
                    <RANKING order="4" place="4" resultid="15050" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3092" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15145" />
                    <RANKING order="2" place="2" resultid="14662" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3093" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15673" />
                    <RANKING order="2" place="2" resultid="14679" />
                    <RANKING order="3" place="3" resultid="15207" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3094" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14857" />
                    <RANKING order="2" place="2" resultid="15735" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3095" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15202" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3096" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15197" />
                    <RANKING order="2" place="-1" resultid="14875" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3097" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14847" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3098" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15512" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3099" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15502" />
                    <RANKING order="2" place="2" resultid="15488" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3100" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15485" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15557" daytime="15:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15558" daytime="15:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="15559" daytime="15:44" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="15560" daytime="15:46" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1092" daytime="15:48" gender="M" number="4" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="8907" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15315" />
                    <RANKING order="2" place="2" resultid="14658" />
                    <RANKING order="3" place="3" resultid="15226" />
                    <RANKING order="4" place="4" resultid="14515" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8908" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15096" />
                    <RANKING order="2" place="2" resultid="15475" />
                    <RANKING order="3" place="3" resultid="14797" />
                    <RANKING order="4" place="4" resultid="14615" />
                    <RANKING order="5" place="-1" resultid="14599" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8909" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15471" />
                    <RANKING order="2" place="2" resultid="14684" />
                    <RANKING order="3" place="3" resultid="15222" />
                    <RANKING order="4" place="4" resultid="14761" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8910" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14522" />
                    <RANKING order="2" place="2" resultid="15129" />
                    <RANKING order="3" place="3" resultid="15714" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8911" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15522" />
                    <RANKING order="2" place="2" resultid="14611" />
                    <RANKING order="3" place="3" resultid="15132" />
                    <RANKING order="4" place="4" resultid="15694" />
                    <RANKING order="5" place="5" resultid="14810" />
                    <RANKING order="6" place="6" resultid="14806" />
                    <RANKING order="7" place="7" resultid="15279" />
                    <RANKING order="8" place="-1" resultid="14819" />
                    <RANKING order="9" place="-1" resultid="15217" />
                    <RANKING order="10" place="-1" resultid="15728" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8912" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15136" />
                    <RANKING order="2" place="2" resultid="14775" />
                    <RANKING order="3" place="3" resultid="15730" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8913" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15212" />
                    <RANKING order="2" place="2" resultid="15288" />
                    <RANKING order="3" place="3" resultid="14733" />
                    <RANKING order="4" place="4" resultid="15724" />
                    <RANKING order="5" place="-1" resultid="15719" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8914" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15326" />
                    <RANKING order="2" place="2" resultid="14564" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8915" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14540" />
                    <RANKING order="2" place="2" resultid="15283" />
                    <RANKING order="3" place="3" resultid="14867" />
                    <RANKING order="4" place="4" resultid="15031" />
                    <RANKING order="5" place="5" resultid="15492" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8916" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14842" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8917" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14605" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8918" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14872" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8919" agemax="89" agemin="85" name="Kategoria M" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15561" daytime="15:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15562" daytime="15:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="15563" daytime="15:52" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="15564" daytime="15:54" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="15565" daytime="15:54" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="15566" daytime="15:56" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="15567" daytime="15:58" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="15568" daytime="16:00" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1105" daytime="16:02" gender="F" number="5" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3113" agemax="29" agemin="25" name="Kategoria A" />
                <AGEGROUP agegroupid="3114" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15676" />
                    <RANKING order="2" place="2" resultid="14728" />
                    <RANKING order="3" place="3" resultid="14752" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3115" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15664" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3116" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15069" />
                    <RANKING order="2" place="2" resultid="14677" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3117" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="15208" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3118" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15009" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3119" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15203" />
                    <RANKING order="2" place="2" resultid="15123" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3120" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15118" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3121" agemax="69" agemin="65" name="Kategoria I" />
                <AGEGROUP agegroupid="3122" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14862" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3123" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15503" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3124" agemax="84" agemin="80" name="Kategoria L" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15569" daytime="16:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15570" daytime="16:06" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="15571" daytime="16:10" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1118" daytime="16:14" gender="M" number="6" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="8920" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14990" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8921" agemax="34" agemin="30" name="Kategoria B" />
                <AGEGROUP agegroupid="8922" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15710" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8923" agemax="44" agemin="40" name="Kategoria D" />
                <AGEGROUP agegroupid="8924" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15236" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8925" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15043" />
                    <RANKING order="2" place="2" resultid="14708" />
                    <RANKING order="3" place="3" resultid="14510" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8926" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15331" />
                    <RANKING order="2" place="2" resultid="15015" />
                    <RANKING order="3" place="3" resultid="15497" />
                    <RANKING order="4" place="4" resultid="15025" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8927" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14693" />
                    <RANKING order="2" place="-1" resultid="15293" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8928" agemax="69" agemin="65" name="Kategoria I" />
                <AGEGROUP agegroupid="8929" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14578" />
                    <RANKING order="2" place="2" resultid="14769" />
                    <RANKING order="3" place="3" resultid="15231" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8930" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14588" />
                    <RANKING order="2" place="2" resultid="15480" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8931" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="8932" agemax="89" agemin="85" name="Kategoria M" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15572" daytime="16:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15573" daytime="16:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="15574" daytime="16:20" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1131" daytime="16:24" gender="F" number="7" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3137" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15038" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3138" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15677" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3139" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15665" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3140" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15146" />
                    <RANKING order="2" place="2" resultid="15241" />
                    <RANKING order="3" place="3" resultid="15690" />
                    <RANKING order="4" place="4" resultid="15305" />
                    <RANKING order="5" place="5" resultid="15163" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3141" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15674" />
                    <RANKING order="2" place="2" resultid="15104" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3142" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15246" />
                    <RANKING order="2" place="2" resultid="15074" />
                    <RANKING order="3" place="3" resultid="15669" />
                    <RANKING order="4" place="4" resultid="15250" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3143" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15079" />
                    <RANKING order="2" place="2" resultid="14560" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3144" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15198" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3145" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14848" />
                    <RANKING order="2" place="2" resultid="14780" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3146" agemax="74" agemin="70" name="Kategoria J" />
                <AGEGROUP agegroupid="3147" agemax="79" agemin="75" name="Kategoria K" />
                <AGEGROUP agegroupid="3148" agemax="84" agemin="80" name="Kategoria L" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15575" daytime="16:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15576" daytime="16:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="15577" daytime="16:28" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="15578" daytime="16:30" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1144" daytime="16:32" gender="M" number="8" order="8" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="8933" agemax="29" agemin="25" name="Kategoria A" />
                <AGEGROUP agegroupid="8934" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14814" />
                    <RANKING order="2" place="2" resultid="14799" />
                    <RANKING order="3" place="3" resultid="14616" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8935" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15740" />
                    <RANKING order="2" place="2" resultid="14685" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8936" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14701" />
                    <RANKING order="2" place="2" resultid="14573" />
                    <RANKING order="3" place="3" resultid="15698" />
                    <RANKING order="4" place="4" resultid="15300" />
                    <RANKING order="5" place="5" resultid="15000" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8937" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14808" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8938" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15044" />
                    <RANKING order="2" place="2" resultid="15055" />
                    <RANKING order="3" place="3" resultid="15451" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8939" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15213" />
                    <RANKING order="2" place="2" resultid="14528" />
                    <RANKING order="3" place="3" resultid="15725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8940" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15294" />
                    <RANKING order="2" place="-1" resultid="14980" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8941" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15255" />
                    <RANKING order="2" place="2" resultid="15284" />
                    <RANKING order="3" place="3" resultid="14546" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8942" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14843" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8943" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14589" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8944" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14873" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8945" agemax="89" agemin="85" name="Kategoria M" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15579" daytime="16:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15580" daytime="16:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="15581" daytime="16:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="15582" daytime="16:36" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="15583" daytime="16:38" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1157" daytime="16:40" gender="F" number="9" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3161" agemax="29" agemin="25" name="Kategoria A" />
                <AGEGROUP agegroupid="3162" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15764" />
                    <RANKING order="2" place="2" resultid="14729" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3163" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14803" />
                    <RANKING order="2" place="2" resultid="14759" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3164" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15467" />
                    <RANKING order="2" place="2" resultid="14984" />
                    <RANKING order="3" place="3" resultid="15242" />
                    <RANKING order="4" place="4" resultid="14969" />
                    <RANKING order="5" place="-1" resultid="15685" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3165" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14680" />
                    <RANKING order="2" place="2" resultid="15158" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3166" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14858" />
                    <RANKING order="2" place="2" resultid="15670" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3167" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15124" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3168" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15119" />
                    <RANKING order="2" place="2" resultid="15084" />
                    <RANKING order="3" place="-1" resultid="14876" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3169" agemax="69" agemin="65" name="Kategoria I" />
                <AGEGROUP agegroupid="3170" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14863" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3171" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14584" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3172" agemax="84" agemin="80" name="Kategoria L" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15584" daytime="16:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15585" daytime="16:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="15586" daytime="16:48" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="15587" daytime="16:54" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1170" daytime="17:00" gender="M" number="10" order="10" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="8946" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14659" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8947" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14815" />
                    <RANKING order="2" place="2" resultid="15022" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8948" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15741" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8949" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15770" />
                    <RANKING order="2" place="2" resultid="15130" />
                    <RANKING order="3" place="3" resultid="15715" />
                    <RANKING order="4" place="4" resultid="15277" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8950" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14811" />
                    <RANKING order="2" place="2" resultid="15280" />
                    <RANKING order="3" place="-1" resultid="14820" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8951" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15137" />
                    <RANKING order="2" place="2" resultid="14776" />
                    <RANKING order="3" place="3" resultid="15446" />
                    <RANKING order="4" place="4" resultid="14974" />
                    <RANKING order="5" place="5" resultid="14709" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8952" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15026" />
                    <RANKING order="2" place="2" resultid="15004" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8953" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14694" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8954" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14868" />
                    <RANKING order="2" place="2" resultid="15032" />
                    <RANKING order="3" place="3" resultid="14547" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8955" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14579" />
                    <RANKING order="2" place="2" resultid="14765" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8956" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14606" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8957" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="8958" agemax="89" agemin="85" name="Kategoria M" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15588" daytime="17:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15589" daytime="17:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="15590" daytime="17:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="15591" daytime="17:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="15592" daytime="17:16" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5376" daytime="17:20" gender="F" number="11" order="11" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5377" agemax="29" agemin="25" name="Kategoria A" />
                <AGEGROUP agegroupid="5378" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15765" />
                    <RANKING order="2" place="2" resultid="14753" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5379" agemax="39" agemin="35" name="Kategoria C" />
                <AGEGROUP agegroupid="5380" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15070" />
                    <RANKING order="2" place="2" resultid="14985" />
                    <RANKING order="3" place="3" resultid="14663" />
                    <RANKING order="4" place="4" resultid="15691" />
                    <RANKING order="5" place="-1" resultid="15686" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5381" agemax="49" agemin="45" name="Kategoria E" />
                <AGEGROUP agegroupid="5382" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15247" />
                    <RANKING order="2" place="2" resultid="15010" />
                    <RANKING order="3" place="3" resultid="15736" />
                    <RANKING order="4" place="4" resultid="15251" />
                    <RANKING order="5" place="5" resultid="15075" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5383" agemax="59" agemin="55" name="Kategoria G" />
                <AGEGROUP agegroupid="5384" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15085" />
                    <RANKING order="2" place="2" resultid="14791" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5385" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14781" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5386" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15513" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5387" agemax="79" agemin="75" name="Kategoria K" />
                <AGEGROUP agegroupid="5388" agemax="84" agemin="80" name="Kategoria L" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15593" daytime="17:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15594" daytime="17:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="15595" daytime="17:26" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5390" daytime="17:30" gender="M" number="12" order="12" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="8959" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15316" />
                    <RANKING order="2" place="2" resultid="14516" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8960" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15476" />
                    <RANKING order="2" place="-1" resultid="14600" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8961" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15223" />
                    <RANKING order="2" place="2" resultid="14825" />
                    <RANKING order="3" place="3" resultid="14762" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8962" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14572" />
                    <RANKING order="2" place="2" resultid="15699" />
                    <RANKING order="3" place="3" resultid="15301" />
                    <RANKING order="4" place="4" resultid="15001" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8963" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15707" />
                    <RANKING order="2" place="2" resultid="15523" />
                    <RANKING order="3" place="3" resultid="15237" />
                    <RANKING order="4" place="4" resultid="15133" />
                    <RANKING order="5" place="5" resultid="14978" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8964" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15447" />
                    <RANKING order="2" place="2" resultid="14975" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8965" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15332" />
                    <RANKING order="2" place="2" resultid="15016" />
                    <RANKING order="3" place="3" resultid="15720" />
                    <RANKING order="4" place="4" resultid="14529" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8966" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15295" />
                    <RANKING order="2" place="2" resultid="15327" />
                    <RANKING order="3" place="3" resultid="14565" />
                    <RANKING order="4" place="4" resultid="15184" />
                    <RANKING order="5" place="5" resultid="15065" />
                    <RANKING order="6" place="6" resultid="14981" />
                    <RANKING order="7" place="-1" resultid="14747" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8967" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15256" />
                    <RANKING order="2" place="2" resultid="15260" />
                    <RANKING order="3" place="3" resultid="14541" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8968" agemax="74" agemin="70" name="Kategoria J" />
                <AGEGROUP agegroupid="8969" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15481" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8970" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="8971" agemax="89" agemin="85" name="Kategoria M" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15596" daytime="17:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15597" daytime="17:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="15598" daytime="17:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="15599" daytime="17:38" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="15600" daytime="17:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="15601" daytime="17:44" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1183" daytime="17:46" gender="F" number="13" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6832" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14715" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6833" agemax="34" agemin="30" name="Kategoria B" />
                <AGEGROUP agegroupid="6834" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15310" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6835" agemax="44" agemin="40" name="Kategoria D" />
                <AGEGROUP agegroupid="6836" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15166" />
                    <RANKING order="2" place="2" resultid="15681" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6837" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14724" />
                    <RANKING order="2" place="2" resultid="15101" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6838" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15080" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6839" agemax="64" agemin="60" name="Kategoria H" />
                <AGEGROUP agegroupid="6840" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14786" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6841" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15109" />
                    <RANKING order="2" place="2" resultid="14853" />
                    <RANKING order="3" place="3" resultid="15508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6842" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15489" />
                    <RANKING order="2" place="2" resultid="14556" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6843" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15486" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15602" daytime="17:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15603" daytime="17:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="15604" daytime="17:50" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6830" daytime="17:52" gender="M" number="14" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="8972" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15227" />
                    <RANKING order="2" place="2" resultid="14991" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8973" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15097" />
                    <RANKING order="2" place="2" resultid="15194" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8974" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14535" />
                    <RANKING order="2" place="2" resultid="14690" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8975" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14702" />
                    <RANKING order="2" place="2" resultid="15141" />
                    <RANKING order="3" place="3" resultid="14523" />
                    <RANKING order="4" place="4" resultid="15179" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8976" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15322" />
                    <RANKING order="2" place="2" resultid="15703" />
                    <RANKING order="3" place="-1" resultid="15695" />
                    <RANKING order="4" place="-1" resultid="15218" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8977" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15152" />
                    <RANKING order="2" place="2" resultid="15189" />
                    <RANKING order="3" place="3" resultid="14739" />
                    <RANKING order="4" place="4" resultid="14519" />
                    <RANKING order="5" place="-1" resultid="15731" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8978" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15498" />
                    <RANKING order="2" place="2" resultid="14772" />
                    <RANKING order="3" place="3" resultid="15060" />
                    <RANKING order="4" place="4" resultid="14734" />
                    <RANKING order="5" place="5" resultid="15289" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8979" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15114" />
                    <RANKING order="2" place="2" resultid="15092" />
                    <RANKING order="3" place="3" resultid="15175" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8980" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15261" />
                    <RANKING order="2" place="2" resultid="15493" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8981" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15232" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8982" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15171" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8983" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14594" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8984" agemax="89" agemin="85" name="Kategoria M" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15605" daytime="17:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15606" daytime="17:54" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="15607" daytime="17:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="15608" daytime="17:58" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="15609" daytime="18:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="15610" daytime="18:02" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6828" daytime="18:04" gender="X" number="15" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6829" agemax="-1" agemin="-1" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15742" />
                    <RANKING order="2" place="2" resultid="15745" />
                    <RANKING order="3" place="3" resultid="15088" />
                    <RANKING order="4" place="4" resultid="14697" />
                    <RANKING order="5" place="5" resultid="15266" />
                    <RANKING order="6" place="6" resultid="15264" />
                    <RANKING order="7" place="7" resultid="15265" />
                    <RANKING order="8" place="8" resultid="15268" />
                    <RANKING order="9" place="9" resultid="14744" />
                    <RANKING order="10" place="10" resultid="15744" />
                    <RANKING order="11" place="11" resultid="14794" />
                    <RANKING order="12" place="-1" resultid="15267" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15611" daytime="18:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15612" daytime="18:06" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2023-04-16" daytime="10:00" endtime="13:47" name="BLOK II" number="2" warmupfrom="09:20" warmupuntil="09:50" maxentriesathlete="3">
          <EVENTS>
            <EVENT eventid="5430" daytime="10:00" gender="F" number="16" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5431" agemax="29" agemin="25" name="Kategoria A" />
                <AGEGROUP agegroupid="5432" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15766" />
                    <RANKING order="2" place="2" resultid="14754" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5433" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15666" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5434" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15071" />
                    <RANKING order="2" place="2" resultid="14986" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5435" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15209" />
                    <RANKING order="2" place="2" resultid="15159" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5436" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15011" />
                    <RANKING order="2" place="2" resultid="15076" />
                    <RANKING order="3" place="3" resultid="15252" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5437" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15125" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5438" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15120" />
                    <RANKING order="2" place="2" resultid="14792" />
                    <RANKING order="3" place="-1" resultid="14877" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5439" agemax="69" agemin="65" name="Kategoria I" />
                <AGEGROUP agegroupid="5440" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14864" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5441" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15504" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5442" agemax="84" agemin="80" name="Kategoria L" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15614" daytime="10:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15615" daytime="10:06" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="15616" daytime="10:14" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5443" daytime="10:20" gender="M" number="17" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="8985" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14517" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8986" agemax="34" agemin="30" name="Kategoria B" />
                <AGEGROUP agegroupid="8987" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15711" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8988" agemax="44" agemin="40" name="Kategoria D" />
                <AGEGROUP agegroupid="8989" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15524" />
                    <RANKING order="2" place="2" resultid="15238" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8990" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15045" />
                    <RANKING order="2" place="2" resultid="15448" />
                    <RANKING order="3" place="3" resultid="14511" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8991" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15017" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8992" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15296" />
                    <RANKING order="2" place="2" resultid="14695" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8993" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14869" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8994" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14766" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8995" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15482" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8996" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="8997" agemax="89" agemin="85" name="Kategoria M" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15617" daytime="10:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15618" daytime="10:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="15619" daytime="10:32" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1198" daytime="10:38" gender="F" number="18" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3185" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14716" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3186" agemax="34" agemin="30" name="Kategoria B" />
                <AGEGROUP agegroupid="3187" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15311" />
                    <RANKING order="2" place="-1" resultid="15051" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3188" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14987" />
                    <RANKING order="2" place="2" resultid="15243" />
                    <RANKING order="3" place="3" resultid="15306" />
                    <RANKING order="4" place="4" resultid="14970" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3189" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14681" />
                    <RANKING order="2" place="2" resultid="15167" />
                    <RANKING order="3" place="3" resultid="15682" />
                    <RANKING order="4" place="4" resultid="15105" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3190" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14859" />
                    <RANKING order="2" place="2" resultid="14725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3191" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14561" />
                    <RANKING order="2" place="-1" resultid="15081" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3192" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14793" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3193" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14787" />
                    <RANKING order="2" place="2" resultid="14849" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3194" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15110" />
                    <RANKING order="2" place="2" resultid="15509" />
                    <RANKING order="3" place="3" resultid="14854" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3195" agemax="79" agemin="75" name="Kategoria K" />
                <AGEGROUP agegroupid="3196" agemax="84" agemin="80" name="Kategoria L" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15620" daytime="10:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15621" daytime="10:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="15622" daytime="10:44" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="15623" daytime="10:46" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1212" daytime="10:50" gender="M" number="19" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="8998" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15228" />
                    <RANKING order="2" place="2" resultid="14993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8999" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15195" />
                    <RANKING order="2" place="2" resultid="14601" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9000" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14536" />
                    <RANKING order="2" place="2" resultid="14691" />
                    <RANKING order="3" place="3" resultid="14826" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9001" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14703" />
                    <RANKING order="2" place="2" resultid="15142" />
                    <RANKING order="3" place="3" resultid="15771" />
                    <RANKING order="4" place="4" resultid="14524" />
                    <RANKING order="5" place="5" resultid="15180" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9002" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15323" />
                    <RANKING order="2" place="2" resultid="15704" />
                    <RANKING order="3" place="3" resultid="14972" />
                    <RANKING order="4" place="-1" resultid="15219" />
                    <RANKING order="5" place="-1" resultid="15708" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9003" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15153" />
                    <RANKING order="2" place="2" resultid="15056" />
                    <RANKING order="3" place="3" resultid="14740" />
                    <RANKING order="4" place="4" resultid="15190" />
                    <RANKING order="5" place="-1" resultid="15454" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9004" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15499" />
                    <RANKING order="2" place="2" resultid="15061" />
                    <RANKING order="3" place="3" resultid="14735" />
                    <RANKING order="4" place="4" resultid="14530" />
                    <RANKING order="5" place="5" resultid="15290" />
                    <RANKING order="6" place="-1" resultid="15214" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9005" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15328" />
                    <RANKING order="2" place="2" resultid="15115" />
                    <RANKING order="3" place="3" resultid="15093" />
                    <RANKING order="4" place="4" resultid="15066" />
                    <RANKING order="5" place="5" resultid="15176" />
                    <RANKING order="6" place="-1" resultid="15185" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9006" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15262" />
                    <RANKING order="2" place="2" resultid="15494" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9007" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="15233" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9008" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15172" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9009" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14595" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9010" agemax="89" agemin="85" name="Kategoria M" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15624" daytime="10:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15625" daytime="10:52" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="15626" daytime="10:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="15627" daytime="10:58" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="15628" daytime="11:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="15629" daytime="11:04" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="15630" daytime="11:08" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1303" daytime="11:12" gender="F" number="20" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3281" agemax="29" agemin="25" name="Kategoria A" />
                <AGEGROUP agegroupid="3282" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15678" />
                    <RANKING order="2" place="2" resultid="14730" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3283" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15312" />
                    <RANKING order="2" place="2" resultid="15052" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3284" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15147" />
                    <RANKING order="2" place="2" resultid="15072" />
                    <RANKING order="3" place="3" resultid="15307" />
                    <RANKING order="4" place="4" resultid="14664" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3285" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15168" />
                    <RANKING order="2" place="2" resultid="15210" />
                    <RANKING order="3" place="3" resultid="15683" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3286" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15737" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3287" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15204" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3288" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15086" />
                    <RANKING order="2" place="2" resultid="15199" />
                    <RANKING order="3" place="-1" resultid="14878" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3289" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14782" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3290" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14855" />
                    <RANKING order="2" place="2" resultid="15510" />
                    <RANKING order="3" place="3" resultid="15514" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3291" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15505" />
                    <RANKING order="2" place="2" resultid="14585" />
                    <RANKING order="3" place="3" resultid="15490" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3292" agemax="84" agemin="80" name="Kategoria L" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15631" daytime="11:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15632" daytime="11:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="15633" daytime="11:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="15634" daytime="11:20" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1316" daytime="11:24" gender="M" number="21" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9011" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15317" />
                    <RANKING order="2" place="2" resultid="14992" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9012" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14602" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9013" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15712" />
                    <RANKING order="2" place="2" resultid="14686" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9014" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15716" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9015" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15696" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9016" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15138" />
                    <RANKING order="2" place="2" resultid="15057" />
                    <RANKING order="3" place="3" resultid="14777" />
                    <RANKING order="4" place="4" resultid="14741" />
                    <RANKING order="5" place="5" resultid="14512" />
                    <RANKING order="6" place="-1" resultid="15732" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9017" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15018" />
                    <RANKING order="2" place="2" resultid="15333" />
                    <RANKING order="3" place="3" resultid="15721" />
                    <RANKING order="4" place="4" resultid="15500" />
                    <RANKING order="5" place="5" resultid="14773" />
                    <RANKING order="6" place="6" resultid="15027" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9018" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15116" />
                    <RANKING order="2" place="-1" resultid="15297" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9019" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15257" />
                    <RANKING order="2" place="2" resultid="15263" />
                    <RANKING order="3" place="3" resultid="14542" />
                    <RANKING order="4" place="4" resultid="15285" />
                    <RANKING order="5" place="5" resultid="15033" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9020" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14580" />
                    <RANKING order="2" place="2" resultid="14767" />
                    <RANKING order="3" place="3" resultid="14844" />
                    <RANKING order="4" place="4" resultid="14770" />
                    <RANKING order="5" place="-1" resultid="15234" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9021" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14590" />
                    <RANKING order="2" place="2" resultid="14607" />
                    <RANKING order="3" place="3" resultid="15483" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9022" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="9023" agemax="89" agemin="85" name="Kategoria M" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15635" daytime="11:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15636" daytime="11:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="15637" daytime="11:28" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="15638" daytime="11:32" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="15639" daytime="11:34" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="15640" daytime="11:38" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5404" daytime="11:40" gender="F" number="22" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5405" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15039" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5406" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15679" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5407" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15667" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5408" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15148" />
                    <RANKING order="2" place="-1" resultid="15687" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5409" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15160" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5410" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15248" />
                    <RANKING order="2" place="2" resultid="15012" />
                    <RANKING order="3" place="3" resultid="15077" />
                    <RANKING order="4" place="4" resultid="15253" />
                    <RANKING order="5" place="-1" resultid="15738" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5411" agemax="59" agemin="55" name="Kategoria G" />
                <AGEGROUP agegroupid="5412" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15087" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5413" agemax="69" agemin="65" name="Kategoria I" />
                <AGEGROUP agegroupid="5414" agemax="74" agemin="70" name="Kategoria J" />
                <AGEGROUP agegroupid="5415" agemax="79" agemin="75" name="Kategoria K" />
                <AGEGROUP agegroupid="5416" agemax="84" agemin="80" name="Kategoria L" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15641" daytime="11:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15642" daytime="11:42" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5417" daytime="11:44" gender="M" number="23" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9024" agemax="29" agemin="25" name="Kategoria A" />
                <AGEGROUP agegroupid="9025" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14816" />
                    <RANKING order="2" place="2" resultid="15477" />
                    <RANKING order="3" place="-1" resultid="14800" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9026" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14827" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9027" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14574" />
                    <RANKING order="2" place="2" resultid="15700" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9028" agemax="49" agemin="45" name="Kategoria E" />
                <AGEGROUP agegroupid="9029" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15046" />
                    <RANKING order="2" place="2" resultid="14710" />
                    <RANKING order="3" place="-1" resultid="15453" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9030" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15334" />
                    <RANKING order="2" place="2" resultid="14531" />
                    <RANKING order="3" place="3" resultid="15005" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9031" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14748" />
                    <RANKING order="2" place="2" resultid="15067" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9032" agemax="69" agemin="65" name="Kategoria I" />
                <AGEGROUP agegroupid="9033" agemax="74" agemin="70" name="Kategoria J" />
                <AGEGROUP agegroupid="9034" agemax="79" agemin="75" name="Kategoria K" />
                <AGEGROUP agegroupid="9035" agemax="84" agemin="80" name="Kategoria L" />
                <AGEGROUP agegroupid="9036" agemax="89" agemin="85" name="Kategoria M" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15643" daytime="11:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15644" daytime="11:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="15645" daytime="11:50" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1225" daytime="11:52" gender="F" number="24" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3209" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15040" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3210" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15767" />
                    <RANKING order="2" place="2" resultid="14731" />
                    <RANKING order="3" place="3" resultid="14755" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3211" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14804" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3212" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15468" />
                    <RANKING order="2" place="2" resultid="15244" />
                    <RANKING order="3" place="3" resultid="14665" />
                    <RANKING order="4" place="4" resultid="15692" />
                    <RANKING order="5" place="-1" resultid="15688" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3213" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14682" />
                    <RANKING order="2" place="2" resultid="15106" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3214" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14860" />
                    <RANKING order="2" place="2" resultid="15671" />
                    <RANKING order="3" place="3" resultid="14726" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3215" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15082" />
                    <RANKING order="2" place="2" resultid="15205" />
                    <RANKING order="3" place="3" resultid="15126" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3216" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15200" />
                    <RANKING order="2" place="2" resultid="15121" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3217" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14850" />
                    <RANKING order="2" place="2" resultid="14788" />
                    <RANKING order="3" place="3" resultid="14783" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3218" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15111" />
                    <RANKING order="2" place="2" resultid="14865" />
                    <RANKING order="3" place="3" resultid="15515" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3219" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14586" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3220" agemax="84" agemin="80" name="Kategoria L" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15646" daytime="11:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15647" daytime="11:54" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="15648" daytime="11:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="15649" daytime="12:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="15650" daytime="12:04" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1238" daytime="12:08" gender="M" number="25" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9037" agemax="29" agemin="25" name="Kategoria A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15318" />
                    <RANKING order="2" place="2" resultid="14660" />
                    <RANKING order="3" place="3" resultid="15229" />
                    <RANKING order="4" place="4" resultid="14518" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9038" agemax="34" agemin="30" name="Kategoria B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14817" />
                    <RANKING order="2" place="2" resultid="15478" />
                    <RANKING order="3" place="3" resultid="14798" />
                    <RANKING order="4" place="-1" resultid="14617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9039" agemax="39" agemin="35" name="Kategoria C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15224" />
                    <RANKING order="2" place="2" resultid="14687" />
                    <RANKING order="3" place="3" resultid="14537" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9040" agemax="44" agemin="40" name="Kategoria D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14575" />
                    <RANKING order="2" place="2" resultid="14704" />
                    <RANKING order="3" place="3" resultid="15772" />
                    <RANKING order="4" place="4" resultid="14525" />
                    <RANKING order="5" place="5" resultid="15717" />
                    <RANKING order="6" place="6" resultid="15181" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9041" agemax="49" agemin="45" name="Kategoria E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14612" />
                    <RANKING order="2" place="2" resultid="15239" />
                    <RANKING order="3" place="3" resultid="14807" />
                    <RANKING order="4" place="-1" resultid="14812" />
                    <RANKING order="5" place="-1" resultid="14821" />
                    <RANKING order="6" place="-1" resultid="15220" />
                    <RANKING order="7" place="-1" resultid="15324" />
                    <RANKING order="8" place="-1" resultid="15525" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9042" agemax="54" agemin="50" name="Kategoria F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15154" />
                    <RANKING order="2" place="2" resultid="15139" />
                    <RANKING order="3" place="3" resultid="14778" />
                    <RANKING order="4" place="4" resultid="15191" />
                    <RANKING order="5" place="5" resultid="15449" />
                    <RANKING order="6" place="-1" resultid="14711" />
                    <RANKING order="7" place="-1" resultid="15733" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9043" agemax="59" agemin="55" name="Kategoria G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15722" />
                    <RANKING order="2" place="2" resultid="15062" />
                    <RANKING order="3" place="3" resultid="15215" />
                    <RANKING order="4" place="4" resultid="15291" />
                    <RANKING order="5" place="5" resultid="15028" />
                    <RANKING order="6" place="6" resultid="15006" />
                    <RANKING order="7" place="7" resultid="15726" />
                    <RANKING order="8" place="8" resultid="14736" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9044" agemax="64" agemin="60" name="Kategoria H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15298" />
                    <RANKING order="2" place="2" resultid="15329" />
                    <RANKING order="3" place="3" resultid="14566" />
                    <RANKING order="4" place="4" resultid="15186" />
                    <RANKING order="5" place="5" resultid="14749" />
                    <RANKING order="6" place="6" resultid="14696" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9045" agemax="69" agemin="65" name="Kategoria I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15258" />
                    <RANKING order="2" place="2" resultid="14543" />
                    <RANKING order="3" place="3" resultid="14870" />
                    <RANKING order="4" place="4" resultid="15286" />
                    <RANKING order="5" place="5" resultid="15034" />
                    <RANKING order="6" place="6" resultid="14548" />
                    <RANKING order="7" place="7" resultid="15495" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9046" agemax="74" agemin="70" name="Kategoria J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14845" />
                    <RANKING order="2" place="2" resultid="14581" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9047" agemax="79" agemin="75" name="Kategoria K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14608" />
                    <RANKING order="2" place="2" resultid="14591" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9048" agemax="84" agemin="80" name="Kategoria L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14596" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9049" agemax="89" agemin="85" name="Kategoria M" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15651" daytime="12:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15652" daytime="12:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="15653" daytime="12:12" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="15654" daytime="12:14" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="15655" daytime="12:16" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="15656" daytime="12:18" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="15657" daytime="12:22" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="15658" daytime="12:24" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="15659" daytime="12:26" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="15660" daytime="12:28" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1290" daytime="12:32" gender="X" number="26" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="14501" agemax="-1" agemin="-1" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="15269" />
                    <RANKING order="2" place="2" resultid="14828" />
                    <RANKING order="3" place="3" resultid="15746" />
                    <RANKING order="4" place="4" resultid="15460" />
                    <RANKING order="5" place="5" resultid="15749" />
                    <RANKING order="6" place="6" resultid="15271" />
                    <RANKING order="7" place="7" resultid="15270" />
                    <RANKING order="8" place="8" resultid="14795" />
                    <RANKING order="9" place="9" resultid="15273" />
                    <RANKING order="10" place="10" resultid="15272" />
                    <RANKING order="11" place="11" resultid="15747" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="15661" daytime="12:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="15662" daytime="12:34" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="JWOR" nation="POL" clubid="14967" name="Ukp &quot;Na Fali&quot; Jawor">
          <ATHLETES>
            <ATHLETE firstname="Paweł" lastname="Jarecki" birthdate="1977-01-20" gender="M" nation="POL" athleteid="14976">
              <RESULTS>
                <RESULT eventid="1066" points="301" swimtime="00:03:40.17" resultid="14977" heatid="15555" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.00" />
                    <SPLIT distance="100" swimtime="00:01:45.65" />
                    <SPLIT distance="150" swimtime="00:02:45.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5390" points="249" swimtime="00:01:35.32" resultid="14978" heatid="15601" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Subocz" birthdate="1963-09-11" gender="M" nation="POL" athleteid="14979">
              <RESULTS>
                <RESULT comment="M-4" eventid="1144" status="DSQ" swimtime="00:00:00.00" resultid="14980" heatid="15583" lane="4" />
                <RESULT eventid="5390" points="181" swimtime="00:02:00.51" resultid="14981" heatid="15600" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Urbańska" birthdate="1980-07-06" gender="F" nation="POL" athleteid="14968">
              <RESULTS>
                <RESULT eventid="1157" points="195" swimtime="00:03:42.82" resultid="14969" heatid="15586" lane="5" />
                <RESULT eventid="1198" points="249" swimtime="00:02:00.26" resultid="14970" heatid="15623" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Florek" birthdate="1976-06-29" gender="M" nation="POL" athleteid="14971">
              <RESULTS>
                <RESULT eventid="1212" points="288" swimtime="00:01:39.94" resultid="14972" heatid="15629" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Wojdyło" birthdate="1973-04-12" gender="M" nation="POL" athleteid="14973">
              <RESULTS>
                <RESULT eventid="1170" points="299" swimtime="00:02:56.44" resultid="14974" heatid="15592" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                    <SPLIT distance="100" swimtime="00:01:21.78" />
                    <SPLIT distance="150" swimtime="00:02:08.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5390" points="274" swimtime="00:01:31.25" resultid="14975" heatid="15600" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LCGW" nation="POL" clubid="14829" name="Landsberg Crew Gorzów Wlkp.">
          <ATHLETES>
            <ATHLETE firstname="Stanislaw" lastname="Kaczmarek" birthdate="1979-01-26" gender="M" nation="POL" athleteid="15768">
              <RESULTS>
                <RESULT eventid="1066" points="621" swimtime="00:02:47.42" resultid="15769" heatid="15552" lane="5" entrytime="00:02:39.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.38" />
                    <SPLIT distance="100" swimtime="00:01:17.40" />
                    <SPLIT distance="150" swimtime="00:02:01.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="630" swimtime="00:02:11.84" resultid="15770" heatid="15588" lane="2" entrytime="00:02:07.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                    <SPLIT distance="100" swimtime="00:01:06.57" />
                    <SPLIT distance="150" swimtime="00:01:39.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="659" swimtime="00:01:13.06" resultid="15771" heatid="15624" lane="5" entrytime="00:01:11.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="653" swimtime="00:00:59.08" resultid="15772" heatid="15651" lane="2" entrytime="00:00:57.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Magdalena" lastname="Kaczmarek" birthdate="1992-08-23" gender="F" nation="POL" athleteid="15763">
              <RESULTS>
                <RESULT eventid="1157" points="776" swimtime="00:02:16.71" resultid="15764" heatid="15584" lane="4" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                    <SPLIT distance="100" swimtime="00:01:06.67" />
                    <SPLIT distance="150" swimtime="00:01:42.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5376" points="774" swimtime="00:01:10.60" resultid="15765" heatid="15593" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5430" points="727" swimtime="00:02:37.44" resultid="15766" heatid="15614" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                    <SPLIT distance="100" swimtime="00:01:14.51" />
                    <SPLIT distance="150" swimtime="00:01:55.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="815" swimtime="00:01:01.52" resultid="15767" heatid="15646" lane="4" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZRYBN" nation="POL" clubid="14513" name="NZ Rybnik">
          <ATHLETES>
            <ATHLETE firstname="Grzegorz" lastname="Kuczera" birthdate="1994-01-01" gender="M" nation="POL" swrid="4180253" athleteid="14514">
              <RESULTS>
                <RESULT eventid="1092" points="537" swimtime="00:00:28.10" resultid="14515" heatid="15562" lane="4" entrytime="00:00:27.90" />
                <RESULT eventid="5390" points="429" swimtime="00:01:13.16" resultid="14516" heatid="15598" lane="3" entrytime="00:01:13.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5443" points="262" swimtime="00:03:01.61" resultid="14517" heatid="15618" lane="3" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.41" />
                    <SPLIT distance="100" swimtime="00:01:28.68" />
                    <SPLIT distance="150" swimtime="00:02:15.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="437" swimtime="00:01:03.97" resultid="14518" heatid="15652" lane="6" entrytime="00:01:03.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02016" nation="POL" region="16" clubid="15029" name="Koszalińskie TKKF">
          <ATHLETES>
            <ATHLETE firstname="Marian" lastname="Lasowy" birthdate="1955-07-15" gender="M" nation="POL" license="502016700001" swrid="4967127" athleteid="15030">
              <RESULTS>
                <RESULT eventid="1092" points="338" swimtime="00:00:39.59" resultid="15031" heatid="15567" lane="4" entrytime="00:00:41.02" entrycourse="SCM" />
                <RESULT eventid="1170" points="334" swimtime="00:03:20.81" resultid="15032" heatid="15590" lane="5" entrytime="00:03:20.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.77" />
                    <SPLIT distance="100" swimtime="00:01:36.69" />
                    <SPLIT distance="150" swimtime="00:02:30.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="224" swimtime="00:00:54.80" resultid="15033" heatid="15638" lane="6" entrytime="00:00:51.57" entrycourse="SCM" />
                <RESULT eventid="1238" points="319" swimtime="00:01:29.42" resultid="15034" heatid="15657" lane="6" entrytime="00:01:31.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03415" nation="POL" clubid="14763" name="UKS Cityzen Poznan">
          <ATHLETES>
            <ATHLETE firstname="Małgorzata" lastname="Łasińska" birthdate="1954-07-13" gender="F" nation="POL" swrid="5471727" athleteid="14779">
              <RESULTS>
                <RESULT eventid="1131" points="196" swimtime="00:01:00.86" resultid="14780" heatid="15577" lane="4" entrytime="00:01:01.75" entrycourse="SCM" />
                <RESULT eventid="5376" points="248" swimtime="00:02:10.32" resultid="14781" heatid="15594" lane="1" entrytime="00:02:09.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="307" swimtime="00:00:59.31" resultid="14782" heatid="15633" lane="4" entrytime="00:00:58.85" entrycourse="SCM" />
                <RESULT eventid="1225" points="169" swimtime="00:02:08.34" resultid="14783" heatid="15648" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Matyszczak" birthdate="1970-12-14" gender="M" nation="POL" swrid="5471729" athleteid="14774">
              <RESULTS>
                <RESULT eventid="1092" points="522" swimtime="00:00:30.41" resultid="14775" heatid="15563" lane="6" entrytime="00:00:30.50" />
                <RESULT eventid="1170" points="370" swimtime="00:02:44.46" resultid="14776" heatid="15589" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.78" />
                    <SPLIT distance="100" swimtime="00:01:17.47" />
                    <SPLIT distance="150" swimtime="00:02:01.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="330" swimtime="00:00:41.02" resultid="14777" heatid="15636" lane="6" entrytime="00:00:40.00" />
                <RESULT eventid="1238" points="408" swimtime="00:01:11.53" resultid="14778" heatid="15654" lane="3" entrytime="00:01:10.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rusłana" lastname="Dembecka" birthdate="1957-10-01" gender="F" nation="POL" athleteid="14784">
              <RESULTS>
                <RESULT eventid="1053" points="380" swimtime="00:04:37.17" resultid="14785" heatid="15550" lane="5" entrytime="00:04:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.90" />
                    <SPLIT distance="100" swimtime="00:02:11.85" />
                    <SPLIT distance="150" swimtime="00:03:25.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="303" swimtime="00:00:57.87" resultid="14786" heatid="15603" lane="2" entrytime="00:00:56.00" />
                <RESULT eventid="1198" points="311" swimtime="00:02:10.46" resultid="14787" heatid="15622" lane="2" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="206" swimtime="00:02:00.10" resultid="14788" heatid="15648" lane="1" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Boryski" birthdate="1951-03-05" gender="M" nation="POL" swrid="4754708" athleteid="14764">
              <RESULTS>
                <RESULT eventid="1170" points="362" swimtime="00:03:27.62" resultid="14765" heatid="15590" lane="6" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.59" />
                    <SPLIT distance="100" swimtime="00:01:41.05" />
                    <SPLIT distance="150" swimtime="00:02:35.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5443" points="489" swimtime="00:03:50.88" resultid="14766" heatid="15618" lane="5" entrytime="00:03:50.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.36" />
                    <SPLIT distance="100" swimtime="00:01:53.62" />
                    <SPLIT distance="150" swimtime="00:02:53.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="402" swimtime="00:00:46.97" resultid="14767" heatid="15638" lane="4" entrytime="00:00:46.04" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Nochowicz" birthdate="1951-06-03" gender="M" nation="POL" swrid="5471731" athleteid="14768">
              <RESULTS>
                <RESULT eventid="1118" points="206" swimtime="00:02:06.98" resultid="14769" heatid="15574" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="187" swimtime="00:01:00.61" resultid="14770" heatid="15639" lane="5" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sławomir" lastname="Cybertowicz" birthdate="1966-01-12" gender="M" nation="POL" swrid="4269915" athleteid="14771">
              <RESULTS>
                <RESULT eventid="6830" points="442" swimtime="00:00:40.03" resultid="14772" heatid="15606" lane="5" entrytime="00:00:37.70" entrycourse="SCM" />
                <RESULT eventid="1316" points="280" swimtime="00:00:44.82" resultid="14773" heatid="15637" lane="1" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Putowska" birthdate="1962-01-22" gender="F" nation="POL" swrid="5416834" athleteid="14789">
              <RESULTS>
                <RESULT eventid="1053" points="402" swimtime="00:04:13.88" resultid="14790" heatid="15550" lane="3" entrytime="00:03:57.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.93" />
                    <SPLIT distance="100" swimtime="00:01:59.46" />
                    <SPLIT distance="150" swimtime="00:03:06.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5376" points="370" swimtime="00:01:50.09" resultid="14791" heatid="15594" lane="5" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5430" points="378" swimtime="00:04:01.11" resultid="14792" heatid="15615" lane="3" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.95" />
                    <SPLIT distance="100" swimtime="00:01:58.47" />
                    <SPLIT distance="150" swimtime="00:03:01.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="393" swimtime="00:01:56.22" resultid="14793" heatid="15621" lane="1" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="6828" swimtime="00:02:44.29" resultid="14794" heatid="15612" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                    <SPLIT distance="100" swimtime="00:01:23.79" />
                    <SPLIT distance="150" swimtime="00:02:13.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14789" number="1" />
                    <RELAYPOSITION athleteid="14764" number="2" />
                    <RELAYPOSITION athleteid="14779" number="3" />
                    <RELAYPOSITION athleteid="14774" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1290" swimtime="00:02:45.81" resultid="14795" heatid="15662" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.21" />
                    <SPLIT distance="100" swimtime="00:01:36.94" />
                    <SPLIT distance="150" swimtime="00:02:14.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14764" number="1" />
                    <RELAYPOSITION athleteid="14789" number="2" />
                    <RELAYPOSITION athleteid="14771" number="3" />
                    <RELAYPOSITION athleteid="14774" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="TMBAR" nation="POL" clubid="14998" name="Team Masters Barracuda">
          <ATHLETES>
            <ATHLETE firstname="Marek" lastname="Gola" birthdate="1981-04-18" gender="M" nation="POL" athleteid="14999">
              <RESULTS>
                <RESULT eventid="1144" points="143" swimtime="00:00:48.01" resultid="15000" heatid="15583" lane="2" />
                <RESULT eventid="5390" points="186" swimtime="00:01:44.78" resultid="15001" heatid="15600" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00211" nation="POL" region="11" clubid="15041" name="KS Górnik Radlin">
          <ATHLETES>
            <ATHLETE firstname="Ryszard" lastname="Kubica" birthdate="1972-02-22" gender="M" nation="POL" license="100211700343" swrid="5398297" athleteid="15042">
              <RESULTS>
                <RESULT eventid="1118" points="453" swimtime="00:01:18.73" resultid="15043" heatid="15572" lane="6" entrytime="00:01:17.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="477" swimtime="00:00:34.29" resultid="15044" heatid="15580" lane="2" entrytime="00:00:32.04" entrycourse="SCM" />
                <RESULT eventid="5443" points="512" swimtime="00:02:53.87" resultid="15045" heatid="15617" lane="1" entrytime="00:02:52.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.64" />
                    <SPLIT distance="100" swimtime="00:01:24.25" />
                    <SPLIT distance="150" swimtime="00:02:09.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5417" points="487" swimtime="00:01:15.80" resultid="15046" heatid="15644" lane="3" entrytime="00:01:13.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02706" nation="POL" region="06" clubid="15302" name="UKS ,,Jasień&apos;&apos; Sucha Beskidzka">
          <ATHLETES>
            <ATHLETE firstname="Aneta" lastname="Pytel" birthdate="1979-02-03" gender="F" nation="POL" license="102706600133" swrid="5582461" athleteid="15303">
              <RESULTS>
                <RESULT eventid="1053" points="280" swimtime="00:04:13.79" resultid="15304" heatid="15550" lane="2" entrytime="00:04:16.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.94" />
                    <SPLIT distance="100" swimtime="00:02:02.38" />
                    <SPLIT distance="150" swimtime="00:03:08.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="191" swimtime="00:00:50.82" resultid="15305" heatid="15578" lane="2" />
                <RESULT eventid="1198" points="266" swimtime="00:01:57.58" resultid="15306" heatid="15621" lane="6" entrytime="00:01:56.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="238" swimtime="00:00:49.25" resultid="15307" heatid="15632" lane="1" entrytime="00:00:48.30" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sabina" lastname="Sikora" birthdate="1984-10-03" gender="F" nation="POL" license="102706600159" swrid="5468086" athleteid="15308">
              <RESULTS>
                <RESULT eventid="1079" points="695" swimtime="00:00:29.55" resultid="15309" heatid="15557" lane="2" entrytime="00:00:29.28" entrycourse="SCM" />
                <RESULT eventid="1183" points="638" swimtime="00:00:36.77" resultid="15310" heatid="15602" lane="4" entrytime="00:00:35.13" entrycourse="SCM" />
                <RESULT eventid="1198" points="576" swimtime="00:01:22.98" resultid="15311" heatid="15620" lane="4" entrytime="00:01:22.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="614" swimtime="00:00:36.33" resultid="15312" heatid="15634" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZŚW" nation="POL" clubid="14532" name="NZ Środa Wielkopolska">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Grzelczak" birthdate="1985-01-01" gender="M" nation="POL" athleteid="14533">
              <RESULTS>
                <RESULT eventid="1066" points="290" swimtime="00:03:32.19" resultid="14534" heatid="15556" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.45" />
                    <SPLIT distance="100" swimtime="00:01:38.98" />
                    <SPLIT distance="150" swimtime="00:02:35.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6830" points="329" swimtime="00:00:41.77" resultid="14535" heatid="15609" lane="1" />
                <RESULT eventid="1212" points="323" swimtime="00:01:32.50" resultid="14536" heatid="15629" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="196" swimtime="00:01:24.97" resultid="14537" heatid="15660" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZJARO" nation="POL" clubid="14544" name="NZ Jarocin">
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Marszałek" birthdate="1954-01-01" gender="M" nation="POL" athleteid="14545">
              <RESULTS>
                <RESULT eventid="1144" points="213" swimtime="00:00:51.17" resultid="14546" heatid="15582" lane="4" entrytime="00:00:50.42" />
                <RESULT eventid="1170" points="287" swimtime="00:03:31.17" resultid="14547" heatid="15591" lane="3" entrytime="00:03:31.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.20" />
                    <SPLIT distance="100" swimtime="00:01:43.47" />
                    <SPLIT distance="150" swimtime="00:02:37.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="239" swimtime="00:01:38.43" resultid="14548" heatid="15658" lane="4" entrytime="00:01:33.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SLOWRO" nation="POL" clubid="15013" name="WKS Sląsk Wrocław">
          <ATHLETES>
            <ATHLETE firstname="Marek" lastname="Rother" birthdate="1968-05-21" gender="M" nation="POL" swrid="4351633" athleteid="15014">
              <RESULTS>
                <RESULT eventid="1118" points="779" swimtime="00:01:10.38" resultid="15015" heatid="15572" lane="2" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5390" points="809" swimtime="00:01:10.53" resultid="15016" heatid="15597" lane="6" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5443" points="860" swimtime="00:02:30.62" resultid="15017" heatid="15617" lane="4" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.83" />
                    <SPLIT distance="100" swimtime="00:01:14.59" />
                    <SPLIT distance="150" swimtime="00:01:53.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="837" swimtime="00:00:31.14" resultid="15018" heatid="15635" lane="5" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00201" nation="POL" region="01" clubid="15035" name="KS AZS AWF Wrocław">
          <ATHLETES>
            <ATHLETE firstname="Dominika" lastname="Sasin" birthdate="1994-05-29" gender="F" nation="POL" license="100201600097" swrid="4236079" athleteid="15036">
              <RESULTS>
                <RESULT eventid="1079" points="744" swimtime="00:00:27.91" resultid="15037" heatid="15557" lane="3" entrytime="00:00:27.16" entrycourse="SCM" />
                <RESULT eventid="1131" points="797" swimtime="00:00:29.75" resultid="15038" heatid="15575" lane="3" entrytime="00:00:28.78" entrycourse="SCM" />
                <RESULT eventid="5404" points="776" swimtime="00:01:06.36" resultid="15039" heatid="15641" lane="3" entrytime="00:01:04.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="793" swimtime="00:01:00.61" resultid="15040" heatid="15646" lane="3" entrytime="00:00:59.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LBL" nation="POL" clubid="14750" name="MASTERS Lublin">
          <ATHLETES>
            <ATHLETE firstname="Paulina" lastname="Kawecka" birthdate="1993-09-06" gender="F" nation="POL" swrid="5118335" athleteid="14751">
              <RESULTS>
                <RESULT eventid="1105" points="310" swimtime="00:01:35.00" resultid="14752" heatid="15570" lane="3" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5376" points="249" swimtime="00:01:42.95" resultid="14753" heatid="15594" lane="4" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5430" points="397" swimtime="00:03:12.63" resultid="14754" heatid="15614" lane="6" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.51" />
                    <SPLIT distance="100" swimtime="00:01:34.87" />
                    <SPLIT distance="150" swimtime="00:02:24.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="256" swimtime="00:01:30.46" resultid="14755" heatid="15648" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SQUAD" nation="POL" clubid="14712" name="Water Squad">
          <ATHLETES>
            <ATHLETE firstname="Karolina" lastname="Szyszkowska" birthdate="1996-11-05" gender="F" nation="POL" swrid="4282341" athleteid="14713">
              <RESULTS>
                <RESULT eventid="1053" points="870" swimtime="00:02:40.95" resultid="14714" heatid="15549" lane="3" entrytime="00:02:40.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.00" />
                    <SPLIT distance="100" swimtime="00:01:17.50" />
                    <SPLIT distance="150" swimtime="00:01:58.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="796" swimtime="00:00:34.08" resultid="14715" heatid="15602" lane="3" entrytime="00:00:34.52" entrycourse="SCM" />
                <RESULT eventid="1198" points="836" swimtime="00:01:14.98" resultid="14716" heatid="15620" lane="3" entrytime="00:01:14.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aneta" lastname="Dolińska" birthdate="1990-07-06" gender="F" nation="POL" swrid="4251116" athleteid="14727">
              <RESULTS>
                <RESULT eventid="1105" points="374" swimtime="00:01:29.25" resultid="14728" heatid="15569" lane="6" entrytime="00:01:29.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="490" swimtime="00:02:39.39" resultid="14729" heatid="15585" lane="3" entrytime="00:02:41.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                    <SPLIT distance="100" swimtime="00:01:15.59" />
                    <SPLIT distance="150" swimtime="00:01:57.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="421" swimtime="00:00:39.79" resultid="14730" heatid="15631" lane="6" entrytime="00:00:40.00" />
                <RESULT eventid="1225" points="527" swimtime="00:01:11.13" resultid="14731" heatid="15646" lane="6" entrytime="00:01:12.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Piaściński" birthdate="1976-09-19" gender="M" nation="POL" athleteid="15521">
              <RESULTS>
                <RESULT eventid="1092" points="614" swimtime="00:00:28.08" resultid="15522" heatid="15562" lane="2" entrytime="00:00:28.00" />
                <RESULT eventid="5390" points="616" swimtime="00:01:10.49" resultid="15523" heatid="15597" lane="5" entrytime="00:01:11.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5443" points="656" swimtime="00:02:31.43" resultid="15524" heatid="15617" lane="2" entrytime="00:02:39.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="100" swimtime="00:01:13.45" />
                    <SPLIT distance="150" swimtime="00:01:52.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" status="DNS" swimtime="00:00:00.00" resultid="15525" heatid="15653" lane="3" entrytime="00:01:04.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Matyszewski" birthdate="1971-10-11" gender="M" nation="POL" swrid="5582459" athleteid="14737">
              <RESULTS>
                <RESULT eventid="1066" points="466" swimtime="00:03:19.57" resultid="14738" heatid="15553" lane="2" entrytime="00:03:21.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.69" />
                    <SPLIT distance="100" swimtime="00:01:33.15" />
                    <SPLIT distance="150" swimtime="00:02:25.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6830" points="453" swimtime="00:00:40.05" resultid="14739" heatid="15606" lane="6" entrytime="00:00:38.92" entrycourse="SCM" />
                <RESULT eventid="1212" points="431" swimtime="00:01:28.84" resultid="14740" heatid="15626" lane="3" entrytime="00:01:30.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="292" swimtime="00:00:42.73" resultid="14741" heatid="15638" lane="3" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Adamowicz" birthdate="1967-07-11" gender="M" nation="POL" swrid="4655152" athleteid="14732">
              <RESULTS>
                <RESULT eventid="1092" points="323" swimtime="00:00:37.92" resultid="14733" heatid="15566" lane="5" entrytime="00:00:37.03" entrycourse="SCM" />
                <RESULT eventid="6830" points="343" swimtime="00:00:43.57" resultid="14734" heatid="15607" lane="1" entrytime="00:00:42.48" entrycourse="SCM" />
                <RESULT eventid="1212" points="321" swimtime="00:01:39.45" resultid="14735" heatid="15627" lane="3" entrytime="00:01:38.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="260" swimtime="00:01:30.82" resultid="14736" heatid="15657" lane="5" entrytime="00:01:28.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Timea" lastname="Balajcza" birthdate="1971-09-22" gender="F" nation="POL" swrid="5240601" athleteid="14722">
              <RESULTS>
                <RESULT eventid="1053" points="692" swimtime="00:03:10.14" resultid="14723" heatid="15549" lane="4" entrytime="00:03:04.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.05" />
                    <SPLIT distance="100" swimtime="00:01:31.38" />
                    <SPLIT distance="150" swimtime="00:02:20.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="773" swimtime="00:00:39.01" resultid="14724" heatid="15602" lane="2" entrytime="00:00:38.05" entrycourse="SCM" />
                <RESULT eventid="1198" points="684" swimtime="00:01:27.49" resultid="14725" heatid="15620" lane="2" entrytime="00:01:27.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="521" swimtime="00:01:15.73" resultid="14726" heatid="15647" lane="2" entrytime="00:01:18.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="6828" swimtime="00:02:18.00" resultid="14744" heatid="15611" lane="2" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                    <SPLIT distance="100" swimtime="00:01:12.57" />
                    <SPLIT distance="150" swimtime="00:01:45.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15521" number="1" />
                    <RELAYPOSITION athleteid="14737" number="2" />
                    <RELAYPOSITION athleteid="14722" number="3" />
                    <RELAYPOSITION athleteid="14727" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1290" swimtime="00:02:13.31" resultid="14828" heatid="15661" lane="3" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                    <SPLIT distance="100" swimtime="00:01:11.20" />
                    <SPLIT distance="150" swimtime="00:01:41.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15521" number="1" />
                    <RELAYPOSITION athleteid="14737" number="2" />
                    <RELAYPOSITION athleteid="14713" number="3" />
                    <RELAYPOSITION athleteid="14727" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="ZABRZ" nation="POL" clubid="14840" name="Weteran  Zabrze">
          <ATHLETES>
            <ATHLETE firstname="Joanna" lastname="Zagała" birthdate="1959-06-24" gender="F" nation="POL" swrid="4934034" athleteid="14874">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="14875" heatid="15558" lane="6" entrytime="00:00:39.07" entrycourse="SCM" />
                <RESULT eventid="1157" status="DNS" swimtime="00:00:00.00" resultid="14876" heatid="15586" lane="4" />
                <RESULT eventid="5430" status="DNS" swimtime="00:00:00.00" resultid="14877" heatid="15616" lane="3" />
                <RESULT eventid="1303" status="DNS" swimtime="00:00:00.00" resultid="14878" heatid="15634" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Twardysko" birthdate="1956-01-16" gender="M" nation="POL" swrid="5464152" athleteid="14866">
              <RESULTS>
                <RESULT eventid="1092" points="434" swimtime="00:00:36.42" resultid="14867" heatid="15566" lane="4" entrytime="00:00:35.10" entrycourse="SCM" />
                <RESULT eventid="1170" points="476" swimtime="00:02:58.50" resultid="14868" heatid="15589" lane="6" entrytime="00:02:55.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.09" />
                    <SPLIT distance="100" swimtime="00:01:21.64" />
                    <SPLIT distance="150" swimtime="00:02:09.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5443" points="391" swimtime="00:03:35.42" resultid="14869" heatid="15618" lane="4" entrytime="00:03:33.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.76" />
                    <SPLIT distance="100" swimtime="00:01:41.90" />
                    <SPLIT distance="150" swimtime="00:02:38.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="463" swimtime="00:01:18.98" resultid="14870" heatid="15655" lane="1" entrytime="00:01:17.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Teresa" lastname="Żylińska" birthdate="1950-10-13" gender="F" nation="POL" swrid="5464154" athleteid="14861">
              <RESULTS>
                <RESULT eventid="1105" points="251" swimtime="00:02:21.19" resultid="14862" heatid="15570" lane="5" entrytime="00:02:15.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="222" swimtime="00:04:36.94" resultid="14863" heatid="15586" lane="3" entrytime="00:04:30.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:12.21" />
                    <SPLIT distance="150" swimtime="00:03:26.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5430" points="274" swimtime="00:05:04.56" resultid="14864" heatid="15615" lane="2" entrytime="00:05:07.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.16" />
                    <SPLIT distance="100" swimtime="00:02:29.49" />
                    <SPLIT distance="150" swimtime="00:03:49.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="199" swimtime="00:02:07.81" resultid="14865" heatid="15649" lane="4" entrytime="00:02:03.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zofia" lastname="Dąbrowska" birthdate="1958-02-05" gender="F" nation="POL" swrid="4934035" athleteid="14846">
              <RESULTS>
                <RESULT eventid="1079" points="397" swimtime="00:00:43.88" resultid="14847" heatid="15559" lane="3" entrytime="00:00:48.00" />
                <RESULT eventid="1131" points="197" swimtime="00:01:00.78" resultid="14848" heatid="15577" lane="3" entrytime="00:00:58.00" />
                <RESULT eventid="1198" points="310" swimtime="00:02:10.67" resultid="14849" heatid="15622" lane="4" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="274" swimtime="00:01:49.14" resultid="14850" heatid="15649" lane="3" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beata" lastname="Sulewska" birthdate="1972-11-02" gender="F" nation="POL" swrid="4792005" athleteid="14856">
              <RESULTS>
                <RESULT eventid="1079" points="689" swimtime="00:00:32.02" resultid="14857" heatid="15560" lane="4" />
                <RESULT eventid="1157" points="747" swimtime="00:02:27.61" resultid="14858" heatid="15584" lane="5" entrytime="00:02:26.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                    <SPLIT distance="100" swimtime="00:01:11.74" />
                    <SPLIT distance="150" swimtime="00:01:49.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="774" swimtime="00:01:23.95" resultid="14859" heatid="15620" lane="5" entrytime="00:01:27.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="661" swimtime="00:01:09.95" resultid="14860" heatid="15646" lane="5" entrytime="00:01:09.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Kosiak" birthdate="1940-04-20" gender="M" nation="POL" athleteid="14871">
              <RESULTS>
                <RESULT eventid="1092" points="333" swimtime="00:00:46.26" resultid="14872" heatid="15567" lane="5" entrytime="00:00:49.00" />
                <RESULT eventid="1144" points="160" swimtime="00:01:06.47" resultid="14873" heatid="15582" lane="2" entrytime="00:01:07.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiesław" lastname="Kornicki" birthdate="1949-01-28" gender="M" nation="POL" swrid="4137183" athleteid="14841">
              <RESULTS>
                <RESULT eventid="1092" points="586" swimtime="00:00:33.92" resultid="14842" heatid="15564" lane="5" entrytime="00:00:32.59" entrycourse="SCM" />
                <RESULT eventid="1144" points="514" swimtime="00:00:39.97" resultid="14843" heatid="15581" lane="2" entrytime="00:00:38.00" entrycourse="SCM" />
                <RESULT eventid="1316" points="348" swimtime="00:00:49.28" resultid="14844" heatid="15638" lane="1" entrytime="00:00:48.00" />
                <RESULT eventid="1238" points="502" swimtime="00:01:21.30" resultid="14845" heatid="15656" lane="6" entrytime="00:01:20.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Genowefa" lastname="Dru.Zyńska" birthdate="1951-02-18" gender="F" nation="POL" athleteid="14851">
              <RESULTS>
                <RESULT eventid="1053" points="234" swimtime="00:05:45.82" resultid="14852" heatid="15551" lane="2" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.24" />
                    <SPLIT distance="100" swimtime="00:02:47.41" />
                    <SPLIT distance="150" swimtime="00:04:17.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="264" swimtime="00:01:07.23" resultid="14853" heatid="15603" lane="5" entrytime="00:01:05.00" />
                <RESULT eventid="1198" points="210" swimtime="00:02:43.23" resultid="14854" heatid="15622" lane="1" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="263" swimtime="00:01:05.23" resultid="14855" heatid="15633" lane="1" entrytime="00:01:20.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03315" nation="POL" region="15" clubid="15127" name="KU AZS UAM Poznań">
          <ATHLETES>
            <ATHLETE firstname="Tomasz" lastname="Juszkiewicz" birthdate="1974-05-10" gender="M" nation="POL" license="503315700077" swrid="5537971" athleteid="15131">
              <RESULTS>
                <RESULT eventid="1092" points="458" swimtime="00:00:30.96" resultid="15132" heatid="15564" lane="4" entrytime="00:00:30.97" entrycourse="SCM" />
                <RESULT eventid="5390" points="275" swimtime="00:01:32.21" resultid="15133" heatid="15600" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Kaczmarek" birthdate="1982-10-03" gender="M" nation="POL" license="503315700221" swrid="5471723" athleteid="15128">
              <RESULTS>
                <RESULT eventid="1092" points="554" swimtime="00:00:28.25" resultid="15129" heatid="15568" lane="4" />
                <RESULT eventid="1170" points="459" swimtime="00:02:26.47" resultid="15130" heatid="15591" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                    <SPLIT distance="100" swimtime="00:01:09.53" />
                    <SPLIT distance="150" swimtime="00:01:48.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01713" nation="POL" region="13" clubid="15019" />
        <CLUB type="CLUB" code="ASTBYD" nation="POL" clubid="14508" name="MKS ASTORIA Bydgoszcz">
          <ATHLETES>
            <ATHLETE firstname="Dariusz" lastname="Kostkowski" birthdate="1970-01-01" gender="M" nation="POL" swrid="5471726" athleteid="14509">
              <RESULTS>
                <RESULT eventid="1118" points="148" swimtime="00:01:54.25" resultid="14510" heatid="15573" lane="6" entrytime="00:01:55.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5443" points="162" swimtime="00:04:15.22" resultid="14511" heatid="15619" lane="3" entrytime="00:04:21.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.46" />
                    <SPLIT distance="100" swimtime="00:02:05.31" />
                    <SPLIT distance="150" swimtime="00:03:10.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="180" swimtime="00:00:50.21" resultid="14512" heatid="15639" lane="3" entrytime="00:00:53.09" entrycourse="SCM" />
                <RESULT eventid="6830" points="282" swimtime="00:00:46.86" resultid="14519" heatid="15608" lane="1" entrytime="00:00:48.74" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="EXOBO" nation="POL" clubid="14603" name="Ks Extreme Team Oborniki">
          <ATHLETES>
            <ATHLETE firstname="Janusz" lastname="Wolniewicz" birthdate="1948-12-22" gender="M" nation="POL" swrid="4754624" athleteid="14604">
              <RESULTS>
                <RESULT eventid="1092" points="516" swimtime="00:00:39.01" resultid="14605" heatid="15567" lane="3" entrytime="00:00:39.14" />
                <RESULT eventid="1170" points="319" swimtime="00:03:52.65" resultid="14606" heatid="15590" lane="2" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.59" />
                    <SPLIT distance="100" swimtime="00:01:42.98" />
                    <SPLIT distance="150" swimtime="00:02:46.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="259" swimtime="00:00:57.10" resultid="14607" heatid="15639" lane="2" entrytime="00:00:58.00" />
                <RESULT eventid="1238" points="405" swimtime="00:01:36.16" resultid="14608" heatid="15657" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04901" nation="POL" region="01" clubid="15094" name="KS Neptun Świdnica">
          <ATHLETES>
            <ATHLETE firstname="Bartłomiej" lastname="Żukowski" birthdate="1993-04-26" gender="M" nation="POL" license="104901700097" swrid="4087259" athleteid="15095">
              <RESULTS>
                <RESULT eventid="1092" points="782" swimtime="00:00:24.02" resultid="15096" heatid="15561" lane="3" entrytime="00:00:23.79" entrycourse="SCM" />
                <RESULT eventid="6830" points="834" swimtime="00:00:29.54" resultid="15097" heatid="15605" lane="3" entrytime="00:00:28.90" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="06306" nation="POL" region="06" clubid="15047" name="Ks Korona 1919">
          <ATHLETES>
            <ATHLETE firstname="Mariola" lastname="Kuliś" birthdate="1966-07-27" gender="F" nation="POL" license="506306600043" swrid="4992797" athleteid="15078">
              <RESULTS>
                <RESULT eventid="1131" points="833" swimtime="00:00:33.95" resultid="15079" heatid="15575" lane="5" entrytime="00:00:33.98" entrycourse="SCM" />
                <RESULT eventid="1183" points="964" swimtime="00:00:38.02" resultid="15080" heatid="15602" lane="5" entrytime="00:00:38.57" entrycourse="SCM" />
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="15081" heatid="15620" lane="1" entrytime="00:01:29.58" entrycourse="SCM" />
                <RESULT eventid="1225" points="658" swimtime="00:01:12.11" resultid="15082" heatid="15650" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adam" lastname="Pycia" birthdate="1966-02-21" gender="M" nation="POL" license="506306700057" swrid="4992712" athleteid="15058">
              <RESULTS>
                <RESULT eventid="1066" points="502" swimtime="00:03:23.74" resultid="15059" heatid="15554" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.69" />
                    <SPLIT distance="100" swimtime="00:01:36.65" />
                    <SPLIT distance="150" swimtime="00:02:29.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6830" points="411" swimtime="00:00:41.00" resultid="15060" heatid="15607" lane="2" entrytime="00:00:40.87" entrycourse="SCM" />
                <RESULT eventid="1212" points="414" swimtime="00:01:31.36" resultid="15061" heatid="15625" lane="6" entrytime="00:01:30.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="580" swimtime="00:01:09.56" resultid="15062" heatid="15653" lane="1" entrytime="00:01:08.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Leńczowska" birthdate="1982-01-15" gender="F" nation="POL" license="506306600071" swrid="4992907" athleteid="15068">
              <RESULTS>
                <RESULT eventid="1105" points="610" swimtime="00:01:20.13" resultid="15069" heatid="15569" lane="5" entrytime="00:01:21.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5376" points="582" swimtime="00:01:21.58" resultid="15070" heatid="15595" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5430" points="607" swimtime="00:02:56.44" resultid="15071" heatid="15616" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.91" />
                    <SPLIT distance="100" swimtime="00:01:26.45" />
                    <SPLIT distance="150" swimtime="00:02:12.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="568" swimtime="00:00:36.88" resultid="15072" heatid="15631" lane="2" entrytime="00:00:36.33" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Macierzewska" birthdate="1960-04-20" gender="F" nation="POL" license="506306600048" swrid="4992827" athleteid="15083">
              <RESULTS>
                <RESULT eventid="1157" points="573" swimtime="00:02:56.63" resultid="15084" heatid="15586" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.07" />
                    <SPLIT distance="100" swimtime="00:01:25.56" />
                    <SPLIT distance="150" swimtime="00:02:12.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5376" points="632" swimtime="00:01:32.16" resultid="15085" heatid="15595" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="630" swimtime="00:00:42.35" resultid="15086" heatid="15632" lane="2" entrytime="00:00:42.48" entrycourse="SCM" />
                <RESULT eventid="5404" points="678" swimtime="00:01:32.70" resultid="15087" heatid="15642" lane="3" entrytime="00:01:31.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Łysiak" birthdate="1973-03-30" gender="M" nation="POL" license="506306700047" swrid="5468085" athleteid="15053">
              <RESULTS>
                <RESULT eventid="1066" status="DNS" swimtime="00:00:00.00" resultid="15054" heatid="15555" lane="5" />
                <RESULT eventid="1144" points="424" swimtime="00:00:35.66" resultid="15055" heatid="15582" lane="5" />
                <RESULT eventid="1212" points="460" swimtime="00:01:26.93" resultid="15056" heatid="15625" lane="4" entrytime="00:01:23.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="401" swimtime="00:00:38.44" resultid="15057" heatid="15639" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulina" lastname="Bielańska" birthdate="1984-04-20" gender="F" nation="POL" license="506306600072" swrid="5468078" athleteid="15048">
              <RESULTS>
                <RESULT eventid="1053" points="178" swimtime="00:04:35.43" resultid="15049" heatid="15551" lane="3" entrytime="00:04:54.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.34" />
                    <SPLIT distance="100" swimtime="00:02:16.18" />
                    <SPLIT distance="150" swimtime="00:03:26.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1079" points="153" swimtime="00:00:48.87" resultid="15050" heatid="15559" lane="4" entrytime="00:00:51.47" entrycourse="LCM" />
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="15051" heatid="15623" lane="2" />
                <RESULT eventid="1303" points="189" swimtime="00:00:53.78" resultid="15052" heatid="15633" lane="3" entrytime="00:00:53.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Janusz" lastname="Toporski" birthdate="1959-10-20" gender="M" nation="POL" license="506306700060" swrid="5484421" athleteid="15063">
              <RESULTS>
                <RESULT eventid="1066" points="447" swimtime="00:03:36.91" resultid="15064" heatid="15555" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.29" />
                    <SPLIT distance="100" swimtime="00:01:46.66" />
                    <SPLIT distance="150" swimtime="00:02:42.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5390" points="274" swimtime="00:01:45.09" resultid="15065" heatid="15601" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="361" swimtime="00:01:43.68" resultid="15066" heatid="15627" lane="6" entrytime="00:01:41.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5417" points="197" swimtime="00:01:55.70" resultid="15067" heatid="15644" lane="5" entrytime="00:01:51.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Janeczko" birthdate="1972-12-23" gender="F" nation="POL" license="506306600033" swrid="4218717" athleteid="15073">
              <RESULTS>
                <RESULT eventid="1131" points="605" swimtime="00:00:36.82" resultid="15074" heatid="15578" lane="3" />
                <RESULT eventid="5376" points="383" swimtime="00:01:35.06" resultid="15075" heatid="15595" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5430" points="390" swimtime="00:03:20.90" resultid="15076" heatid="15616" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.64" />
                    <SPLIT distance="100" swimtime="00:01:39.56" />
                    <SPLIT distance="150" swimtime="00:02:32.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5404" points="382" swimtime="00:01:33.16" resultid="15077" heatid="15642" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="6828" swimtime="00:02:05.51" resultid="15088" heatid="15611" lane="4" entrytime="00:02:04.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.80" />
                    <SPLIT distance="100" swimtime="00:01:02.68" />
                    <SPLIT distance="150" swimtime="00:01:34.63" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15058" number="1" />
                    <RELAYPOSITION athleteid="15078" number="2" />
                    <RELAYPOSITION athleteid="15068" number="3" />
                    <RELAYPOSITION athleteid="15053" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="NZWROC" nation="POL" region="01" clubid="14520" name="NZ Wrocław">
          <ATHLETES>
            <ATHLETE firstname="Małgorzata" lastname="Bołtuć" birthdate="1983-06-13" gender="F" nation="POL" athleteid="14983">
              <RESULTS>
                <RESULT eventid="1157" points="477" swimtime="00:02:45.48" resultid="14984" heatid="15585" lane="4" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.79" />
                    <SPLIT distance="100" swimtime="00:01:20.05" />
                    <SPLIT distance="150" swimtime="00:02:02.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5376" points="398" swimtime="00:01:32.61" resultid="14985" heatid="15593" lane="5" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5430" points="444" swimtime="00:03:15.74" resultid="14986" heatid="15614" lane="5" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.77" />
                    <SPLIT distance="100" swimtime="00:01:36.09" />
                    <SPLIT distance="150" swimtime="00:02:26.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="352" swimtime="00:01:47.13" resultid="14987" heatid="15621" lane="2" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" lastname="Wciórka" birthdate="1982-01-01" gender="M" nation="POL" athleteid="14521">
              <RESULTS>
                <RESULT eventid="1092" points="591" swimtime="00:00:27.65" resultid="14522" heatid="15563" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="6830" points="572" swimtime="00:00:35.02" resultid="14523" heatid="15606" lane="3" entrytime="00:00:36.00" />
                <RESULT eventid="1212" points="475" swimtime="00:01:21.49" resultid="14524" heatid="15625" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="527" swimtime="00:01:03.46" resultid="14525" heatid="15653" lane="4" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alina" lastname="Piekarska" birthdate="1947-07-15" gender="F" nation="POL" athleteid="14555">
              <RESULTS>
                <RESULT eventid="1183" points="39" swimtime="00:02:18.70" resultid="14556" heatid="15604" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="POZNAŃ" nation="POL" clubid="15444" name="NZ Poznań">
          <ATHLETES>
            <ATHLETE firstname="Mateusz" lastname="Kędzior" birthdate="1973-11-08" gender="M" nation="POL" athleteid="15445">
              <RESULTS>
                <RESULT eventid="1170" points="362" swimtime="00:02:45.72" resultid="15446" heatid="15589" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.12" />
                    <SPLIT distance="100" swimtime="00:01:20.96" />
                    <SPLIT distance="150" swimtime="00:02:03.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5390" points="286" swimtime="00:01:30.03" resultid="15447" heatid="15599" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5443" points="321" swimtime="00:03:23.22" resultid="15448" heatid="15617" lane="6" entrytime="00:03:15.00" />
                <RESULT eventid="1238" points="376" swimtime="00:01:13.54" resultid="15449" heatid="15654" lane="5" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="FOKA" nation="POL" clubid="14570" name="Foka Masters TEAM">
          <ATHLETES>
            <ATHLETE firstname="Krzysztof" lastname="Kęsik" birthdate="1979-09-21" gender="M" nation="POL" athleteid="14571">
              <RESULTS>
                <RESULT eventid="5390" points="768" swimtime="00:01:05.30" resultid="14572" heatid="15596" lane="2" entrytime="00:01:04.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="693" swimtime="00:00:28.39" resultid="14573" heatid="15579" lane="4" entrytime="00:00:27.84" />
                <RESULT eventid="5417" points="722" swimtime="00:01:03.11" resultid="14574" heatid="15643" lane="2" entrytime="00:01:03.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="681" swimtime="00:00:58.27" resultid="14575" heatid="15651" lane="1" entrytime="00:00:58.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZBIEL" nation="POL" region="01" clubid="14988" name="NZ Bielawa">
          <ATHLETES>
            <ATHLETE firstname="Patryk" lastname="Źródlak" birthdate="1997-10-31" gender="M" nation="POL" athleteid="14989">
              <RESULTS>
                <RESULT eventid="1118" points="233" swimtime="00:01:29.39" resultid="14990" heatid="15574" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6830" points="313" swimtime="00:00:41.58" resultid="14991" heatid="15610" lane="4" />
                <RESULT eventid="1316" points="315" swimtime="00:00:36.78" resultid="14992" heatid="15640" lane="3" />
                <RESULT eventid="1212" points="312" swimtime="00:01:31.36" resultid="14993" heatid="15628" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAPOL" nation="POL" clubid="14618" name="KS Masters Polkowice">
          <ATHLETES>
            <ATHLETE firstname="Emilia" lastname="Kawula" birthdate="1941-10-02" gender="F" nation="POL" athleteid="15484">
              <RESULTS>
                <RESULT eventid="1079" points="84" swimtime="00:01:36.22" resultid="15485" heatid="15559" lane="1" />
                <RESULT eventid="1183" points="47" swimtime="00:02:16.44" resultid="15486" heatid="15604" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kazimierz" lastname="Rosik" birthdate="1955-11-11" gender="M" nation="POL" athleteid="15491">
              <RESULTS>
                <RESULT eventid="1092" points="274" swimtime="00:00:42.45" resultid="15492" heatid="15567" lane="2" entrytime="00:00:42.90" entrycourse="SCM" />
                <RESULT eventid="6830" points="281" swimtime="00:00:51.53" resultid="15493" heatid="15608" lane="6" entrytime="00:00:50.40" entrycourse="SCM" />
                <RESULT eventid="1212" points="298" swimtime="00:01:55.11" resultid="15494" heatid="15630" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="220" swimtime="00:01:41.17" resultid="15495" heatid="15659" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pavlo" lastname="Vechirko" birthdate="1968-01-02" gender="M" nation="POL" athleteid="15496">
              <RESULTS>
                <RESULT eventid="1118" points="562" swimtime="00:01:18.43" resultid="15497" heatid="15572" lane="1" entrytime="00:01:16.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6830" points="487" swimtime="00:00:38.76" resultid="15498" heatid="15606" lane="4" entrytime="00:00:37.00" entrycourse="SCM" />
                <RESULT eventid="1212" points="508" swimtime="00:01:25.36" resultid="15499" heatid="15625" lane="2" entrytime="00:01:24.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="498" swimtime="00:00:37.02" resultid="15500" heatid="15635" lane="6" entrytime="00:00:35.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Janina" lastname="Zając" birthdate="1946-08-16" gender="F" nation="POL" athleteid="15501">
              <RESULTS>
                <RESULT eventid="1079" points="109" swimtime="00:01:12.21" resultid="15502" heatid="15559" lane="5" entrytime="00:01:11.00" entrycourse="SCM" />
                <RESULT eventid="1105" points="136" swimtime="00:03:02.08" resultid="15503" heatid="15571" lane="3" entrytime="00:02:56.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:31.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5430" points="167" swimtime="00:06:07.83" resultid="15504" heatid="15615" lane="5" entrytime="00:06:10.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:29.11" />
                    <SPLIT distance="100" swimtime="00:02:58.49" />
                    <SPLIT distance="150" swimtime="00:04:35.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="102" swimtime="00:01:33.19" resultid="15505" heatid="15633" lane="6" entrytime="00:01:24.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Józefa" lastname="Wołoszczuk" birthdate="1953-01-23" gender="F" nation="POL" athleteid="15511">
              <RESULTS>
                <RESULT eventid="1079" points="140" swimtime="00:01:04.18" resultid="15512" heatid="15559" lane="2" entrytime="00:01:06.00" entrycourse="SCM" />
                <RESULT eventid="5376" points="105" swimtime="00:02:56.36" resultid="15513" heatid="15594" lane="6" entrytime="00:02:58.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="195" swimtime="00:01:12.01" resultid="15514" heatid="15633" lane="5" entrytime="00:01:11.00" entrycourse="SCM" />
                <RESULT eventid="1225" points="133" swimtime="00:02:26.03" resultid="15515" heatid="15649" lane="2" entrytime="00:02:18.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gizela" lastname="Wójcik" birthdate="1949-11-16" gender="F" nation="POL" athleteid="15506">
              <RESULTS>
                <RESULT eventid="1053" points="250" swimtime="00:05:38.08" resultid="15507" heatid="15551" lane="4" entrytime="00:05:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.38" />
                    <SPLIT distance="100" swimtime="00:02:39.69" />
                    <SPLIT distance="150" swimtime="00:04:07.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="199" swimtime="00:01:13.90" resultid="15508" heatid="15603" lane="1" entrytime="00:01:12.00" entrycourse="SCM" />
                <RESULT eventid="1198" points="222" swimtime="00:02:40.18" resultid="15509" heatid="15622" lane="6" entrytime="00:02:39.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="207" swimtime="00:01:10.60" resultid="15510" heatid="15633" lane="2" entrytime="00:01:09.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zdzisława" lastname="Pachom" birthdate="1945-10-10" gender="F" nation="POL" athleteid="15487">
              <RESULTS>
                <RESULT eventid="1079" points="56" swimtime="00:01:29.96" resultid="15488" heatid="15560" lane="3" />
                <RESULT eventid="1183" points="64" swimtime="00:01:57.63" resultid="15489" heatid="15604" lane="4" />
                <RESULT eventid="1303" points="74" swimtime="00:01:43.74" resultid="15490" heatid="15634" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bogdan" lastname="Jawor" birthdate="1947-04-23" gender="M" nation="POL" athleteid="15479">
              <RESULTS>
                <RESULT eventid="1118" points="273" swimtime="00:02:05.79" resultid="15480" heatid="15574" lane="2" entrytime="00:02:14.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5390" points="262" swimtime="00:02:10.44" resultid="15481" heatid="15600" lane="3" entrytime="00:02:07.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5443" points="273" swimtime="00:04:37.60" resultid="15482" heatid="15619" lane="4" entrytime="00:04:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.45" />
                    <SPLIT distance="100" swimtime="00:02:14.13" />
                    <SPLIT distance="150" swimtime="00:03:26.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="249" swimtime="00:00:57.84" resultid="15483" heatid="15639" lane="1" entrytime="00:01:01.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00115" nation="POL" region="15" clubid="15098" name="KS Warta Poznań">
          <ATHLETES>
            <ATHLETE firstname="Przemysław" lastname="Waraczewski" birthdate="1962-04-19" gender="M" nation="POL" license="100115700344" swrid="4992781" athleteid="15112">
              <RESULTS>
                <RESULT eventid="1066" points="652" swimtime="00:03:11.33" resultid="15113" heatid="15553" lane="4" entrytime="00:03:08.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.42" />
                    <SPLIT distance="100" swimtime="00:01:30.53" />
                    <SPLIT distance="150" swimtime="00:02:21.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6830" points="592" swimtime="00:00:38.99" resultid="15114" heatid="15606" lane="1" entrytime="00:00:38.55" entrycourse="SCM" />
                <RESULT eventid="1212" points="627" swimtime="00:01:26.29" resultid="15115" heatid="15625" lane="1" entrytime="00:01:26.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="446" swimtime="00:00:41.10" resultid="15116" heatid="15640" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Krupińska" birthdate="1953-05-24" gender="F" nation="POL" license="500115600520" swrid="4992790" athleteid="15107">
              <RESULTS>
                <RESULT eventid="1053" points="540" swimtime="00:04:21.81" resultid="15108" heatid="15550" lane="4" entrytime="00:04:11.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.92" />
                    <SPLIT distance="100" swimtime="00:02:06.32" />
                    <SPLIT distance="150" swimtime="00:03:14.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="493" swimtime="00:00:54.66" resultid="15109" heatid="15603" lane="3" entrytime="00:00:51.00" entrycourse="SCM" />
                <RESULT eventid="1198" points="504" swimtime="00:02:01.97" resultid="15110" heatid="15622" lane="3" entrytime="00:01:59.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="235" swimtime="00:02:00.90" resultid="15111" heatid="15648" lane="6" entrytime="00:01:55.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sylwia" lastname="Gorockiewicz" birthdate="1975-03-29" gender="F" nation="POL" license="500115600525" swrid="4837788" athleteid="15102">
              <RESULTS>
                <RESULT eventid="1053" points="208" swimtime="00:04:45.40" resultid="15103" heatid="15550" lane="1" entrytime="00:04:41.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.48" />
                    <SPLIT distance="100" swimtime="00:02:16.65" />
                    <SPLIT distance="150" swimtime="00:03:32.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="114" swimtime="00:01:01.86" resultid="15104" heatid="15578" lane="4" />
                <RESULT eventid="1198" points="212" swimtime="00:02:09.92" resultid="15105" heatid="15622" lane="5" entrytime="00:02:10.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="96" swimtime="00:02:09.84" resultid="15106" heatid="15649" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewa" lastname="Szała" birthdate="1959-03-19" gender="F" nation="POL" license="500115600674" swrid="4302573" athleteid="15117">
              <RESULTS>
                <RESULT eventid="1105" points="772" swimtime="00:01:28.40" resultid="15118" heatid="15571" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="591" swimtime="00:02:54.83" resultid="15119" heatid="15587" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.62" />
                    <SPLIT distance="100" swimtime="00:01:24.30" />
                    <SPLIT distance="150" swimtime="00:02:09.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5430" points="759" swimtime="00:03:11.11" resultid="15120" heatid="15616" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.52" />
                    <SPLIT distance="100" swimtime="00:01:32.77" />
                    <SPLIT distance="150" swimtime="00:02:22.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="583" swimtime="00:01:21.51" resultid="15121" heatid="15649" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Kotecka" birthdate="1965-05-08" gender="F" nation="POL" license="100115600357" swrid="4754727" athleteid="15122">
              <RESULTS>
                <RESULT eventid="1105" points="397" swimtime="00:01:41.22" resultid="15123" heatid="15570" lane="4" entrytime="00:01:41.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="453" swimtime="00:02:59.29" resultid="15124" heatid="15587" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.78" />
                    <SPLIT distance="100" swimtime="00:01:27.19" />
                    <SPLIT distance="150" swimtime="00:02:13.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5430" points="399" swimtime="00:03:33.29" resultid="15125" heatid="15614" lane="1" entrytime="00:03:28.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.34" />
                    <SPLIT distance="100" swimtime="00:01:43.60" />
                    <SPLIT distance="150" swimtime="00:02:39.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="421" swimtime="00:01:23.63" resultid="15126" heatid="15650" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabela" lastname="Skurczyńska" birthdate="1971-10-13" gender="F" nation="POL" license="500115600746" athleteid="15099">
              <RESULTS>
                <RESULT eventid="1053" points="348" swimtime="00:03:58.94" resultid="15100" heatid="15549" lane="6" entrytime="00:03:57.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.08" />
                    <SPLIT distance="100" swimtime="00:01:52.03" />
                    <SPLIT distance="150" swimtime="00:02:56.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="394" swimtime="00:00:48.82" resultid="15101" heatid="15602" lane="6" entrytime="00:00:48.55" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04303" nation="POL" region="03" clubid="15134" name="Masters Avia Świdnik">
          <ATHLETES>
            <ATHLETE firstname="Cezary" lastname="Lipiński" birthdate="1972-04-11" gender="M" nation="POL" license="104303700002" swrid="5449345" athleteid="15135">
              <RESULTS>
                <RESULT eventid="1092" points="620" swimtime="00:00:28.72" resultid="15136" heatid="15562" lane="6" entrytime="00:00:28.27" entrycourse="SCM" />
                <RESULT eventid="1170" points="543" swimtime="00:02:24.76" resultid="15137" heatid="15588" lane="6" entrytime="00:02:20.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                    <SPLIT distance="100" swimtime="00:01:09.35" />
                    <SPLIT distance="150" swimtime="00:01:47.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="406" swimtime="00:00:38.30" resultid="15138" heatid="15640" lane="5" />
                <RESULT eventid="1238" points="554" swimtime="00:01:04.64" resultid="15139" heatid="15652" lane="3" entrytime="00:01:02.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jakub" lastname="Kozłowski" birthdate="1982-07-01" gender="M" nation="POL" license="504303700014" athleteid="15140">
              <RESULTS>
                <RESULT eventid="6830" points="707" swimtime="00:00:32.63" resultid="15141" heatid="15610" lane="3" />
                <RESULT eventid="1212" points="679" swimtime="00:01:12.34" resultid="15142" heatid="15629" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="BIAŁYS" nation="POL" clubid="14562" name="MKS Juvenia Białystok">
          <ATHLETES>
            <ATHLETE firstname="Dominika" lastname="Michalik" birthdate="1979-01-01" gender="F" nation="POL" athleteid="15466">
              <RESULTS>
                <RESULT eventid="1157" points="715" swimtime="00:02:24.56" resultid="15467" heatid="15584" lane="2" entrytime="00:02:24.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                    <SPLIT distance="100" swimtime="00:01:09.83" />
                    <SPLIT distance="150" swimtime="00:01:46.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="695" swimtime="00:01:06.01" resultid="15468" heatid="15646" lane="2" entrytime="00:01:06.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Żmiejko" birthdate="1963-01-01" gender="M" nation="POL" swrid="4186249" athleteid="14563">
              <RESULTS>
                <RESULT eventid="1092" points="783" swimtime="00:00:29.11" resultid="14564" heatid="15562" lane="1" entrytime="00:00:28.13" entrycourse="SCM" />
                <RESULT eventid="5390" points="859" swimtime="00:01:11.81" resultid="14565" heatid="15597" lane="2" entrytime="00:01:11.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="821" swimtime="00:01:03.93" resultid="14566" heatid="15652" lane="4" entrytime="00:01:02.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="08001" nation="POL" region="01" clubid="15274" name="Sport Active">
          <ATHLETES>
            <ATHLETE firstname="Wojciech" lastname="Mroczko" birthdate="1978-01-30" gender="M" nation="POL" license="508001700025" athleteid="15278">
              <RESULTS>
                <RESULT eventid="1092" points="261" swimtime="00:00:37.33" resultid="15279" heatid="15568" lane="3" />
                <RESULT eventid="1170" points="238" swimtime="00:03:05.01" resultid="15280" heatid="15591" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.74" />
                    <SPLIT distance="100" swimtime="00:01:27.72" />
                    <SPLIT distance="150" swimtime="00:02:16.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Cygal" birthdate="1980-09-10" gender="M" nation="POL" license="508001700040" athleteid="15275">
              <RESULTS>
                <RESULT eventid="1066" points="241" swimtime="00:03:49.37" resultid="15276" heatid="15555" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.13" />
                    <SPLIT distance="100" swimtime="00:01:45.96" />
                    <SPLIT distance="150" swimtime="00:02:48.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="156" swimtime="00:03:29.85" resultid="15277" heatid="15592" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.80" />
                    <SPLIT distance="100" swimtime="00:01:36.65" />
                    <SPLIT distance="150" swimtime="00:02:33.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="10414" nation="POL" region="14" clubid="15023" name="Klub Sportowy Mako">
          <ATHLETES>
            <ATHLETE firstname="Marek" lastname="Piórkowski" birthdate="1965-07-28" gender="M" nation="POL" license="510414700072" swrid="5506637" athleteid="15024">
              <RESULTS>
                <RESULT eventid="1118" points="229" swimtime="00:01:45.71" resultid="15025" heatid="15573" lane="1" entrytime="00:01:49.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="260" swimtime="00:03:18.54" resultid="15026" heatid="15590" lane="1" entrytime="00:03:21.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.65" />
                    <SPLIT distance="100" swimtime="00:01:32.49" />
                    <SPLIT distance="150" swimtime="00:02:25.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="239" swimtime="00:00:47.27" resultid="15027" heatid="15638" lane="5" entrytime="00:00:47.37" entrycourse="SCM" />
                <RESULT eventid="1238" points="313" swimtime="00:01:25.39" resultid="15028" heatid="15657" lane="2" entrytime="00:01:28.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="07611" nation="POL" region="11" clubid="15313" name="UKS DRAGON Sosnowiec">
          <ATHLETES>
            <ATHLETE firstname="Paweł" lastname="Jankowski" birthdate="1995-08-14" gender="M" nation="POL" license="107611700057" swrid="4112623" athleteid="15314">
              <RESULTS>
                <RESULT eventid="1092" points="830" swimtime="00:00:24.30" resultid="15315" heatid="15561" lane="4" entrytime="00:00:23.82" />
                <RESULT eventid="5390" points="819" swimtime="00:00:58.99" resultid="15316" heatid="15596" lane="3" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="884" swimtime="00:00:26.10" resultid="15317" heatid="15635" lane="3" entrytime="00:00:26.07" />
                <RESULT eventid="1238" points="822" swimtime="00:00:51.85" resultid="15318" heatid="15651" lane="3" entrytime="00:00:51.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOTYL" nation="POL" clubid="14557" name="Motyl Mosir Stalowa Wola">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Petecka" birthdate="1967-04-17" gender="F" nation="POL" swrid="4992840" athleteid="14558">
              <RESULTS>
                <RESULT eventid="1053" points="568" swimtime="00:03:43.70" resultid="14559" heatid="15549" lane="5" entrytime="00:03:38.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.53" />
                    <SPLIT distance="100" swimtime="00:01:47.12" />
                    <SPLIT distance="150" swimtime="00:02:45.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="446" swimtime="00:00:41.80" resultid="14560" heatid="15576" lane="5" entrytime="00:00:42.00" />
                <RESULT eventid="1198" points="502" swimtime="00:01:44.69" resultid="14561" heatid="15621" lane="4" entrytime="00:01:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="03311" nation="POL" clubid="14699" name="Uks Wodnik 29 Katowice">
          <ATHLETES>
            <ATHLETE firstname="Michał" lastname="Spławiński" birthdate="1981-05-16" gender="M" nation="POL" swrid="4060309" athleteid="14700">
              <RESULTS>
                <RESULT eventid="1144" points="724" swimtime="00:00:27.98" resultid="14701" heatid="15579" lane="1" entrytime="00:00:28.90" />
                <RESULT eventid="6830" points="761" swimtime="00:00:31.84" resultid="14702" heatid="15605" lane="1" entrytime="00:00:32.50" />
                <RESULT eventid="1212" points="703" swimtime="00:01:11.51" resultid="14703" heatid="15624" lane="6" entrytime="00:01:14.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="655" swimtime="00:00:59.02" resultid="14704" heatid="15652" lane="1" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZOLES" nation="POL" region="01" clubid="15472" name="NZ Oleśnica">
          <ATHLETES>
            <ATHLETE firstname="Piotr" lastname="Krzekotowski" birthdate="1966-01-01" gender="M" nation="POL" swrid="5416779" athleteid="15002">
              <RESULTS>
                <RESULT eventid="1066" points="343" swimtime="00:03:51.32" resultid="15003" heatid="15554" lane="2" entrytime="00:03:59.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.62" />
                    <SPLIT distance="100" swimtime="00:01:50.00" />
                    <SPLIT distance="150" swimtime="00:02:49.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="257" swimtime="00:03:19.29" resultid="15004" heatid="15591" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.05" />
                    <SPLIT distance="100" swimtime="00:01:35.66" />
                    <SPLIT distance="150" swimtime="00:03:18.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5417" points="179" swimtime="00:01:51.76" resultid="15005" heatid="15645" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="304" swimtime="00:01:26.23" resultid="15006" heatid="15658" lane="3" entrytime="00:01:32.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="GÓRRAD" nation="POL" clubid="14526" name="Górnik Radlin">
          <ATHLETES>
            <ATHLETE firstname="Marian" lastname="Otlik" birthdate="1966-09-08" gender="M" nation="POL" swrid="4831502" athleteid="14527">
              <RESULTS>
                <RESULT eventid="1144" points="402" swimtime="00:00:37.99" resultid="14528" heatid="15581" lane="3" entrytime="00:00:36.40" entrycourse="SCM" />
                <RESULT eventid="5390" points="432" swimtime="00:01:26.92" resultid="14529" heatid="15598" lane="6" entrytime="00:01:25.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="295" swimtime="00:01:42.30" resultid="14530" heatid="15629" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5417" points="337" swimtime="00:01:30.60" resultid="14531" heatid="15645" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" clubid="15774" name="Aqua Sfera Masters Olsztyn">
          <ATHLETES>
            <ATHLETE firstname="Mieszko" lastname="Palmi-Kukiełko" birthdate="1993-09-15" gender="M" nation="POL" license="101713700006" swrid="4073437" athleteid="15020">
              <RESULTS>
                <RESULT eventid="1066" points="688" swimtime="00:02:39.12" resultid="15021" heatid="15552" lane="2" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                    <SPLIT distance="100" swimtime="00:01:14.65" />
                    <SPLIT distance="150" swimtime="00:01:56.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="599" swimtime="00:02:06.36" resultid="15022" heatid="15588" lane="4" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.23" />
                    <SPLIT distance="100" swimtime="00:01:01.26" />
                    <SPLIT distance="150" swimtime="00:01:34.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="8CHRZ" nation="POL" clubid="14538" name="Uks Sp 8 Chrzanów">
          <ATHLETES>
            <ATHLETE firstname="Alfred" lastname="Zabrzański" birthdate="1954-05-12" gender="M" nation="POL" swrid="4477631" athleteid="14539">
              <RESULTS>
                <RESULT eventid="1092" points="554" swimtime="00:00:33.57" resultid="14540" heatid="15564" lane="1" entrytime="00:00:32.97" entrycourse="SCM" />
                <RESULT eventid="5390" points="369" swimtime="00:01:38.63" resultid="14541" heatid="15599" lane="4" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="434" swimtime="00:00:43.99" resultid="14542" heatid="15637" lane="6" entrytime="00:00:43.81" />
                <RESULT eventid="1238" points="526" swimtime="00:01:15.68" resultid="14543" heatid="15655" lane="5" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SLEZA" nation="POL" clubid="14879" name="Swim Club Masters Ślęza">
          <ATHLETES>
            <ATHLETE firstname="Joanna" lastname="Chojcan" birthdate="1986-08-04" gender="F" nation="POL" athleteid="15663">
              <RESULTS>
                <RESULT eventid="1105" points="645" swimtime="00:01:16.28" resultid="15664" heatid="15569" lane="4" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="529" swimtime="00:00:35.15" resultid="15665" heatid="15576" lane="4" entrytime="00:00:37.00" />
                <RESULT eventid="5430" points="613" swimtime="00:02:48.08" resultid="15666" heatid="15614" lane="4" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.71" />
                    <SPLIT distance="100" swimtime="00:01:20.34" />
                    <SPLIT distance="150" swimtime="00:02:03.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5404" points="522" swimtime="00:01:19.18" resultid="15667" heatid="15641" lane="1" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Ducki" birthdate="1967-02-03" gender="M" nation="POL" athleteid="15718">
              <RESULTS>
                <RESULT comment="O-4" eventid="1092" status="DSQ" swimtime="00:00:00.00" resultid="15719" heatid="15563" lane="2" entrytime="00:00:29.70" />
                <RESULT eventid="5390" points="555" swimtime="00:01:19.98" resultid="15720" heatid="15598" lane="4" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="537" swimtime="00:00:36.10" resultid="15721" heatid="15636" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="1238" points="635" swimtime="00:01:07.50" resultid="15722" heatid="15653" lane="5" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Perek" birthdate="1980-07-01" gender="F" nation="POL" athleteid="15689">
              <RESULTS>
                <RESULT eventid="1131" points="194" swimtime="00:00:50.57" resultid="15690" heatid="15576" lane="6" entrytime="00:00:45.00" />
                <RESULT eventid="5376" points="232" swimtime="00:01:50.74" resultid="15691" heatid="15594" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="225" swimtime="00:01:36.07" resultid="15692" heatid="15648" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Bąkowski" birthdate="1984-06-20" gender="M" nation="POL" athleteid="15709">
              <RESULTS>
                <RESULT eventid="1118" points="420" swimtime="00:01:14.65" resultid="15710" heatid="15572" lane="5" entrytime="00:01:14.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5443" points="411" swimtime="00:02:43.48" resultid="15711" heatid="15617" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.14" />
                    <SPLIT distance="100" swimtime="00:01:17.94" />
                    <SPLIT distance="150" swimtime="00:02:00.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="366" swimtime="00:00:34.21" resultid="15712" heatid="15635" lane="1" entrytime="00:00:34.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Radosław" lastname="Stefurak" birthdate="1974-09-07" gender="M" nation="POL" athleteid="15701">
              <RESULTS>
                <RESULT eventid="1066" points="488" swimtime="00:03:07.50" resultid="15702" heatid="15553" lane="3" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.51" />
                    <SPLIT distance="100" swimtime="00:01:29.19" />
                    <SPLIT distance="150" swimtime="00:02:17.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6830" points="479" swimtime="00:00:38.71" resultid="15703" heatid="15606" lane="2" entrytime="00:00:37.00" />
                <RESULT eventid="1212" points="431" swimtime="00:01:27.41" resultid="15704" heatid="15625" lane="3" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Michalczuk" birthdate="1970-03-05" gender="M" nation="POL" athleteid="15729">
              <RESULTS>
                <RESULT eventid="1092" points="384" swimtime="00:00:33.68" resultid="15730" heatid="15564" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="6830" status="DNS" swimtime="00:00:00.00" resultid="15731" heatid="15607" lane="4" entrytime="00:00:39.00" />
                <RESULT eventid="1316" status="DNS" swimtime="00:00:00.00" resultid="15732" heatid="15637" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1238" status="DNS" swimtime="00:00:00.00" resultid="15733" heatid="15654" lane="1" entrytime="00:01:13.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Hanuza" birthdate="1984-06-17" gender="M" nation="POL" athleteid="15739">
              <RESULTS>
                <RESULT eventid="1144" points="531" swimtime="00:00:29.18" resultid="15740" heatid="15579" lane="6" entrytime="00:00:28.95" />
                <RESULT eventid="1170" points="522" swimtime="00:02:18.44" resultid="15741" heatid="15588" lane="1" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                    <SPLIT distance="100" swimtime="00:01:07.23" />
                    <SPLIT distance="150" swimtime="00:01:43.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnieszka" lastname="Dusza" birthdate="1983-10-11" gender="F" nation="POL" athleteid="15684">
              <RESULTS>
                <RESULT eventid="1157" status="DNS" swimtime="00:00:00.00" resultid="15685" heatid="15585" lane="1" entrytime="00:02:58.00" />
                <RESULT eventid="5376" status="DNS" swimtime="00:00:00.00" resultid="15686" heatid="15593" lane="1" entrytime="00:01:34.00" />
                <RESULT eventid="5404" status="DNS" swimtime="00:00:00.00" resultid="15687" heatid="15642" lane="2" entrytime="00:01:35.00" />
                <RESULT eventid="1225" status="DNS" swimtime="00:00:00.00" resultid="15688" heatid="15647" lane="5" entrytime="00:01:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dorota" lastname="Batóg" birthdate="1972-03-11" gender="F" nation="POL" athleteid="15734">
              <RESULTS>
                <RESULT eventid="1079" points="573" swimtime="00:00:34.06" resultid="15735" heatid="15558" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="5376" points="462" swimtime="00:01:29.27" resultid="15736" heatid="15594" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="421" swimtime="00:00:41.73" resultid="15737" heatid="15632" lane="4" entrytime="00:00:42.00" />
                <RESULT eventid="5404" status="DNS" swimtime="00:00:00.00" resultid="15738" heatid="15642" lane="4" entrytime="00:01:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Kolenkiewicz" birthdate="1977-12-13" gender="M" nation="POL" athleteid="15705">
              <RESULTS>
                <RESULT eventid="1066" points="741" swimtime="00:02:43.16" resultid="15706" heatid="15552" lane="1" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                    <SPLIT distance="100" swimtime="00:01:17.14" />
                    <SPLIT distance="150" swimtime="00:01:59.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5390" points="666" swimtime="00:01:08.68" resultid="15707" heatid="15596" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="15708" heatid="15624" lane="1" entrytime="00:01:14.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta" lastname="Burandt" birthdate="1972-01-01" gender="F" nation="POL" athleteid="15668">
              <RESULTS>
                <RESULT eventid="1131" points="565" swimtime="00:00:37.67" resultid="15669" heatid="15576" lane="2" entrytime="00:00:37.15" />
                <RESULT eventid="1157" points="498" swimtime="00:02:48.95" resultid="15670" heatid="15584" lane="6" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.64" />
                    <SPLIT distance="100" swimtime="00:01:18.08" />
                    <SPLIT distance="150" swimtime="00:02:02.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="545" swimtime="00:01:14.57" resultid="15671" heatid="15647" lane="3" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paweł" lastname="Chudoba" birthdate="1981-03-04" gender="M" nation="POL" athleteid="15697">
              <RESULTS>
                <RESULT eventid="1144" points="675" swimtime="00:00:28.64" resultid="15698" heatid="15579" lane="2" entrytime="00:00:28.50" />
                <RESULT eventid="5390" points="600" swimtime="00:01:10.89" resultid="15699" heatid="15596" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5417" points="673" swimtime="00:01:04.60" resultid="15700" heatid="15643" lane="5" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolina" lastname="Wawrzyńczak" birthdate="1990-09-11" gender="F" nation="POL" athleteid="15675">
              <RESULTS>
                <RESULT eventid="1105" points="590" swimtime="00:01:16.65" resultid="15676" heatid="15569" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="546" swimtime="00:00:34.49" resultid="15677" heatid="15575" lane="1" entrytime="00:00:34.00" />
                <RESULT eventid="1303" points="609" swimtime="00:00:35.18" resultid="15678" heatid="15631" lane="4" entrytime="00:00:35.60" />
                <RESULT eventid="5404" points="512" swimtime="00:01:18.23" resultid="15679" heatid="15641" lane="5" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oksana" lastname="Fiedor-Wojciechowska" birthdate="1975-05-22" gender="F" nation="POL" athleteid="15680">
              <RESULTS>
                <RESULT eventid="1183" points="397" swimtime="00:00:47.30" resultid="15681" heatid="15603" lane="4" entrytime="00:00:55.00" />
                <RESULT eventid="1198" points="407" swimtime="00:01:44.61" resultid="15682" heatid="15621" lane="5" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="199" swimtime="00:00:52.14" resultid="15683" heatid="15632" lane="5" entrytime="00:00:47.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Podulka" birthdate="1975-02-02" gender="F" nation="POL" athleteid="15672">
              <RESULTS>
                <RESULT eventid="1079" points="610" swimtime="00:00:31.73" resultid="15673" heatid="15557" lane="1" entrytime="00:00:32.16" />
                <RESULT eventid="1131" points="523" swimtime="00:00:37.26" resultid="15674" heatid="15576" lane="3" entrytime="00:00:36.38" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dawid" lastname="Ogorzałek" birthdate="1977-04-04" gender="M" nation="POL" athleteid="15727">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="15728" heatid="15566" lane="6" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Romanowicz" birthdate="1975-05-16" gender="M" nation="POL" athleteid="15693">
              <RESULTS>
                <RESULT eventid="1092" points="394" swimtime="00:00:32.55" resultid="15694" heatid="15565" lane="6" entrytime="00:00:35.00" />
                <RESULT comment="K-1" eventid="6830" status="DSQ" swimtime="00:00:00.00" resultid="15695" heatid="15608" lane="5" entrytime="00:00:45.00" />
                <RESULT eventid="1316" points="337" swimtime="00:00:40.04" resultid="15696" heatid="15636" lane="1" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Wójcik" birthdate="1981-02-02" gender="M" nation="POL" athleteid="15713">
              <RESULTS>
                <RESULT eventid="1092" points="349" swimtime="00:00:32.94" resultid="15714" heatid="15564" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="1170" points="219" swimtime="00:03:07.36" resultid="15715" heatid="15589" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                    <SPLIT distance="100" swimtime="00:01:25.95" />
                    <SPLIT distance="150" swimtime="00:02:16.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="191" swimtime="00:00:47.07" resultid="15716" heatid="15637" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1238" points="279" swimtime="00:01:18.44" resultid="15717" heatid="15655" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wojciech" lastname="Basiuk" birthdate="1968-03-14" gender="M" nation="POL" athleteid="15723">
              <RESULTS>
                <RESULT eventid="1092" points="220" swimtime="00:00:43.09" resultid="15724" heatid="15566" lane="2" entrytime="00:00:37.00" />
                <RESULT eventid="1144" points="196" swimtime="00:00:48.23" resultid="15725" heatid="15581" lane="1" entrytime="00:00:40.00" />
                <RESULT eventid="1238" points="273" swimtime="00:01:29.43" resultid="15726" heatid="15657" lane="4" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="6828" swimtime="00:01:58.39" resultid="15742" heatid="15612" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.71" />
                    <SPLIT distance="100" swimtime="00:00:58.96" />
                    <SPLIT distance="150" swimtime="00:01:26.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15697" number="1" />
                    <RELAYPOSITION athleteid="15663" number="2" />
                    <RELAYPOSITION athleteid="15705" number="3" />
                    <RELAYPOSITION athleteid="15672" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1290" swimtime="00:02:16.69" resultid="15746" heatid="15661" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                    <SPLIT distance="100" swimtime="00:01:15.72" />
                    <SPLIT distance="150" swimtime="00:01:44.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15705" number="1" />
                    <RELAYPOSITION athleteid="15663" number="2" />
                    <RELAYPOSITION athleteid="15697" number="3" />
                    <RELAYPOSITION athleteid="15672" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="6828" swimtime="00:02:04.86" resultid="15745" heatid="15611" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                    <SPLIT distance="100" swimtime="00:01:02.16" />
                    <SPLIT distance="150" swimtime="00:01:31.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15709" number="1" />
                    <RELAYPOSITION athleteid="15675" number="2" />
                    <RELAYPOSITION athleteid="15718" number="3" />
                    <RELAYPOSITION athleteid="15668" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1290" swimtime="00:02:24.94" resultid="15749" heatid="15661" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.70" />
                    <SPLIT distance="100" swimtime="00:01:17.93" />
                    <SPLIT distance="150" swimtime="00:01:51.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15718" number="1" />
                    <RELAYPOSITION athleteid="15693" number="2" />
                    <RELAYPOSITION athleteid="15675" number="3" />
                    <RELAYPOSITION athleteid="15668" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="6828" swimtime="00:02:21.90" resultid="15744" heatid="15611" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                    <SPLIT distance="100" swimtime="00:01:06.89" />
                    <SPLIT distance="150" swimtime="00:01:49.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15734" number="1" />
                    <RELAYPOSITION athleteid="15693" number="2" />
                    <RELAYPOSITION athleteid="15680" number="3" />
                    <RELAYPOSITION athleteid="15701" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1290" swimtime="00:03:03.92" resultid="15747" heatid="15661" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.60" />
                    <SPLIT distance="100" swimtime="00:01:42.12" />
                    <SPLIT distance="150" swimtime="00:02:33.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15689" number="1" />
                    <RELAYPOSITION athleteid="15680" number="2" />
                    <RELAYPOSITION athleteid="15723" number="3" />
                    <RELAYPOSITION athleteid="15727" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="ZDZIE" nation="POL" clubid="15007" name="MASTERS Zdzieszowice">
          <ATHLETES>
            <ATHLETE firstname="Dorota" lastname="Woźniak" birthdate="1973-09-18" gender="F" nation="POL" swrid="4992846" athleteid="15008">
              <RESULTS>
                <RESULT eventid="1105" points="506" swimtime="00:01:24.25" resultid="15009" heatid="15569" lane="1" entrytime="00:01:24.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5376" points="537" swimtime="00:01:24.92" resultid="15010" heatid="15593" lane="2" entrytime="00:01:25.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5430" points="504" swimtime="00:03:04.43" resultid="15011" heatid="15614" lane="2" entrytime="00:03:03.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.59" />
                    <SPLIT distance="100" swimtime="00:01:29.91" />
                    <SPLIT distance="150" swimtime="00:02:17.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5404" points="482" swimtime="00:01:26.22" resultid="15012" heatid="15641" lane="6" entrytime="00:01:27.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LARISW" nation="POL" clubid="14822" name="Lub. Akademia Rat. i Sportów Wod.">
          <ATHLETES>
            <ATHLETE firstname="Paweł" lastname="Krupiński" birthdate="1987-02-05" gender="M" nation="POL" swrid="5568771" athleteid="14823">
              <RESULTS>
                <RESULT eventid="1066" points="261" swimtime="00:03:39.87" resultid="14824" heatid="15553" lane="6" entrytime="00:03:38.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.81" />
                    <SPLIT distance="100" swimtime="00:01:42.50" />
                    <SPLIT distance="150" swimtime="00:02:40.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5390" points="230" swimtime="00:01:32.66" resultid="14825" heatid="15599" lane="5" entrytime="00:01:34.12" entrycourse="SCM" />
                <RESULT eventid="1212" points="264" swimtime="00:01:38.91" resultid="14826" heatid="15627" lane="4" entrytime="00:01:40.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5417" points="193" swimtime="00:01:35.45" resultid="14827" heatid="15645" lane="3" entrytime="00:01:59.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02211" nation="POL" region="11" clubid="15149" name="MUKS Gilus Gilowice">
          <ATHLETES>
            <ATHLETE firstname="Sławomir" lastname="Formas" birthdate="1969-11-05" gender="M" nation="POL" license="502211700187" swrid="4292540" athleteid="15150">
              <RESULTS>
                <RESULT eventid="1066" points="1048" swimtime="00:02:32.30" resultid="15151" heatid="15552" lane="4" entrytime="00:02:30.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                    <SPLIT distance="100" swimtime="00:01:10.99" />
                    <SPLIT distance="150" swimtime="00:01:50.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6830" points="956" swimtime="00:00:31.22" resultid="15152" heatid="15605" lane="2" entrytime="00:00:30.65" entrycourse="SCM" />
                <RESULT eventid="1212" points="980" swimtime="00:01:07.60" resultid="15153" heatid="15624" lane="4" entrytime="00:01:07.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="713" swimtime="00:00:59.40" resultid="15154" heatid="15659" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00612" nation="POL" region="12" clubid="15089" name="KS KSZO Ostrowiec Św.">
          <ATHLETES>
            <ATHLETE firstname="Stanisław" lastname="Sejmicki" birthdate="1961-05-04" gender="M" nation="POL" license="500612700426" swrid="5558380" athleteid="15090">
              <RESULTS>
                <RESULT eventid="1066" points="441" swimtime="00:03:37.97" resultid="15091" heatid="15554" lane="4" entrytime="00:03:44.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.94" />
                    <SPLIT distance="100" swimtime="00:01:44.94" />
                    <SPLIT distance="150" swimtime="00:02:41.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6830" points="429" swimtime="00:00:43.39" resultid="15092" heatid="15608" lane="2" entrytime="00:00:44.35" entrycourse="SCM" />
                <RESULT eventid="1212" points="443" swimtime="00:01:36.87" resultid="15093" heatid="15626" lane="6" entrytime="00:01:37.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DWCZ" nation="POL" clubid="14706" name="UKS Dwójeczka Częstochowa">
          <ATHLETES>
            <ATHLETE firstname="Ireneusz" lastname="Stachurski" birthdate="1969-07-22" gender="M" nation="POL" swrid="5464094" athleteid="14707">
              <RESULTS>
                <RESULT eventid="1118" points="243" swimtime="00:01:36.91" resultid="14708" heatid="15573" lane="4" entrytime="00:01:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="295" swimtime="00:02:57.36" resultid="14709" heatid="15589" lane="1" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                    <SPLIT distance="100" swimtime="00:01:24.46" />
                    <SPLIT distance="150" swimtime="00:02:12.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5417" points="193" swimtime="00:01:43.08" resultid="14710" heatid="15644" lane="2" entrytime="00:01:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" status="DNS" swimtime="00:00:00.00" resultid="14711" heatid="15656" lane="4" entrytime="00:01:18.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="701" nation="POL" clubid="14675" name="MKS 9 Dzierżoniów">
          <ATHLETES>
            <ATHLETE firstname="Rafał" lastname="Kwaśny" birthdate="1984-04-02" gender="M" nation="POL" athleteid="14688">
              <RESULTS>
                <RESULT eventid="1066" points="306" swimtime="00:03:28.49" resultid="14689" heatid="15555" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.71" />
                    <SPLIT distance="100" swimtime="00:01:38.58" />
                    <SPLIT distance="150" swimtime="00:02:34.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6830" points="285" swimtime="00:00:43.82" resultid="14690" heatid="15610" lane="2" />
                <RESULT eventid="1212" points="296" swimtime="00:01:35.20" resultid="14691" heatid="15628" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ryszard" lastname="Gendziel" birthdate="1986-03-19" gender="M" nation="POL" athleteid="14683">
              <RESULTS>
                <RESULT eventid="1092" points="394" swimtime="00:00:30.05" resultid="14684" heatid="15567" lane="1" />
                <RESULT eventid="1144" points="317" swimtime="00:00:34.63" resultid="14685" heatid="15583" lane="3" />
                <RESULT eventid="1316" points="236" swimtime="00:00:39.58" resultid="14686" heatid="15640" lane="2" />
                <RESULT eventid="1238" points="312" swimtime="00:01:12.79" resultid="14687" heatid="15658" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agata" lastname="Nowak" birthdate="1977-04-09" gender="F" nation="POL" athleteid="14678">
              <RESULTS>
                <RESULT eventid="1079" points="480" swimtime="00:00:34.36" resultid="14679" heatid="15557" lane="6" entrytime="00:00:32.58" />
                <RESULT eventid="1157" points="441" swimtime="00:02:51.31" resultid="14680" heatid="15584" lane="3" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.89" />
                    <SPLIT distance="100" swimtime="00:01:20.32" />
                    <SPLIT distance="150" swimtime="00:02:05.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="485" swimtime="00:01:38.62" resultid="14681" heatid="15620" lane="6" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="483" swimtime="00:01:16.00" resultid="14682" heatid="15647" lane="4" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dariusz" lastname="Piec" birthdate="1962-01-23" gender="M" nation="POL" athleteid="14692">
              <RESULTS>
                <RESULT eventid="1118" points="312" swimtime="00:01:39.66" resultid="14693" heatid="15573" lane="2" entrytime="00:01:43.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="367" swimtime="00:03:10.48" resultid="14694" heatid="15590" lane="4" entrytime="00:03:02.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.81" />
                    <SPLIT distance="100" swimtime="00:01:29.56" />
                    <SPLIT distance="150" swimtime="00:02:19.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5443" points="364" swimtime="00:03:39.82" resultid="14695" heatid="15618" lane="2" entrytime="00:03:45.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.27" />
                    <SPLIT distance="100" swimtime="00:01:47.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="355" swimtime="00:01:24.48" resultid="14696" heatid="15657" lane="3" entrytime="00:01:24.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewa" lastname="Fit" birthdate="1982-10-28" gender="F" nation="POL" athleteid="14676">
              <RESULTS>
                <RESULT eventid="1105" points="570" swimtime="00:01:21.96" resultid="14677" heatid="15569" lane="2" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zuzanna" lastname="Pisarska" birthdate="1981-11-06" gender="F" nation="POL" license="100701600113" swrid="5464072" athleteid="15144">
              <RESULTS>
                <RESULT eventid="1079" points="869" swimtime="00:00:27.53" resultid="15145" heatid="15557" lane="4" entrytime="00:00:27.38" entrycourse="SCM" />
                <RESULT comment="Wynik plepszy od rekordu Polski" eventid="1131" points="1031" swimtime="00:00:29.00" resultid="15146" heatid="15575" lane="4" entrytime="00:00:29.09" entrycourse="SCM" />
                <RESULT comment="Wynik lepszy od rekordu Polski" eventid="1303" points="951" swimtime="00:00:31.06" resultid="15147" heatid="15631" lane="3" entrytime="00:00:31.09" entrycourse="SCM" />
                <RESULT comment="Wynik lepszy od rekordu Polski" eventid="5404" points="892" swimtime="00:01:07.10" resultid="15148" heatid="15641" lane="4" entrytime="00:01:07.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="6828" swimtime="00:02:05.85" resultid="14697" heatid="15611" lane="3" entrytime="00:01:59.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                    <SPLIT distance="100" swimtime="00:01:08.11" />
                    <SPLIT distance="150" swimtime="00:01:38.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14676" number="1" />
                    <RELAYPOSITION athleteid="14688" number="2" />
                    <RELAYPOSITION athleteid="14683" number="3" />
                    <RELAYPOSITION athleteid="15144" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1290" swimtime="00:02:23.18" resultid="15460" heatid="15661" lane="4" entrytime="00:02:15.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                    <SPLIT distance="100" swimtime="00:01:13.18" />
                    <SPLIT distance="150" swimtime="00:01:49.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15144" number="1" />
                    <RELAYPOSITION athleteid="14688" number="2" />
                    <RELAYPOSITION athleteid="14683" number="3" />
                    <RELAYPOSITION athleteid="14678" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="15469" name="5Styl Warszawa">
          <ATHLETES>
            <ATHLETE firstname="Andrzej" lastname="Dubiel" birthdate="1987-01-15" gender="M" nation="POL" athleteid="15470">
              <RESULTS>
                <RESULT eventid="1092" points="707" swimtime="00:00:24.72" resultid="15471" heatid="15561" lane="1" entrytime="00:00:25.50" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00607" nation="POL" region="07" clubid="15281" name="Towarzystwo Pływackie ,,Masters&apos;&apos; Opole">
          <ATHLETES>
            <ATHLETE firstname="Jerzy" lastname="Minkiewicz" birthdate="1956-05-31" gender="M" nation="POL" license="100607700031" swrid="4183581" athleteid="15282">
              <RESULTS>
                <RESULT eventid="1092" points="545" swimtime="00:00:33.76" resultid="15283" heatid="15565" lane="4" entrytime="00:00:34.00" />
                <RESULT eventid="1144" points="446" swimtime="00:00:39.99" resultid="15284" heatid="15580" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="1316" points="418" swimtime="00:00:44.56" resultid="15285" heatid="15637" lane="5" entrytime="00:00:41.00" />
                <RESULT eventid="1238" points="460" swimtime="00:01:19.16" resultid="15286" heatid="15654" lane="6" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Vogel" birthdate="1981-09-20" gender="M" nation="POL" license="100607700016" swrid="5506641" athleteid="15299">
              <RESULTS>
                <RESULT eventid="1144" points="625" swimtime="00:00:29.39" resultid="15300" heatid="15579" lane="5" entrytime="00:00:28.87" entrycourse="SCM" />
                <RESULT eventid="5390" points="592" swimtime="00:01:11.24" resultid="15301" heatid="15597" lane="3" entrytime="00:01:10.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Mandziuk" birthdate="1965-04-11" gender="M" nation="POL" license="100607700033" athleteid="15287">
              <RESULTS>
                <RESULT eventid="1092" points="337" swimtime="00:00:37.40" resultid="15288" heatid="15565" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="6830" points="186" swimtime="00:00:53.35" resultid="15289" heatid="15609" lane="3" entrytime="00:00:52.00" />
                <RESULT eventid="1212" points="173" swimtime="00:02:02.22" resultid="15290" heatid="15628" lane="4" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="331" swimtime="00:01:23.82" resultid="15291" heatid="15656" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zbigniew" lastname="Januszkiewicz" birthdate="1962-08-18" gender="M" nation="POL" license="100607700003" swrid="4843497" athleteid="15292">
              <RESULTS>
                <RESULT eventid="1118" status="DNS" swimtime="00:00:00.00" resultid="15293" heatid="15572" lane="3" entrytime="00:01:05.46" entrycourse="SCM" />
                <RESULT eventid="1144" points="971" swimtime="00:00:29.43" resultid="15294" heatid="15580" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="5390" points="974" swimtime="00:01:08.88" resultid="15295" heatid="15597" lane="1" entrytime="00:01:11.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5443" points="1225" swimtime="00:02:26.74" resultid="15296" heatid="15617" lane="3" entrytime="00:02:23.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                    <SPLIT distance="100" swimtime="00:01:12.54" />
                    <SPLIT distance="150" swimtime="00:01:49.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" status="DNS" swimtime="00:00:00.00" resultid="15297" heatid="15635" lane="4" entrytime="00:00:30.77" entrycourse="SCM" />
                <RESULT eventid="1238" points="996" swimtime="00:00:59.94" resultid="15298" heatid="15652" lane="2" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KRAK" nation="POL" clubid="14756" name="JK TEAM Kraków">
          <ATHLETES>
            <ATHLETE firstname="Agata" lastname="Jasik" birthdate="1984-01-01" gender="F" nation="POL" swrid="5484408" athleteid="14757">
              <RESULTS>
                <RESULT eventid="1079" points="355" swimtime="00:00:36.95" resultid="14758" heatid="15558" lane="3" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1157" points="388" swimtime="00:02:55.66" resultid="14759" heatid="15585" lane="2" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.19" />
                    <SPLIT distance="100" swimtime="00:01:23.06" />
                    <SPLIT distance="150" swimtime="00:02:09.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ryszard" lastname="Zając" birthdate="1984-01-01" gender="M" nation="POL" swrid="5468089" athleteid="14760">
              <RESULTS>
                <RESULT eventid="1092" points="266" swimtime="00:00:34.23" resultid="14761" heatid="15565" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="5390" points="203" swimtime="00:01:36.61" resultid="14762" heatid="15599" lane="1" entrytime="00:01:40.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="04214" nation="POL" region="14" clubid="15319" name="Warsaw Masters Team">
          <ATHLETES>
            <ATHLETE firstname="Leszek" lastname="Madej" birthdate="1960-06-17" gender="M" nation="POL" license="504214700005" swrid="4183799" athleteid="15325">
              <RESULTS>
                <RESULT eventid="1092" points="867" swimtime="00:00:28.14" resultid="15326" heatid="15562" lane="3" entrytime="00:00:27.89" entrycourse="SCM" />
                <RESULT eventid="5390" points="876" swimtime="00:01:11.34" resultid="15327" heatid="15597" lane="4" entrytime="00:01:11.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="790" swimtime="00:01:19.90" resultid="15328" heatid="15630" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="926" swimtime="00:01:01.42" resultid="15329" heatid="15652" lane="5" entrytime="00:01:02.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Skośkiewicz" birthdate="1966-05-05" gender="M" nation="POL" license="504214700002" swrid="4183802" athleteid="15330">
              <RESULTS>
                <RESULT eventid="1118" points="788" swimtime="00:01:10.10" resultid="15331" heatid="15572" lane="4" entrytime="00:01:10.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5390" points="869" swimtime="00:01:08.87" resultid="15332" heatid="15596" lane="6" entrytime="00:01:10.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="724" swimtime="00:00:32.68" resultid="15333" heatid="15635" lane="2" entrytime="00:00:32.30" entrycourse="SCM" />
                <RESULT eventid="5417" points="751" swimtime="00:01:09.39" resultid="15334" heatid="15643" lane="6" entrytime="00:01:10.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bartosz" lastname="Ostrowski" birthdate="1977-05-14" gender="M" nation="POL" license="504214700091" swrid="5506635" athleteid="15320">
              <RESULTS>
                <RESULT eventid="1066" points="588" swimtime="00:02:56.19" resultid="15321" heatid="15552" lane="6" entrytime="00:02:48.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.46" />
                    <SPLIT distance="100" swimtime="00:01:20.46" />
                    <SPLIT distance="150" swimtime="00:02:08.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6830" points="833" swimtime="00:00:32.19" resultid="15322" heatid="15605" lane="5" entrytime="00:00:31.89" entrycourse="SCM" />
                <RESULT eventid="1212" points="737" swimtime="00:01:13.12" resultid="15323" heatid="15624" lane="2" entrytime="00:01:10.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" status="DNS" swimtime="00:00:00.00" resultid="15324" heatid="15651" lane="6" entrytime="00:00:59.13" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="REKIN" nation="POL" region="01" clubid="14597" name="KS REKIN Świebodzice">
          <ATHLETES>
            <ATHLETE firstname="Maciej" lastname="Jaroński" birthdate="1991-05-09" gender="M" nation="POL" swrid="4192553" athleteid="14598">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="14599" heatid="15563" lane="5" entrytime="00:00:30.11" />
                <RESULT eventid="5390" status="DNS" swimtime="00:00:00.00" resultid="14600" heatid="15598" lane="2" entrytime="00:01:20.02" />
                <RESULT eventid="1212" points="342" swimtime="00:01:27.66" resultid="14601" heatid="15626" lane="4" entrytime="00:01:35.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="419" swimtime="00:00:35.39" resultid="14602" heatid="15636" lane="3" entrytime="00:00:36.19" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02805" nation="POL" region="05" clubid="15155" name="MUKS Zgierz">
          <ATHLETES>
            <ATHLETE firstname="Małgorzata" lastname="Ścibiorek" birthdate="1971-09-12" gender="F" nation="POL" license="502805600026" swrid="4992745" athleteid="15245">
              <RESULTS>
                <RESULT eventid="1131" points="861" swimtime="00:00:32.74" resultid="15246" heatid="15575" lane="2" entrytime="00:00:32.28" entrycourse="SCM" />
                <RESULT eventid="5376" points="756" swimtime="00:01:15.79" resultid="15247" heatid="15593" lane="4" entrytime="00:01:14.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5404" points="762" swimtime="00:01:14.03" resultid="15248" heatid="15641" lane="2" entrytime="00:01:12.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabela" lastname="Wypych - Staszewska" birthdate="1970-08-16" gender="F" nation="POL" license="502805600164" athleteid="15249">
              <RESULTS>
                <RESULT eventid="1131" points="485" swimtime="00:00:39.63" resultid="15250" heatid="15577" lane="5" />
                <RESULT eventid="5376" points="423" swimtime="00:01:31.95" resultid="15251" heatid="15595" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5430" points="344" swimtime="00:03:29.52" resultid="15252" heatid="15615" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.15" />
                    <SPLIT distance="100" swimtime="00:01:39.73" />
                    <SPLIT distance="150" swimtime="00:02:34.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5404" points="365" swimtime="00:01:34.60" resultid="15253" heatid="15642" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafał" lastname="Maciejewski" birthdate="1974-04-11" gender="M" nation="POL" license="502805700028" swrid="5373991" athleteid="15216">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="15217" heatid="15566" lane="3" entrytime="00:00:35.10" entrycourse="SCM" />
                <RESULT eventid="6830" status="DNS" swimtime="00:00:00.00" resultid="15218" heatid="15608" lane="4" entrytime="00:00:44.00" entrycourse="SCM" />
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="15219" heatid="15627" lane="5" entrytime="00:01:41.45" entrycourse="SCM" />
                <RESULT eventid="1238" status="DNS" swimtime="00:00:00.00" resultid="15220" heatid="15656" lane="2" entrytime="00:01:19.64" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandra" lastname="Ławniczak" birthdate="1979-09-13" gender="F" nation="POL" athleteid="14661">
              <RESULTS>
                <RESULT eventid="1079" points="268" swimtime="00:00:40.76" resultid="14662" heatid="15558" lane="1" entrytime="00:00:39.00" />
                <RESULT eventid="5376" points="271" swimtime="00:01:45.22" resultid="14663" heatid="15593" lane="6" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="232" swimtime="00:00:49.67" resultid="14664" heatid="15631" lane="1" entrytime="00:00:39.00" />
                <RESULT eventid="1225" points="258" swimtime="00:01:31.81" resultid="14665" heatid="15648" lane="4" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" lastname="Matczak" birthdate="1989-08-12" gender="M" nation="POL" license="102805700157" swrid="4071609" athleteid="15192">
              <RESULTS>
                <RESULT eventid="1066" points="915" swimtime="00:02:24.70" resultid="15193" heatid="15552" lane="3" entrytime="00:02:21.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                    <SPLIT distance="100" swimtime="00:01:10.60" />
                    <SPLIT distance="150" swimtime="00:01:47.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6830" points="766" swimtime="00:00:30.39" resultid="15194" heatid="15605" lane="4" entrytime="00:00:29.77" entrycourse="SCM" />
                <RESULT eventid="1212" points="762" swimtime="00:01:07.13" resultid="15195" heatid="15624" lane="3" entrytime="00:01:04.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robert" lastname="Szalbierz" birthdate="1968-08-06" gender="M" nation="POL" license="502805700034" swrid="5373990" athleteid="15211">
              <RESULTS>
                <RESULT eventid="1092" points="596" swimtime="00:00:30.93" resultid="15212" heatid="15564" lane="3" entrytime="00:00:30.81" entrycourse="SCM" />
                <RESULT eventid="1144" points="522" swimtime="00:00:34.82" resultid="15213" heatid="15580" lane="1" entrytime="00:00:34.23" entrycourse="SCM" />
                <RESULT comment="K-1" eventid="1212" status="DSQ" swimtime="00:00:00.00" resultid="15214" heatid="15629" lane="3" />
                <RESULT eventid="1238" points="522" swimtime="00:01:12.07" resultid="15215" heatid="15659" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Justyna" lastname="Barańska" birthdate="1977-01-05" gender="F" nation="POL" license="502805600055" swrid="4655158" athleteid="15164">
              <RESULTS>
                <RESULT eventid="1053" points="468" swimtime="00:03:37.89" resultid="15165" heatid="15549" lane="2" entrytime="00:03:36.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.06" />
                    <SPLIT distance="100" swimtime="00:01:44.67" />
                    <SPLIT distance="150" swimtime="00:02:41.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="400" swimtime="00:00:47.16" resultid="15166" heatid="15602" lane="1" entrytime="00:00:45.35" entrycourse="SCM" />
                <RESULT eventid="1198" points="435" swimtime="00:01:42.27" resultid="15167" heatid="15621" lane="3" entrytime="00:01:39.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="262" swimtime="00:00:47.60" resultid="15168" heatid="15634" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wiktor" lastname="Morozowski" birthdate="1973-05-09" gender="M" nation="POL" license="102805700051" swrid="5416829" athleteid="15187">
              <RESULTS>
                <RESULT eventid="1066" status="DNS" swimtime="00:00:00.00" resultid="15188" heatid="15553" lane="5" entrytime="00:03:27.10" entrycourse="SCM" />
                <RESULT eventid="6830" points="465" swimtime="00:00:39.70" resultid="15189" heatid="15607" lane="3" entrytime="00:00:38.93" entrycourse="SCM" />
                <RESULT eventid="1212" points="392" swimtime="00:01:31.68" resultid="15190" heatid="15630" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="386" swimtime="00:01:12.91" resultid="15191" heatid="15658" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roman" lastname="Wiczel" birthdate="1948-01-22" gender="M" nation="POL" license="502805700021" swrid="4876444" athleteid="15169">
              <RESULTS>
                <RESULT eventid="1066" points="713" swimtime="00:03:38.86" resultid="15170" heatid="15553" lane="1" entrytime="00:03:34.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.75" />
                    <SPLIT distance="100" swimtime="00:01:45.90" />
                    <SPLIT distance="150" swimtime="00:02:43.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6830" points="732" swimtime="00:00:43.48" resultid="15171" heatid="15608" lane="3" entrytime="00:00:43.37" entrycourse="SCM" />
                <RESULT comment="Wynik lepszy od rekordu Polski" eventid="1212" points="717" swimtime="00:01:36.91" resultid="15172" heatid="15626" lane="1" entrytime="00:01:37.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stanisław" lastname="Sikorski" birthdate="1951-05-03" gender="M" nation="POL" license="502805700036" swrid="5582462" athleteid="15230">
              <RESULTS>
                <RESULT eventid="1118" points="161" swimtime="00:02:17.83" resultid="15231" heatid="15574" lane="4" entrytime="00:02:07.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6830" points="309" swimtime="00:00:52.55" resultid="15232" heatid="15609" lane="4" entrytime="00:00:53.03" entrycourse="SCM" />
                <RESULT comment="K-15" eventid="1212" status="DSQ" swimtime="00:00:00.00" resultid="15233" heatid="15628" lane="2" entrytime="00:02:04.07" entrycourse="SCM" />
                <RESULT comment="O-5" eventid="1316" status="DSQ" swimtime="00:00:00.00" resultid="15234" heatid="15639" lane="4" entrytime="00:00:57.12" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dorota" lastname="Kajdos" birthdate="1976-06-25" gender="F" nation="POL" license="502805600148" swrid="5558379" athleteid="15206">
              <RESULTS>
                <RESULT eventid="1079" points="247" swimtime="00:00:42.87" resultid="15207" heatid="15560" lane="2" />
                <RESULT comment="G-8" eventid="1105" status="DSQ" swimtime="00:00:00.00" resultid="15208" heatid="15570" lane="2" entrytime="00:01:56.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5430" points="309" swimtime="00:03:47.41" resultid="15209" heatid="15615" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.70" />
                    <SPLIT distance="100" swimtime="00:01:50.97" />
                    <SPLIT distance="150" swimtime="00:02:50.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="241" swimtime="00:00:48.98" resultid="15210" heatid="15632" lane="6" entrytime="00:00:49.96" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dagmara" lastname="Luzniakowska" birthdate="1980-04-29" gender="F" nation="POL" license="102805600154" swrid="5582458" athleteid="15240">
              <RESULTS>
                <RESULT eventid="1131" points="255" swimtime="00:00:46.17" resultid="15241" heatid="15576" lane="1" entrytime="00:00:43.42" entrycourse="SCM" />
                <RESULT eventid="1157" points="406" swimtime="00:02:54.56" resultid="15242" heatid="15585" lane="5" entrytime="00:02:55.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.05" />
                    <SPLIT distance="100" swimtime="00:01:24.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="347" swimtime="00:01:47.68" resultid="15243" heatid="15623" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="415" swimtime="00:01:18.37" resultid="15244" heatid="15647" lane="1" entrytime="00:01:20.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrzej" lastname="Sypniewski" birthdate="1957-02-01" gender="M" nation="POL" license="102805700035" swrid="5373999" athleteid="15259">
              <RESULTS>
                <RESULT eventid="5390" points="564" swimtime="00:01:25.62" resultid="15260" heatid="15598" lane="5" entrytime="00:01:20.67" entrycourse="SCM" />
                <RESULT eventid="6830" points="487" swimtime="00:00:42.94" resultid="15261" heatid="15609" lane="5" />
                <RESULT eventid="1212" points="503" swimtime="00:01:36.72" resultid="15262" heatid="15626" lane="5" entrytime="00:01:37.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="577" swimtime="00:00:40.01" resultid="15263" heatid="15636" lane="2" entrytime="00:00:39.37" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zdzisław" lastname="Jasiński" birthdate="1960-07-23" gender="M" nation="POL" license="502805700027" swrid="5374015" athleteid="15182">
              <RESULTS>
                <RESULT eventid="1066" points="442" swimtime="00:03:37.72" resultid="15183" heatid="15554" lane="3" entrytime="00:03:43.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.01" />
                    <SPLIT distance="100" swimtime="00:01:45.26" />
                    <SPLIT distance="150" swimtime="00:02:43.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5390" points="401" swimtime="00:01:32.53" resultid="15184" heatid="15599" lane="2" entrytime="00:01:32.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.34" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="O-1" eventid="1212" status="DSQ" swimtime="00:00:00.00" resultid="15185" heatid="15627" lane="2" entrytime="00:01:40.89" entrycourse="SCM" />
                <RESULT eventid="1238" points="504" swimtime="00:01:15.21" resultid="15186" heatid="15655" lane="6" entrytime="00:01:17.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Pietruszewski - Gil" birthdate="1986-12-17" gender="M" nation="POL" license="502805700163" athleteid="15221">
              <RESULTS>
                <RESULT eventid="1092" points="350" swimtime="00:00:31.25" resultid="15222" heatid="15568" lane="2" />
                <RESULT eventid="5390" points="329" swimtime="00:01:22.24" resultid="15223" heatid="15601" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="351" swimtime="00:01:09.96" resultid="15224" heatid="15659" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Urszula" lastname="Mróz" birthdate="1962-03-03" gender="F" nation="POL" license="502805600024" swrid="4754660" athleteid="15196">
              <RESULTS>
                <RESULT eventid="1079" points="749" swimtime="00:00:34.14" resultid="15197" heatid="15558" lane="4" entrytime="00:00:33.30" entrycourse="SCM" />
                <RESULT eventid="1131" points="779" swimtime="00:00:36.33" resultid="15198" heatid="15575" lane="6" entrytime="00:00:35.04" entrycourse="SCM" />
                <RESULT eventid="1303" points="620" swimtime="00:00:42.56" resultid="15199" heatid="15632" lane="3" entrytime="00:00:40.40" entrycourse="SCM" />
                <RESULT eventid="1225" points="709" swimtime="00:01:16.40" resultid="15200" heatid="15647" lane="6" entrytime="00:01:22.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Piotr" lastname="Gołębiowski" birthdate="1996-05-20" gender="M" nation="POL" license="502805700155" swrid="4115580" athleteid="15225">
              <RESULTS>
                <RESULT eventid="1092" points="605" swimtime="00:00:27.00" resultid="15226" heatid="15561" lane="6" entrytime="00:00:27.61" entrycourse="SCM" />
                <RESULT eventid="6830" points="551" swimtime="00:00:34.46" resultid="15227" heatid="15605" lane="6" entrytime="00:00:35.23" entrycourse="SCM" />
                <RESULT eventid="1212" points="542" swimtime="00:01:16.04" resultid="15228" heatid="15629" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="549" swimtime="00:00:59.31" resultid="15229" heatid="15660" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Dziedziczak" birthdate="1977-02-04" gender="M" nation="POL" license="502805700153" swrid="5558378" athleteid="15235">
              <RESULTS>
                <RESULT eventid="1118" points="265" swimtime="00:01:32.46" resultid="15236" heatid="15574" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5390" points="344" swimtime="00:01:25.60" resultid="15237" heatid="15598" lane="1" entrytime="00:01:22.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5443" points="305" swimtime="00:03:15.44" resultid="15238" heatid="15619" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="420" swimtime="00:01:10.61" resultid="15239" heatid="15654" lane="4" entrytime="00:01:11.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" lastname="Rembowska-Świeboda" birthdate="1968-06-27" gender="F" nation="POL" license="102805600031" swrid="5439505" athleteid="15201">
              <RESULTS>
                <RESULT eventid="1079" points="609" swimtime="00:00:33.88" resultid="15202" heatid="15558" lane="5" entrytime="00:00:34.90" entrycourse="SCM" />
                <RESULT eventid="1105" points="696" swimtime="00:01:23.96" resultid="15203" heatid="15571" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="682" swimtime="00:00:38.45" resultid="15204" heatid="15631" lane="5" entrytime="00:00:38.96" entrycourse="SCM" />
                <RESULT eventid="1225" points="570" swimtime="00:01:15.63" resultid="15205" heatid="15650" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" lastname="Ścibiorek" birthdate="1997-02-19" gender="M" nation="POL" swrid="4287843" athleteid="14657">
              <RESULTS>
                <RESULT eventid="1092" points="661" swimtime="00:00:26.21" resultid="14658" heatid="15561" lane="2" entrytime="00:00:25.00" />
                <RESULT eventid="1170" points="616" swimtime="00:02:10.61" resultid="14659" heatid="15588" lane="5" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.89" />
                    <SPLIT distance="100" swimtime="00:01:02.34" />
                    <SPLIT distance="150" swimtime="00:01:36.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="591" swimtime="00:00:57.86" resultid="14660" heatid="15651" lane="5" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monika" lastname="Klarecka" birthdate="1977-06-06" gender="F" nation="POL" license="502805600152" swrid="5464091" athleteid="15156">
              <RESULTS>
                <RESULT eventid="1053" points="385" swimtime="00:03:52.51" resultid="15157" heatid="15549" lane="1" entrytime="00:03:50.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.91" />
                    <SPLIT distance="100" swimtime="00:01:52.95" />
                    <SPLIT distance="150" swimtime="00:02:52.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="306" swimtime="00:03:13.54" resultid="15158" heatid="15585" lane="6" entrytime="00:03:16.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.60" />
                    <SPLIT distance="100" swimtime="00:01:33.49" />
                    <SPLIT distance="150" swimtime="00:02:24.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5430" points="250" swimtime="00:04:04.06" resultid="15159" heatid="15615" lane="4" entrytime="00:04:11.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.24" />
                    <SPLIT distance="100" swimtime="00:02:01.95" />
                    <SPLIT distance="150" swimtime="00:03:04.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5404" points="242" swimtime="00:01:45.93" resultid="15160" heatid="15642" lane="5" entrytime="00:01:41.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tadeusz" lastname="Obiedziński" birthdate="1959-05-12" gender="M" nation="POL" license="502805700040" swrid="4992722" athleteid="15173">
              <RESULTS>
                <RESULT eventid="1066" points="283" swimtime="00:04:12.55" resultid="15174" heatid="15554" lane="5" entrytime="00:03:59.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.21" />
                    <SPLIT distance="100" swimtime="00:01:58.72" />
                    <SPLIT distance="150" swimtime="00:03:08.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6830" points="414" swimtime="00:00:43.91" resultid="15175" heatid="15607" lane="6" entrytime="00:00:43.34" entrycourse="SCM" />
                <RESULT eventid="1212" points="357" swimtime="00:01:44.11" resultid="15176" heatid="15627" lane="1" entrytime="00:01:41.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Włodzimierz" lastname="Przytulski" birthdate="1957-01-09" gender="M" nation="POL" license="502805700049" swrid="4754657" athleteid="15254">
              <RESULTS>
                <RESULT eventid="1144" points="690" swimtime="00:00:34.57" resultid="15255" heatid="15580" lane="5" entrytime="00:00:33.46" entrycourse="SCM" />
                <RESULT eventid="5390" points="614" swimtime="00:01:23.20" resultid="15256" heatid="15600" lane="5" />
                <RESULT eventid="1316" points="587" swimtime="00:00:39.79" resultid="15257" heatid="15636" lane="5" entrytime="00:00:39.37" entrycourse="SCM" />
                <RESULT eventid="1238" points="618" swimtime="00:01:11.71" resultid="15258" heatid="15658" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jarosław" lastname="Woźniak" birthdate="1980-09-30" gender="M" nation="POL" license="502805700158" swrid="5506643" athleteid="15177">
              <RESULTS>
                <RESULT eventid="1066" points="268" swimtime="00:03:41.43" resultid="15178" heatid="15556" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.39" />
                    <SPLIT distance="100" swimtime="00:01:41.20" />
                    <SPLIT distance="150" swimtime="00:02:41.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6830" points="404" swimtime="00:00:39.33" resultid="15179" heatid="15607" lane="5" entrytime="00:00:42.18" entrycourse="SCM" />
                <RESULT eventid="1212" points="316" swimtime="00:01:33.28" resultid="15180" heatid="15626" lane="2" entrytime="00:01:36.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="263" swimtime="00:01:19.95" resultid="15181" heatid="15656" lane="1" entrytime="00:01:20.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Wiśniewska" birthdate="1981-02-26" gender="F" nation="POL" license="502805600123" swrid="5464096" athleteid="15161">
              <RESULTS>
                <RESULT eventid="1053" points="226" swimtime="00:04:32.69" resultid="15162" heatid="15550" lane="6" entrytime="00:04:51.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.27" />
                    <SPLIT distance="100" swimtime="00:02:13.42" />
                    <SPLIT distance="150" swimtime="00:03:25.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="159" swimtime="00:00:53.99" resultid="15163" heatid="15577" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="6828" swimtime="00:02:11.50" resultid="15264" heatid="15611" lane="5" entrytime="00:02:07.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                    <SPLIT distance="100" swimtime="00:01:06.24" />
                    <SPLIT distance="150" swimtime="00:01:37.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15254" number="1" />
                    <RELAYPOSITION athleteid="15259" number="2" />
                    <RELAYPOSITION athleteid="15245" number="3" />
                    <RELAYPOSITION athleteid="15196" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1290" swimtime="00:02:05.61" resultid="15269" heatid="15661" lane="5" entrytime="00:02:25.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.79" />
                    <SPLIT distance="100" swimtime="00:01:10.67" />
                    <SPLIT distance="150" swimtime="00:01:38.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15254" number="1" />
                    <RELAYPOSITION athleteid="15192" number="2" />
                    <RELAYPOSITION athleteid="14657" number="3" />
                    <RELAYPOSITION athleteid="15225" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="6828" swimtime="00:02:16.67" resultid="15265" heatid="15612" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                    <SPLIT distance="100" swimtime="00:01:07.04" />
                    <SPLIT distance="150" swimtime="00:01:39.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15201" number="1" />
                    <RELAYPOSITION athleteid="15187" number="2" />
                    <RELAYPOSITION athleteid="15211" number="3" />
                    <RELAYPOSITION athleteid="15240" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1290" swimtime="00:02:34.51" resultid="15270" heatid="15662" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.25" />
                    <SPLIT distance="100" swimtime="00:01:25.75" />
                    <SPLIT distance="150" swimtime="00:01:59.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15201" number="1" />
                    <RELAYPOSITION athleteid="15164" number="2" />
                    <RELAYPOSITION athleteid="15245" number="3" />
                    <RELAYPOSITION athleteid="15196" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="6828" swimtime="00:02:11.25" resultid="15266" heatid="15612" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.50" />
                    <SPLIT distance="100" swimtime="00:01:01.25" />
                    <SPLIT distance="150" swimtime="00:01:45.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15206" number="1" />
                    <RELAYPOSITION athleteid="15192" number="2" />
                    <RELAYPOSITION athleteid="15249" number="3" />
                    <RELAYPOSITION athleteid="15225" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1290" swimtime="00:02:26.68" resultid="15271" heatid="15662" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.08" />
                    <SPLIT distance="100" swimtime="00:01:21.15" />
                    <SPLIT distance="150" swimtime="00:01:55.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15259" number="1" />
                    <RELAYPOSITION athleteid="15187" number="2" />
                    <RELAYPOSITION athleteid="15211" number="3" />
                    <RELAYPOSITION athleteid="15221" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="6828" status="DNS" swimtime="00:00:00.00" resultid="15267" heatid="15612" lane="6" />
                <RESULT eventid="1290" swimtime="00:02:53.11" resultid="15272" heatid="15662" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15206" number="1" />
                    <RELAYPOSITION athleteid="15182" number="2" />
                    <RELAYPOSITION athleteid="15177" number="3" />
                    <RELAYPOSITION athleteid="15156" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="5">
              <RESULTS>
                <RESULT eventid="6828" swimtime="00:02:17.37" resultid="15268" heatid="15612" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                    <SPLIT distance="100" swimtime="00:01:13.27" />
                    <SPLIT distance="150" swimtime="00:01:51.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15182" number="1" />
                    <RELAYPOSITION athleteid="15164" number="2" />
                    <RELAYPOSITION athleteid="14661" number="3" />
                    <RELAYPOSITION athleteid="14657" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1290" swimtime="00:02:47.06" resultid="15273" heatid="15662" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.09" />
                    <SPLIT distance="100" swimtime="00:01:31.72" />
                    <SPLIT distance="150" swimtime="00:02:11.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14661" number="1" />
                    <RELAYPOSITION athleteid="15173" number="2" />
                    <RELAYPOSITION athleteid="15249" number="3" />
                    <RELAYPOSITION athleteid="15240" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="NZ" nation="POL" clubid="14609" name="NZ">
          <ATHLETES>
            <ATHLETE firstname="Dominik" lastname="Rudzki" birthdate="1992-06-21" gender="M" nation="POL" athleteid="15474">
              <RESULTS>
                <RESULT eventid="1092" points="597" swimtime="00:00:26.28" resultid="15475" heatid="15561" lane="5" entrytime="00:00:25.40" />
                <RESULT eventid="5390" points="590" swimtime="00:01:05.55" resultid="15476" heatid="15596" lane="4" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5417" points="583" swimtime="00:01:03.00" resultid="15477" heatid="15643" lane="4" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="606" swimtime="00:00:57.93" resultid="15478" heatid="15651" lane="4" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artur" lastname="Malina" birthdate="1970-02-10" gender="M" nation="POL" athleteid="15450">
              <RESULTS>
                <RESULT eventid="1144" points="119" swimtime="00:00:54.38" resultid="15451" heatid="15581" lane="6" entrytime="00:00:45.00" />
                <RESULT eventid="1066" points="279" swimtime="00:03:56.61" resultid="15452" heatid="15556" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.63" />
                    <SPLIT distance="100" swimtime="00:01:49.63" />
                    <SPLIT distance="150" swimtime="00:02:53.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5417" status="DNS" swimtime="00:00:00.00" resultid="15453" heatid="15644" lane="1" entrytime="00:01:52.00" />
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="15454" heatid="15628" lane="3" entrytime="00:01:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Bądkowski" birthdate="1978-01-01" gender="M" nation="POL" athleteid="14809">
              <RESULTS>
                <RESULT eventid="1092" points="377" swimtime="00:00:33.02" resultid="14810" heatid="15563" lane="1" entrytime="00:00:30.50" />
                <RESULT eventid="1170" points="350" swimtime="00:02:42.77" resultid="14811" heatid="15589" lane="3" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                    <SPLIT distance="100" swimtime="00:01:17.97" />
                    <SPLIT distance="150" swimtime="00:02:00.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" status="DNS" swimtime="00:00:00.00" resultid="14812" heatid="15653" lane="6" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katarzyna" lastname="Koba-Gołaszewska" birthdate="1986-01-01" gender="F" nation="POL" athleteid="14801">
              <RESULTS>
                <RESULT eventid="1079" points="614" swimtime="00:00:30.80" resultid="14802" heatid="15557" lane="5" entrytime="00:00:30.50" />
                <RESULT eventid="1157" points="514" swimtime="00:02:39.91" resultid="14803" heatid="15584" lane="1" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                    <SPLIT distance="100" swimtime="00:01:18.18" />
                    <SPLIT distance="150" swimtime="00:01:59.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="590" swimtime="00:01:08.88" resultid="14804" heatid="15646" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Łukasz" lastname="Szymański" birthdate="1978-01-02" gender="M" nation="POL" athleteid="14610">
              <RESULTS>
                <RESULT eventid="1092" points="483" swimtime="00:00:30.42" resultid="14611" heatid="15563" lane="3" entrytime="00:00:28.76" />
                <RESULT eventid="1238" points="542" swimtime="00:01:04.90" resultid="14612" heatid="15653" lane="2" entrytime="00:01:06.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maciej" lastname="Wilk" birthdate="1991-01-01" gender="M" nation="POL" athleteid="14796">
              <RESULTS>
                <RESULT eventid="1092" points="457" swimtime="00:00:28.73" resultid="14797" heatid="15562" lane="5" entrytime="00:00:28.00" />
                <RESULT eventid="1238" points="445" swimtime="00:01:04.21" resultid="14798" heatid="15660" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="417" swimtime="00:00:30.60" resultid="14799" heatid="15580" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="5417" status="DNS" swimtime="00:00:00.00" resultid="14800" heatid="15643" lane="1" entrytime="00:01:08.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marek" lastname="Wydmuch" birthdate="1962-04-11" gender="M" nation="POL" athleteid="14745">
              <RESULTS>
                <RESULT eventid="1066" points="363" swimtime="00:03:52.47" resultid="14746" heatid="15554" lane="1" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:21.14" />
                    <SPLIT distance="100" swimtime="00:00:54.77" />
                    <SPLIT distance="150" swimtime="00:01:55.21" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Z3/G-8" eventid="5390" status="DSQ" swimtime="00:00:00.00" resultid="14747" heatid="15599" lane="6" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5417" points="238" swimtime="00:01:48.72" resultid="14748" heatid="15644" lane="4" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="369" swimtime="00:01:23.40" resultid="14749" heatid="15654" lane="2" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jacek" lastname="Sokulski" birthdate="1991-01-01" gender="M" nation="POL" swrid="4062177" athleteid="14813">
              <RESULTS>
                <RESULT eventid="1144" points="706" swimtime="00:00:25.68" resultid="14814" heatid="15579" lane="3" entrytime="00:00:24.35" entrycourse="SCM" />
                <RESULT eventid="1170" points="654" swimtime="00:02:02.67" resultid="14815" heatid="15588" lane="3" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.63" />
                    <SPLIT distance="100" swimtime="00:01:01.61" />
                    <SPLIT distance="150" swimtime="00:01:34.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5417" points="643" swimtime="00:01:00.96" resultid="14816" heatid="15643" lane="3" entrytime="00:00:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="801" swimtime="00:00:52.79" resultid="14817" heatid="15658" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Grzegorz" lastname="Paszkiewicz" birthdate="1975-01-01" gender="M" nation="POL" athleteid="14805">
              <RESULTS>
                <RESULT eventid="1092" points="305" swimtime="00:00:35.46" resultid="14806" heatid="15565" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1238" points="276" swimtime="00:01:21.22" resultid="14807" heatid="15655" lane="3" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="252" swimtime="00:00:40.65" resultid="14808" heatid="15581" lane="5" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michał" lastname="Szymaniak" birthdate="1993-09-06" gender="M" nation="POL" athleteid="14614">
              <RESULTS>
                <RESULT eventid="1092" points="302" swimtime="00:00:32.98" resultid="14615" heatid="15565" lane="3" entrytime="00:00:33.55" />
                <RESULT eventid="1144" points="213" swimtime="00:00:38.28" resultid="14616" heatid="15581" lane="4" entrytime="00:00:37.89" />
                <RESULT eventid="1238" status="DNS" swimtime="00:00:00.00" resultid="14617" heatid="15655" lane="2" entrytime="00:01:15.82" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rajmund" lastname="Grys" birthdate="1977-01-01" gender="M" nation="POL" athleteid="14818">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="14819" heatid="15566" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="1170" status="DNS" swimtime="00:00:00.00" resultid="14820" heatid="15590" lane="3" entrytime="00:03:00.00" />
                <RESULT eventid="1238" status="DNS" swimtime="00:00:00.00" resultid="14821" heatid="15656" lane="5" entrytime="00:01:20.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="RAAS" nation="POL" clubid="14576" name="Rydułtowska Akademia Aktyw. Seniora">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Lippa" birthdate="1946-02-02" gender="F" nation="POL" swrid="5484413" athleteid="14582">
              <RESULTS>
                <RESULT eventid="1053" points="99" swimtime="00:07:46.25" resultid="14583" heatid="15551" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:44.09" />
                    <SPLIT distance="100" swimtime="00:03:44.77" />
                    <SPLIT distance="150" swimtime="00:05:46.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="71" swimtime="00:07:14.11" resultid="14584" heatid="15587" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:36.77" />
                    <SPLIT distance="100" swimtime="00:03:30.12" />
                    <SPLIT distance="150" swimtime="00:05:25.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="74" swimtime="00:01:43.55" resultid="14585" heatid="15634" lane="3" entrytime="00:01:38.15" entrycourse="SCM" />
                <RESULT eventid="1225" points="46" swimtime="00:03:40.22" resultid="14586" heatid="15649" lane="5" entrytime="00:03:09.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:37.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rudolf" lastname="Bugla" birthdate="1940-05-16" gender="M" nation="POL" swrid="4831499" athleteid="14592">
              <RESULTS>
                <RESULT eventid="1066" points="196" swimtime="00:06:13.67" resultid="14593" heatid="15555" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.98" />
                    <SPLIT distance="100" swimtime="00:02:59.24" />
                    <SPLIT distance="150" swimtime="00:04:38.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6830" points="141" swimtime="00:01:22.46" resultid="14594" heatid="15609" lane="2" entrytime="00:01:05.90" entrycourse="SCM" />
                <RESULT eventid="1212" points="154" swimtime="00:03:00.72" resultid="14595" heatid="15628" lane="5" entrytime="00:02:45.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="76" swimtime="00:02:53.42" resultid="14596" heatid="15659" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernard" lastname="Poloczek" birthdate="1947-02-25" gender="M" nation="POL" swrid="4792004" athleteid="14587">
              <RESULTS>
                <RESULT eventid="1118" points="494" swimtime="00:01:43.23" resultid="14588" heatid="15573" lane="5" entrytime="00:01:45.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="397" swimtime="00:00:46.23" resultid="14589" heatid="15582" lane="3" entrytime="00:00:45.23" entrycourse="SCM" />
                <RESULT eventid="1316" points="520" swimtime="00:00:45.25" resultid="14590" heatid="15638" lane="2" entrytime="00:00:46.57" entrycourse="SCM" />
                <RESULT eventid="1238" points="397" swimtime="00:01:36.75" resultid="14591" heatid="15659" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jerzy" lastname="Ciecior" birthdate="1953-11-24" gender="M" nation="POL" swrid="4934027" athleteid="14577">
              <RESULTS>
                <RESULT eventid="1118" points="442" swimtime="00:01:38.56" resultid="14578" heatid="15573" lane="3" entrytime="00:01:37.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="444" swimtime="00:03:13.91" resultid="14579" heatid="15592" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.45" />
                    <SPLIT distance="100" swimtime="00:01:33.83" />
                    <SPLIT distance="150" swimtime="00:02:25.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="598" swimtime="00:00:41.15" resultid="14580" heatid="15637" lane="2" entrytime="00:00:40.65" entrycourse="SCM" />
                <RESULT eventid="1238" points="493" swimtime="00:01:21.75" resultid="14581" heatid="15660" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>

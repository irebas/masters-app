<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Miejski Klub Plywacki" version="11.37565">
    <CONTACT name="Swimrankings" street="Weltpoststrasse 5" city="Bern" zip="3015" country="CH" phone="+41 99 999 99 99" fax="+41 99 999 99 99" email="sales@swimrankings.net" internet="http://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Szczecin" name="Otwarte Mistrzostwa Polski w Pływaniu Masters" course="LCM" deadline="2015-06-05" nation="POL" timing="AUTOMATIC">
      <AGEDATE value="2015-06-28" type="YEAR" />
      <POOL lanemax="9" />
      <POINTTABLE pointtableid="1121" name="DSV Master Performance Table" version="2013" />
      <SESSIONS>
        <SESSION date="2015-06-26" daytime="15:00" name="I Blok" number="1" warmupfrom="14:00">
          <EVENTS>
            <EVENT eventid="1090" daytime="16:09" gender="F" number="3" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2259" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5264" />
                    <RANKING order="2" place="2" resultid="4667" />
                    <RANKING order="3" place="3" resultid="2847" />
                    <RANKING order="4" place="4" resultid="4614" />
                    <RANKING order="5" place="5" resultid="4055" />
                    <RANKING order="6" place="-1" resultid="3590" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2260" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5411" />
                    <RANKING order="2" place="2" resultid="5036" />
                    <RANKING order="3" place="3" resultid="3762" />
                    <RANKING order="4" place="4" resultid="5208" />
                    <RANKING order="5" place="5" resultid="3984" />
                    <RANKING order="6" place="6" resultid="4326" />
                    <RANKING order="7" place="7" resultid="4660" />
                    <RANKING order="8" place="8" resultid="3103" />
                    <RANKING order="9" place="9" resultid="3978" />
                    <RANKING order="10" place="10" resultid="4597" />
                    <RANKING order="11" place="11" resultid="4632" />
                    <RANKING order="12" place="12" resultid="3056" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2261" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3966" />
                    <RANKING order="2" place="2" resultid="3470" />
                    <RANKING order="3" place="3" resultid="3973" />
                    <RANKING order="4" place="4" resultid="4820" />
                    <RANKING order="5" place="5" resultid="2941" />
                    <RANKING order="6" place="6" resultid="3886" />
                    <RANKING order="7" place="-1" resultid="4586" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2262" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3117" />
                    <RANKING order="2" place="2" resultid="4907" />
                    <RANKING order="3" place="3" resultid="2130" />
                    <RANKING order="4" place="4" resultid="4878" />
                    <RANKING order="5" place="5" resultid="5196" />
                    <RANKING order="6" place="6" resultid="4776" />
                    <RANKING order="7" place="-1" resultid="5406" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2263" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4995" />
                    <RANKING order="2" place="2" resultid="5399" />
                    <RANKING order="3" place="3" resultid="2946" />
                    <RANKING order="4" place="4" resultid="3945" />
                    <RANKING order="5" place="5" resultid="3740" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2264" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3873" />
                    <RANKING order="2" place="2" resultid="5170" />
                    <RANKING order="3" place="3" resultid="4262" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2265" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5064" />
                    <RANKING order="2" place="2" resultid="5008" />
                    <RANKING order="3" place="3" resultid="3286" />
                    <RANKING order="4" place="4" resultid="3669" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2266" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5372" />
                    <RANKING order="2" place="2" resultid="5278" />
                    <RANKING order="3" place="3" resultid="3881" />
                    <RANKING order="4" place="4" resultid="4496" />
                    <RANKING order="5" place="5" resultid="5753" />
                    <RANKING order="6" place="6" resultid="3048" />
                    <RANKING order="7" place="7" resultid="3745" />
                    <RANKING order="8" place="8" resultid="3446" />
                    <RANKING order="9" place="9" resultid="5283" />
                    <RANKING order="10" place="10" resultid="4445" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2267" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5364" />
                    <RANKING order="2" place="2" resultid="3432" />
                    <RANKING order="3" place="3" resultid="3622" />
                    <RANKING order="4" place="4" resultid="3415" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2268" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5270" />
                    <RANKING order="2" place="2" resultid="3909" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2269" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="2270" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4954" />
                    <RANKING order="2" place="2" resultid="4008" />
                    <RANKING order="3" place="3" resultid="2226" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2271" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="2272" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2273" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7954" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7955" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7956" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7957" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7958" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7959" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7960" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1075" daytime="15:21" gender="M" number="2" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2244" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3704" />
                    <RANKING order="2" place="2" resultid="4581" />
                    <RANKING order="3" place="3" resultid="4205" />
                    <RANKING order="4" place="4" resultid="3143" />
                    <RANKING order="5" place="5" resultid="4307" />
                    <RANKING order="6" place="6" resultid="3713" />
                    <RANKING order="7" place="-1" resultid="3581" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2245" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5042" />
                    <RANKING order="2" place="2" resultid="4647" />
                    <RANKING order="3" place="3" resultid="5027" />
                    <RANKING order="4" place="4" resultid="3338" />
                    <RANKING order="5" place="5" resultid="3604" />
                    <RANKING order="6" place="-1" resultid="2880" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2246" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4638" />
                    <RANKING order="2" place="2" resultid="4294" />
                    <RANKING order="3" place="3" resultid="2789" />
                    <RANKING order="4" place="4" resultid="4281" />
                    <RANKING order="5" place="5" resultid="4142" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2247" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4827" />
                    <RANKING order="2" place="2" resultid="3655" />
                    <RANKING order="3" place="3" resultid="5047" />
                    <RANKING order="4" place="4" resultid="3123" />
                    <RANKING order="5" place="5" resultid="4164" />
                    <RANKING order="6" place="6" resultid="2817" />
                    <RANKING order="7" place="7" resultid="3775" />
                    <RANKING order="8" place="8" resultid="4792" />
                    <RANKING order="9" place="9" resultid="4158" />
                    <RANKING order="10" place="10" resultid="3064" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2248" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4230" />
                    <RANKING order="2" place="2" resultid="3135" />
                    <RANKING order="3" place="3" resultid="4717" />
                    <RANKING order="4" place="4" resultid="4913" />
                    <RANKING order="5" place="5" resultid="3956" />
                    <RANKING order="6" place="6" resultid="3863" />
                    <RANKING order="7" place="7" resultid="4246" />
                    <RANKING order="8" place="8" resultid="4050" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2249" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4524" />
                    <RANKING order="2" place="2" resultid="4516" />
                    <RANKING order="3" place="3" resultid="2810" />
                    <RANKING order="4" place="4" resultid="3841" />
                    <RANKING order="5" place="5" resultid="5163" />
                    <RANKING order="6" place="6" resultid="4036" />
                    <RANKING order="7" place="7" resultid="4416" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2250" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5477" />
                    <RANKING order="2" place="2" resultid="3780" />
                    <RANKING order="3" place="3" resultid="4709" />
                    <RANKING order="4" place="4" resultid="3939" />
                    <RANKING order="5" place="5" resultid="3680" />
                    <RANKING order="6" place="6" resultid="4723" />
                    <RANKING order="7" place="7" resultid="3153" />
                    <RANKING order="8" place="8" resultid="2833" />
                    <RANKING order="9" place="-1" resultid="5429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2251" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3084" />
                    <RANKING order="2" place="2" resultid="4255" />
                    <RANKING order="3" place="3" resultid="5055" />
                    <RANKING order="4" place="4" resultid="5300" />
                    <RANKING order="5" place="5" resultid="2155" />
                    <RANKING order="6" place="6" resultid="5031" />
                    <RANKING order="7" place="7" resultid="2164" />
                    <RANKING order="8" place="8" resultid="2171" />
                    <RANKING order="9" place="-1" resultid="4187" />
                    <RANKING order="10" place="-1" resultid="4555" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2252" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2964" />
                    <RANKING order="2" place="2" resultid="3496" />
                    <RANKING order="3" place="3" resultid="5292" />
                    <RANKING order="4" place="4" resultid="3003" />
                    <RANKING order="5" place="5" resultid="4408" />
                    <RANKING order="6" place="6" resultid="4806" />
                    <RANKING order="7" place="7" resultid="3568" />
                    <RANKING order="8" place="8" resultid="3751" />
                    <RANKING order="9" place="9" resultid="3271" />
                    <RANKING order="10" place="10" resultid="4762" />
                    <RANKING order="11" place="11" resultid="3518" />
                    <RANKING order="12" place="12" resultid="4399" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2253" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4239" />
                    <RANKING order="2" place="2" resultid="3789" />
                    <RANKING order="3" place="3" resultid="5022" />
                    <RANKING order="4" place="4" resultid="3899" />
                    <RANKING order="5" place="5" resultid="3406" />
                    <RANKING order="6" place="6" resultid="4969" />
                    <RANKING order="7" place="7" resultid="3645" />
                    <RANKING order="8" place="8" resultid="4366" />
                    <RANKING order="9" place="-1" resultid="3637" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2254" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2116" />
                    <RANKING order="2" place="2" resultid="2106" />
                    <RANKING order="3" place="3" resultid="3891" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2255" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3422" />
                    <RANKING order="2" place="2" resultid="4425" />
                    <RANKING order="3" place="3" resultid="2769" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2256" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="2257" agemax="89" agemin="85" name="Kat. M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4084" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2258" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7945" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7946" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7947" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7948" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7949" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7950" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7951" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7952" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7953" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1120" daytime="16:45" gender="F" number="5" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2289" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4620" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2290" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2957" />
                    <RANKING order="2" place="2" resultid="5087" />
                    <RANKING order="3" place="-1" resultid="4768" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2291" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3098" />
                    <RANKING order="2" place="2" resultid="3507" />
                    <RANKING order="3" place="3" resultid="3091" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2292" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4869" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2293" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5139" />
                    <RANKING order="2" place="2" resultid="5400" />
                    <RANKING order="3" place="3" resultid="3946" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2294" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3021" />
                    <RANKING order="2" place="2" resultid="4864" />
                    <RANKING order="3" place="3" resultid="3042" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2295" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3287" />
                    <RANKING order="2" place="2" resultid="3396" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2296" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4547" />
                    <RANKING order="2" place="2" resultid="4497" />
                    <RANKING order="3" place="3" resultid="4454" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2297" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3623" />
                    <RANKING order="2" place="2" resultid="5101" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2298" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2888" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2299" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="2300" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4955" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2301" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="2302" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2303" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8136" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8137" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8138" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1165" daytime="19:00" gender="M" number="8" order="8" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2334" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4308" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2335" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3008" />
                    <RANKING order="2" place="2" resultid="4182" />
                    <RANKING order="3" place="3" resultid="3303" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2336" agemax="34" agemin="30" name="Kat. B" />
                <AGEGROUP agegroupid="2337" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3656" />
                    <RANKING order="2" place="2" resultid="2818" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2338" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4887" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2339" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5453" />
                    <RANKING order="2" place="2" resultid="3716" />
                    <RANKING order="3" place="3" resultid="3842" />
                    <RANKING order="4" place="4" resultid="4940" />
                    <RANKING order="5" place="5" resultid="5164" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2340" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4334" />
                    <RANKING order="2" place="2" resultid="4724" />
                    <RANKING order="3" place="3" resultid="5152" />
                    <RANKING order="4" place="4" resultid="3809" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2341" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4692" />
                    <RANKING order="2" place="2" resultid="3728" />
                    <RANKING order="3" place="3" resultid="4556" />
                    <RANKING order="4" place="4" resultid="5423" />
                    <RANKING order="5" place="5" resultid="3734" />
                    <RANKING order="6" place="6" resultid="3203" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2342" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3497" />
                    <RANKING order="2" place="2" resultid="4409" />
                    <RANKING order="3" place="3" resultid="5322" />
                    <RANKING order="4" place="4" resultid="3853" />
                    <RANKING order="5" place="5" resultid="3211" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2343" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3790" />
                    <RANKING order="2" place="2" resultid="6438" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2344" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2117" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2345" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2099" />
                    <RANKING order="2" place="2" resultid="3927" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2346" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3178" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2347" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2348" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8143" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8144" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8145" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8146" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1150" daytime="18:27" gender="F" number="7" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2319" agemax="24" agemin="20" name="Kat. 0" />
                <AGEGROUP agegroupid="2320" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3057" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2321" agemax="34" agemin="30" name="Kat. B" />
                <AGEGROUP agegroupid="2322" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5758" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2323" agemax="44" agemin="40" name="Kat. D" />
                <AGEGROUP agegroupid="2324" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3109" />
                    <RANKING order="2" place="2" resultid="4699" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2325" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3691" />
                    <RANKING order="2" place="2" resultid="4563" />
                    <RANKING order="3" place="3" resultid="5093" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2326" agemax="59" agemin="55" name="Kat. G" />
                <AGEGROUP agegroupid="2327" agemax="64" agemin="60" name="Kat. H" />
                <AGEGROUP agegroupid="2328" agemax="69" agemin="65" name="Kat. I" />
                <AGEGROUP agegroupid="2329" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5134" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2330" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="2331" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="2332" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2333" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8142" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1135" daytime="17:38" gender="M" number="6" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2304" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4436" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2305" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3001" />
                    <RANKING order="2" place="2" resultid="5244" />
                    <RANKING order="3" place="3" resultid="3356" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2306" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2790" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2307" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4503" />
                    <RANKING order="2" place="2" resultid="2905" />
                    <RANKING order="3" place="3" resultid="4132" />
                    <RANKING order="4" place="4" resultid="3065" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2308" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3013" />
                    <RANKING order="2" place="2" resultid="4921" />
                    <RANKING order="3" place="3" resultid="3957" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2309" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4061" />
                    <RANKING order="2" place="2" resultid="5440" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2310" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5434" />
                    <RANKING order="2" place="2" resultid="3685" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2311" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2156" />
                    <RANKING order="2" place="2" resultid="2912" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2312" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3519" />
                    <RANKING order="2" place="2" resultid="3272" />
                    <RANKING order="3" place="3" resultid="5288" />
                    <RANKING order="4" place="4" resultid="4400" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2313" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3900" />
                    <RANKING order="2" place="2" resultid="4970" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2314" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="2315" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="2316" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4015" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2317" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2318" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8139" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8140" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8141" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1058" daytime="15:00" gender="F" number="1" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1062" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4613" />
                    <RANKING order="2" place="2" resultid="3597" />
                    <RANKING order="3" place="-1" resultid="3589" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1063" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2783" />
                    <RANKING order="2" place="2" resultid="4325" />
                    <RANKING order="3" place="3" resultid="3983" />
                    <RANKING order="4" place="4" resultid="4531" />
                    <RANKING order="5" place="5" resultid="4631" />
                    <RANKING order="6" place="6" resultid="3102" />
                    <RANKING order="7" place="-1" resultid="4607" />
                    <RANKING order="8" place="-1" resultid="4767" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1064" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4819" />
                    <RANKING order="2" place="2" resultid="4073" />
                    <RANKING order="3" place="3" resultid="5205" />
                    <RANKING order="4" place="4" resultid="3506" />
                    <RANKING order="5" place="5" resultid="4538" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3116" />
                    <RANKING order="2" place="2" resultid="4877" />
                    <RANKING order="3" place="3" resultid="2129" />
                    <RANKING order="4" place="4" resultid="4775" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5000" />
                    <RANKING order="2" place="2" resultid="3739" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4261" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1068" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5388" />
                    <RANKING order="2" place="2" resultid="5007" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4546" />
                    <RANKING order="2" place="2" resultid="5371" />
                    <RANKING order="3" place="3" resultid="3047" />
                    <RANKING order="4" place="4" resultid="4453" />
                    <RANKING order="5" place="5" resultid="3445" />
                    <RANKING order="6" place="6" resultid="3744" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5359" />
                    <RANKING order="2" place="2" resultid="3431" />
                    <RANKING order="3" place="3" resultid="3414" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3908" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1072" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="1073" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="1074" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="2243" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="1059" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7941" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7942" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7943" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7944" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1105" daytime="16:24" gender="M" number="4" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2274" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3770" />
                    <RANKING order="2" place="2" resultid="4385" />
                    <RANKING order="3" place="3" resultid="4320" />
                    <RANKING order="4" place="4" resultid="4206" />
                    <RANKING order="5" place="5" resultid="3705" />
                    <RANKING order="6" place="6" resultid="3714" />
                    <RANKING order="7" place="7" resultid="4435" />
                    <RANKING order="8" place="-1" resultid="3582" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2275" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2881" />
                    <RANKING order="2" place="2" resultid="4270" />
                    <RANKING order="3" place="3" resultid="4218" />
                    <RANKING order="4" place="4" resultid="4222" />
                    <RANKING order="5" place="5" resultid="4079" />
                    <RANKING order="6" place="6" resultid="4648" />
                    <RANKING order="7" place="7" resultid="5252" />
                    <RANKING order="8" place="8" resultid="3355" />
                    <RANKING order="9" place="9" resultid="3350" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2276" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2137" />
                    <RANKING order="2" place="2" resultid="4295" />
                    <RANKING order="3" place="3" resultid="5258" />
                    <RANKING order="4" place="4" resultid="4639" />
                    <RANKING order="5" place="5" resultid="4288" />
                    <RANKING order="6" place="6" resultid="5223" />
                    <RANKING order="7" place="7" resultid="3148" />
                    <RANKING order="8" place="-1" resultid="4592" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2277" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4828" />
                    <RANKING order="2" place="2" resultid="3464" />
                    <RANKING order="3" place="3" resultid="5048" />
                    <RANKING order="4" place="4" resultid="3169" />
                    <RANKING order="5" place="5" resultid="4578" />
                    <RANKING order="6" place="6" resultid="4165" />
                    <RANKING order="7" place="7" resultid="5313" />
                    <RANKING order="8" place="8" resultid="4755" />
                    <RANKING order="9" place="9" resultid="2904" />
                    <RANKING order="10" place="10" resultid="4793" />
                    <RANKING order="11" place="11" resultid="2864" />
                    <RANKING order="12" place="12" resultid="5215" />
                    <RANKING order="13" place="13" resultid="4177" />
                    <RANKING order="14" place="14" resultid="3364" />
                    <RANKING order="15" place="15" resultid="2970" />
                    <RANKING order="16" place="16" resultid="4100" />
                    <RANKING order="17" place="-1" resultid="4131" />
                    <RANKING order="18" place="-1" resultid="4137" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2278" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4231" />
                    <RANKING order="2" place="2" resultid="3136" />
                    <RANKING order="3" place="3" resultid="2213" />
                    <RANKING order="4" place="4" resultid="5187" />
                    <RANKING order="5" place="4" resultid="5219" />
                    <RANKING order="6" place="6" resultid="3297" />
                    <RANKING order="7" place="7" resultid="4920" />
                    <RANKING order="8" place="8" resultid="4212" />
                    <RANKING order="9" place="9" resultid="4914" />
                    <RANKING order="10" place="10" resultid="4394" />
                    <RANKING order="11" place="11" resultid="3129" />
                    <RANKING order="12" place="12" resultid="4894" />
                    <RANKING order="13" place="13" resultid="4381" />
                    <RANKING order="14" place="14" resultid="4743" />
                    <RANKING order="15" place="15" resultid="4247" />
                    <RANKING order="16" place="16" resultid="3370" />
                    <RANKING order="17" place="17" resultid="4886" />
                    <RANKING order="18" place="18" resultid="4654" />
                    <RANKING order="19" place="19" resultid="4470" />
                    <RANKING order="20" place="-1" resultid="3801" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2279" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2778" />
                    <RANKING order="2" place="2" resultid="2952" />
                    <RANKING order="3" place="3" resultid="2741" />
                    <RANKING order="4" place="4" resultid="5183" />
                    <RANKING order="5" place="5" resultid="3281" />
                    <RANKING order="6" place="6" resultid="5158" />
                    <RANKING order="7" place="7" resultid="2811" />
                    <RANKING order="8" place="8" resultid="4939" />
                    <RANKING order="9" place="9" resultid="4417" />
                    <RANKING order="10" place="10" resultid="2854" />
                    <RANKING order="11" place="-1" resultid="4900" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2280" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5081" />
                    <RANKING order="2" place="2" resultid="3698" />
                    <RANKING order="3" place="3" resultid="5478" />
                    <RANKING order="4" place="4" resultid="3781" />
                    <RANKING order="5" place="5" resultid="3940" />
                    <RANKING order="6" place="6" resultid="2834" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2281" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3085" />
                    <RANKING order="2" place="2" resultid="4490" />
                    <RANKING order="3" place="3" resultid="5056" />
                    <RANKING order="4" place="4" resultid="4948" />
                    <RANKING order="5" place="5" resultid="2754" />
                    <RANKING order="6" place="6" resultid="5764" />
                    <RANKING order="7" place="7" resultid="4691" />
                    <RANKING order="8" place="8" resultid="5301" />
                    <RANKING order="9" place="9" resultid="3202" />
                    <RANKING order="10" place="10" resultid="5416" />
                    <RANKING order="11" place="11" resultid="3727" />
                    <RANKING order="12" place="12" resultid="6025" />
                    <RANKING order="13" place="-1" resultid="4963" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2282" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4476" />
                    <RANKING order="2" place="2" resultid="4807" />
                    <RANKING order="3" place="3" resultid="3752" />
                    <RANKING order="4" place="4" resultid="4813" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2283" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5115" />
                    <RANKING order="2" place="2" resultid="5015" />
                    <RANKING order="3" place="3" resultid="2797" />
                    <RANKING order="4" place="4" resultid="3386" />
                    <RANKING order="5" place="5" resultid="4367" />
                    <RANKING order="6" place="6" resultid="5110" />
                    <RANKING order="7" place="7" resultid="6018" />
                    <RANKING order="8" place="8" resultid="3646" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2284" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2107" />
                    <RANKING order="2" place="2" resultid="2183" />
                    <RANKING order="3" place="3" resultid="3892" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2285" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3423" />
                    <RANKING order="2" place="2" resultid="4426" />
                    <RANKING order="3" place="3" resultid="2770" />
                    <RANKING order="4" place="4" resultid="4023" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2286" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="2287" agemax="89" agemin="85" name="Kat. M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4085" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2288" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7961" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7962" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7963" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7964" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7965" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7966" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7967" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7968" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7969" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7970" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7971" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7972" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2015-06-27" daytime="09:00" name="II Blok" number="2" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="1228" daytime="10:06" gender="M" number="12" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2394" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4582" />
                    <RANKING order="2" place="2" resultid="3144" />
                    <RANKING order="3" place="3" resultid="3771" />
                    <RANKING order="4" place="-1" resultid="3194" />
                    <RANKING order="5" place="-1" resultid="3584" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2395" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3546" />
                    <RANKING order="2" place="2" resultid="2873" />
                    <RANKING order="3" place="3" resultid="3073" />
                    <RANKING order="4" place="4" resultid="5340" />
                    <RANKING order="5" place="5" resultid="5043" />
                    <RANKING order="6" place="6" resultid="5246" />
                    <RANKING order="7" place="7" resultid="3358" />
                    <RANKING order="8" place="8" resultid="4272" />
                    <RANKING order="9" place="9" resultid="5254" />
                    <RANKING order="10" place="10" resultid="5028" />
                    <RANKING order="11" place="11" resultid="3605" />
                    <RANKING order="12" place="12" resultid="3340" />
                    <RANKING order="13" place="-1" resultid="2895" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2396" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5259" />
                    <RANKING order="2" place="2" resultid="2842" />
                    <RANKING order="3" place="3" resultid="4296" />
                    <RANKING order="4" place="4" resultid="2791" />
                    <RANKING order="5" place="5" resultid="4283" />
                    <RANKING order="6" place="6" resultid="5224" />
                    <RANKING order="7" place="7" resultid="4290" />
                    <RANKING order="8" place="-1" resultid="4143" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2397" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4830" />
                    <RANKING order="2" place="2" resultid="5050" />
                    <RANKING order="3" place="3" resultid="3170" />
                    <RANKING order="4" place="4" resultid="5315" />
                    <RANKING order="5" place="5" resultid="3776" />
                    <RANKING order="6" place="6" resultid="4167" />
                    <RANKING order="7" place="7" resultid="4159" />
                    <RANKING order="8" place="8" resultid="3918" />
                    <RANKING order="9" place="9" resultid="4102" />
                    <RANKING order="10" place="-1" resultid="4149" />
                    <RANKING order="11" place="-1" resultid="4154" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2398" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6411" />
                    <RANKING order="2" place="2" resultid="2214" />
                    <RANKING order="3" place="3" resultid="5347" />
                    <RANKING order="4" place="4" resultid="4923" />
                    <RANKING order="5" place="5" resultid="4915" />
                    <RANKING order="6" place="6" resultid="3958" />
                    <RANKING order="7" place="7" resultid="2802" />
                    <RANKING order="8" place="8" resultid="5220" />
                    <RANKING order="9" place="9" resultid="5188" />
                    <RANKING order="10" place="10" resultid="4895" />
                    <RANKING order="11" place="11" resultid="2151" />
                    <RANKING order="12" place="12" resultid="4051" />
                    <RANKING order="13" place="13" resultid="3077" />
                    <RANKING order="14" place="14" resultid="3308" />
                    <RANKING order="15" place="15" resultid="3390" />
                    <RANKING order="16" place="16" resultid="3372" />
                    <RANKING order="17" place="17" resultid="3803" />
                    <RANKING order="18" place="18" resultid="4029" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2399" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2742" />
                    <RANKING order="2" place="2" resultid="4063" />
                    <RANKING order="3" place="3" resultid="5442" />
                    <RANKING order="4" place="4" resultid="4902" />
                    <RANKING order="5" place="5" resultid="3630" />
                    <RANKING order="6" place="6" resultid="4419" />
                    <RANKING order="7" place="7" resultid="3613" />
                    <RANKING order="8" place="-1" resultid="5309" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2400" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3941" />
                    <RANKING order="2" place="2" resultid="4710" />
                    <RANKING order="3" place="3" resultid="3783" />
                    <RANKING order="4" place="4" resultid="3681" />
                    <RANKING order="5" place="5" resultid="5082" />
                    <RANKING order="6" place="6" resultid="5430" />
                    <RANKING order="7" place="7" resultid="5153" />
                    <RANKING order="8" place="8" resultid="3575" />
                    <RANKING order="9" place="9" resultid="5746" />
                    <RANKING order="10" place="10" resultid="3811" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2401" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6033" />
                    <RANKING order="2" place="2" resultid="2765" />
                    <RANKING order="3" place="3" resultid="4949" />
                    <RANKING order="4" place="4" resultid="5032" />
                    <RANKING order="5" place="5" resultid="5417" />
                    <RANKING order="6" place="6" resultid="4856" />
                    <RANKING order="7" place="7" resultid="2755" />
                    <RANKING order="8" place="8" resultid="5303" />
                    <RANKING order="9" place="9" resultid="3205" />
                    <RANKING order="10" place="10" resultid="2172" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2402" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3569" />
                    <RANKING order="2" place="2" resultid="3004" />
                    <RANKING order="3" place="3" resultid="3402" />
                    <RANKING order="4" place="3" resultid="5293" />
                    <RANKING order="5" place="5" resultid="3753" />
                    <RANKING order="6" place="6" resultid="4737" />
                    <RANKING order="7" place="7" resultid="3485" />
                    <RANKING order="8" place="8" resultid="4401" />
                    <RANKING order="9" place="9" resultid="4814" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2403" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4991" />
                    <RANKING order="2" place="2" resultid="5023" />
                    <RANKING order="3" place="3" resultid="3407" />
                    <RANKING order="4" place="4" resultid="3647" />
                    <RANKING order="5" place="5" resultid="6020" />
                    <RANKING order="6" place="-1" resultid="3639" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2404" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2109" />
                    <RANKING order="2" place="2" resultid="2184" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2405" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3424" />
                    <RANKING order="2" place="2" resultid="5125" />
                    <RANKING order="3" place="3" resultid="4427" />
                    <RANKING order="4" place="4" resultid="2771" />
                    <RANKING order="5" place="5" resultid="3929" />
                    <RANKING order="6" place="6" resultid="4024" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2406" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3381" />
                    <RANKING order="2" place="2" resultid="3180" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2407" agemax="89" agemin="85" name="Kat. M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4087" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2408" agemax="94" agemin="90" name="Kat. N">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5077" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8000" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8001" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8002" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8003" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8004" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8005" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8006" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="8007" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="8008" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="8009" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="8010" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1181" daytime="09:00" gender="F" number="9" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2349" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4108" />
                    <RANKING order="2" place="2" resultid="5265" />
                    <RANKING order="3" place="3" resultid="2848" />
                    <RANKING order="4" place="4" resultid="3550" />
                    <RANKING order="5" place="5" resultid="4615" />
                    <RANKING order="6" place="-1" resultid="3591" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2350" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5412" />
                    <RANKING order="2" place="2" resultid="3763" />
                    <RANKING order="3" place="3" resultid="5037" />
                    <RANKING order="4" place="4" resultid="2930" />
                    <RANKING order="5" place="5" resultid="4661" />
                    <RANKING order="6" place="6" resultid="5209" />
                    <RANKING order="7" place="7" resultid="4532" />
                    <RANKING order="8" place="8" resultid="4598" />
                    <RANKING order="9" place="9" resultid="5237" />
                    <RANKING order="10" place="10" resultid="2901" />
                    <RANKING order="11" place="11" resultid="3058" />
                    <RANKING order="12" place="12" resultid="5088" />
                    <RANKING order="13" place="13" resultid="2936" />
                    <RANKING order="14" place="-1" resultid="4327" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2351" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2869" />
                    <RANKING order="2" place="2" resultid="3967" />
                    <RANKING order="3" place="3" resultid="4587" />
                    <RANKING order="4" place="4" resultid="3092" />
                    <RANKING order="5" place="5" resultid="4539" />
                    <RANKING order="6" place="6" resultid="3508" />
                    <RANKING order="7" place="7" resultid="2942" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2352" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5759" />
                    <RANKING order="2" place="2" resultid="4908" />
                    <RANKING order="3" place="3" resultid="4879" />
                    <RANKING order="4" place="4" resultid="5197" />
                    <RANKING order="5" place="5" resultid="4777" />
                    <RANKING order="6" place="6" resultid="4093" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2353" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5140" />
                    <RANKING order="2" place="2" resultid="5401" />
                    <RANKING order="3" place="3" resultid="3947" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2354" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3874" />
                    <RANKING order="2" place="2" resultid="3110" />
                    <RANKING order="3" place="3" resultid="5176" />
                    <RANKING order="4" place="4" resultid="4678" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2355" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5065" />
                    <RANKING order="2" place="2" resultid="5009" />
                    <RANKING order="3" place="3" resultid="5378" />
                    <RANKING order="4" place="4" resultid="3288" />
                    <RANKING order="5" place="5" resultid="3692" />
                    <RANKING order="6" place="6" resultid="5094" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2356" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5373" />
                    <RANKING order="2" place="2" resultid="3882" />
                    <RANKING order="3" place="3" resultid="4498" />
                    <RANKING order="4" place="4" resultid="4548" />
                    <RANKING order="5" place="5" resultid="3746" />
                    <RANKING order="6" place="6" resultid="3049" />
                    <RANKING order="7" place="7" resultid="5754" />
                    <RANKING order="8" place="8" resultid="5284" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2357" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5365" />
                    <RANKING order="2" place="2" resultid="3433" />
                    <RANKING order="3" place="3" resultid="3624" />
                    <RANKING order="4" place="4" resultid="5102" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2358" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5271" />
                    <RANKING order="2" place="2" resultid="5146" />
                    <RANKING order="3" place="3" resultid="2805" />
                    <RANKING order="4" place="4" resultid="2889" />
                    <RANKING order="5" place="5" resultid="3910" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2359" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3440" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2360" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4956" />
                    <RANKING order="2" place="2" resultid="5354" />
                    <RANKING order="3" place="3" resultid="4001" />
                    <RANKING order="4" place="4" resultid="4009" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2361" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="2362" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2363" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7973" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7974" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7975" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7976" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7977" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7978" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7979" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1258" daytime="10:40" gender="M" number="14" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2424" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3707" />
                    <RANKING order="2" place="2" resultid="4321" />
                    <RANKING order="3" place="3" resultid="4309" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2425" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4183" />
                    <RANKING order="2" place="2" resultid="4649" />
                    <RANKING order="3" place="3" resultid="3009" />
                    <RANKING order="4" place="-1" resultid="4627" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2426" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4297" />
                    <RANKING order="2" place="2" resultid="4786" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2427" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3657" />
                    <RANKING order="2" place="2" resultid="2820" />
                    <RANKING order="3" place="3" resultid="3066" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2428" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4233" />
                    <RANKING order="2" place="2" resultid="3298" />
                    <RANKING order="3" place="3" resultid="3865" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2429" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4037" />
                    <RANKING order="2" place="2" resultid="2855" />
                    <RANKING order="3" place="-1" resultid="2953" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2430" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3686" />
                    <RANKING order="2" place="2" resultid="4726" />
                    <RANKING order="3" place="3" resultid="2835" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2431" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3086" />
                    <RANKING order="2" place="2" resultid="5058" />
                    <RANKING order="3" place="3" resultid="4693" />
                    <RANKING order="4" place="4" resultid="2165" />
                    <RANKING order="5" place="5" resultid="2173" />
                    <RANKING order="6" place="-1" resultid="4557" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2432" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3499" />
                    <RANKING order="2" place="2" resultid="3520" />
                    <RANKING order="3" place="3" resultid="4763" />
                    <RANKING order="4" place="4" resultid="3754" />
                    <RANKING order="5" place="5" resultid="3273" />
                    <RANKING order="6" place="6" resultid="4402" />
                    <RANKING order="7" place="7" resultid="3312" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2433" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3791" />
                    <RANKING order="2" place="2" resultid="3408" />
                    <RANKING order="3" place="3" resultid="3902" />
                    <RANKING order="4" place="4" resultid="4971" />
                    <RANKING order="5" place="5" resultid="5017" />
                    <RANKING order="6" place="6" resultid="4368" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2434" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2119" />
                    <RANKING order="2" place="2" resultid="2185" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2435" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4428" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2436" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="2437" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2438" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8013" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8014" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8015" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8016" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8017" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1318" daytime="12:10" gender="M" number="18" order="10" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1319" agemax="119" agemin="100" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="2978" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1320" agemax="159" agemin="120" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4301" />
                    <RANKING order="2" place="2" resultid="5227" />
                    <RANKING order="3" place="3" resultid="2980" />
                    <RANKING order="4" place="4" resultid="4171" />
                    <RANKING order="5" place="5" resultid="3375" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1321" agemax="199" agemin="160" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6431" />
                    <RANKING order="2" place="2" resultid="6171" />
                    <RANKING order="3" place="3" resultid="3159" />
                    <RANKING order="4" place="4" resultid="5070" />
                    <RANKING order="5" place="5" resultid="3867" />
                    <RANKING order="6" place="6" resultid="6038" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1322" agemax="239" agemin="200" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2979" />
                    <RANKING order="2" place="2" resultid="5463" />
                    <RANKING order="3" place="-1" resultid="3722" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1323" agemax="279" agemin="240" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4858" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1324" agemax="-1" agemin="280" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3950" />
                    <RANKING order="2" place="-1" resultid="3456" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8030" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8031" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1288" daytime="11:29" gender="M" number="16" order="8" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2454" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4310" />
                    <RANKING order="2" place="2" resultid="4438" />
                    <RANKING order="3" place="3" resultid="3195" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2455" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2896" />
                    <RANKING order="2" place="2" resultid="3606" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2456" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6028" />
                    <RANKING order="2" place="2" resultid="3345" />
                    <RANKING order="3" place="3" resultid="4277" />
                    <RANKING order="4" place="4" resultid="3676" />
                    <RANKING order="5" place="-1" resultid="4641" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2457" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5201" />
                    <RANKING order="2" place="2" resultid="3658" />
                    <RANKING order="3" place="3" resultid="4757" />
                    <RANKING order="4" place="4" resultid="3465" />
                    <RANKING order="5" place="5" resultid="3858" />
                    <RANKING order="6" place="6" resultid="4570" />
                    <RANKING order="7" place="7" resultid="4505" />
                    <RANKING order="8" place="8" resultid="4794" />
                    <RANKING order="9" place="9" resultid="3365" />
                    <RANKING order="10" place="10" resultid="3067" />
                    <RANKING order="11" place="-1" resultid="3171" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2458" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4718" />
                    <RANKING order="2" place="2" resultid="6428" />
                    <RANKING order="3" place="3" resultid="3959" />
                    <RANKING order="4" place="4" resultid="3324" />
                    <RANKING order="5" place="5" resultid="4249" />
                    <RANKING order="6" place="-1" resultid="3014" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2459" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5159" />
                    <RANKING order="2" place="2" resultid="4518" />
                    <RANKING order="3" place="3" resultid="2812" />
                    <RANKING order="4" place="4" resultid="4986" />
                    <RANKING order="5" place="5" resultid="3717" />
                    <RANKING order="6" place="6" resultid="3848" />
                    <RANKING order="7" place="7" resultid="4942" />
                    <RANKING order="8" place="8" resultid="3631" />
                    <RANKING order="9" place="-1" resultid="5165" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2460" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4851" />
                    <RANKING order="2" place="2" resultid="4711" />
                    <RANKING order="3" place="3" resultid="5747" />
                    <RANKING order="4" place="4" resultid="2836" />
                    <RANKING order="5" place="-1" resultid="4335" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2461" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4257" />
                    <RANKING order="2" place="2" resultid="2756" />
                    <RANKING order="3" place="3" resultid="3729" />
                    <RANKING order="4" place="4" resultid="2158" />
                    <RANKING order="5" place="5" resultid="2166" />
                    <RANKING order="6" place="6" resultid="2914" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2462" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2965" />
                    <RANKING order="2" place="2" resultid="5294" />
                    <RANKING order="3" place="3" resultid="4410" />
                    <RANKING order="4" place="4" resultid="3274" />
                    <RANKING order="5" place="5" resultid="5324" />
                    <RANKING order="6" place="6" resultid="4068" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2463" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4240" />
                    <RANKING order="2" place="2" resultid="4972" />
                    <RANKING order="3" place="3" resultid="3648" />
                    <RANKING order="4" place="4" resultid="3923" />
                    <RANKING order="5" place="5" resultid="4369" />
                    <RANKING order="6" place="6" resultid="4800" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2464" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="2465" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3425" />
                    <RANKING order="2" place="2" resultid="4844" />
                    <RANKING order="3" place="3" resultid="2772" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2466" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4017" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2467" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2468" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8022" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8023" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8024" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8025" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8026" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8027" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8028" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1213" daytime="09:53" gender="F" number="11" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2379" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4109" />
                    <RANKING order="2" place="2" resultid="3598" />
                    <RANKING order="3" place="3" resultid="3551" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2380" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3764" />
                    <RANKING order="2" place="2" resultid="2931" />
                    <RANKING order="3" place="3" resultid="3985" />
                    <RANKING order="4" place="4" resultid="2784" />
                    <RANKING order="5" place="5" resultid="4662" />
                    <RANKING order="6" place="6" resultid="3979" />
                    <RANKING order="7" place="7" resultid="4633" />
                    <RANKING order="8" place="8" resultid="2937" />
                    <RANKING order="9" place="-1" resultid="4608" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2381" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3974" />
                    <RANKING order="2" place="2" resultid="2920" />
                    <RANKING order="3" place="3" resultid="3490" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2382" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5407" />
                    <RANKING order="2" place="2" resultid="4511" />
                    <RANKING order="3" place="3" resultid="4870" />
                    <RANKING order="4" place="4" resultid="4778" />
                    <RANKING order="5" place="5" resultid="4880" />
                    <RANKING order="6" place="6" resultid="4094" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2383" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2947" />
                    <RANKING order="2" place="2" resultid="4200" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2384" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3875" />
                    <RANKING order="2" place="2" resultid="5177" />
                    <RANKING order="3" place="3" resultid="4679" />
                    <RANKING order="4" place="4" resultid="2750" />
                    <RANKING order="5" place="5" resultid="4700" />
                    <RANKING order="6" place="6" resultid="3043" />
                    <RANKING order="7" place="7" resultid="4043" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2385" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5066" />
                    <RANKING order="2" place="2" resultid="5389" />
                    <RANKING order="3" place="3" resultid="2860" />
                    <RANKING order="4" place="4" resultid="4564" />
                    <RANKING order="5" place="5" resultid="3670" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2386" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5279" />
                    <RANKING order="2" place="2" resultid="3935" />
                    <RANKING order="3" place="3" resultid="3050" />
                    <RANKING order="4" place="4" resultid="4455" />
                    <RANKING order="5" place="5" resultid="3447" />
                    <RANKING order="6" place="6" resultid="4446" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2387" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5360" />
                    <RANKING order="2" place="2" resultid="5366" />
                    <RANKING order="3" place="3" resultid="4196" />
                    <RANKING order="4" place="4" resultid="3434" />
                    <RANKING order="5" place="5" resultid="2828" />
                    <RANKING order="6" place="6" resultid="5103" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2388" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5272" />
                    <RANKING order="2" place="2" resultid="3911" />
                    <RANKING order="3" place="3" resultid="2890" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2389" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5135" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2390" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5355" />
                    <RANKING order="2" place="2" resultid="4010" />
                    <RANKING order="3" place="3" resultid="2227" />
                    <RANKING order="4" place="4" resultid="4002" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2391" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3017" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2392" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2393" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7994" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7995" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7996" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7997" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7998" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7999" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1273" daytime="11:07" gender="F" number="15" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2439" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4668" />
                    <RANKING order="2" place="2" resultid="4056" />
                    <RANKING order="3" place="3" resultid="3599" />
                    <RANKING order="4" place="-1" resultid="2849" />
                    <RANKING order="5" place="-1" resultid="3592" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2440" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2958" />
                    <RANKING order="2" place="2" resultid="4533" />
                    <RANKING order="3" place="3" resultid="5210" />
                    <RANKING order="4" place="4" resultid="2925" />
                    <RANKING order="5" place="5" resultid="4769" />
                    <RANKING order="6" place="6" resultid="5238" />
                    <RANKING order="7" place="-1" resultid="4328" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2441" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4074" />
                    <RANKING order="2" place="2" resultid="5192" />
                    <RANKING order="3" place="3" resultid="3509" />
                    <RANKING order="4" place="-1" resultid="2921" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2442" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4871" />
                    <RANKING order="2" place="2" resultid="2131" />
                    <RANKING order="3" place="3" resultid="3118" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2443" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5001" />
                    <RANKING order="2" place="2" resultid="4685" />
                    <RANKING order="3" place="3" resultid="5394" />
                    <RANKING order="4" place="4" resultid="4115" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2444" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5171" />
                    <RANKING order="2" place="2" resultid="3022" />
                    <RANKING order="3" place="3" resultid="4044" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2445" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5010" />
                    <RANKING order="2" place="2" resultid="4565" />
                    <RANKING order="3" place="3" resultid="3397" />
                    <RANKING order="4" place="4" resultid="3671" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2446" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4549" />
                    <RANKING order="2" place="2" resultid="2746" />
                    <RANKING order="3" place="3" resultid="4456" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2447" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3417" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2448" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5147" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2449" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="2450" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4957" />
                    <RANKING order="2" place="2" resultid="2228" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2451" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="2452" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2453" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8018" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8019" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8020" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8021" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1198" daytime="09:19" gender="M" number="10" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2364" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4207" />
                    <RANKING order="2" place="2" resultid="3706" />
                    <RANKING order="3" place="3" resultid="4386" />
                    <RANKING order="4" place="4" resultid="4437" />
                    <RANKING order="5" place="5" resultid="3796" />
                    <RANKING order="6" place="-1" resultid="3583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2365" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4376" />
                    <RANKING order="2" place="2" resultid="4219" />
                    <RANKING order="3" place="3" resultid="2882" />
                    <RANKING order="4" place="4" resultid="2822" />
                    <RANKING order="5" place="5" resultid="4080" />
                    <RANKING order="6" place="6" resultid="4271" />
                    <RANKING order="7" place="7" resultid="5253" />
                    <RANKING order="8" place="8" resultid="5245" />
                    <RANKING order="9" place="9" resultid="3357" />
                    <RANKING order="10" place="10" resultid="3339" />
                    <RANKING order="11" place="11" resultid="4626" />
                    <RANKING order="12" place="12" resultid="3351" />
                    <RANKING order="13" place="-1" resultid="3304" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2366" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4640" />
                    <RANKING order="2" place="2" resultid="4934" />
                    <RANKING order="3" place="3" resultid="4282" />
                    <RANKING order="4" place="4" resultid="4289" />
                    <RANKING order="5" place="-1" resultid="2125" />
                    <RANKING order="6" place="-1" resultid="3149" />
                    <RANKING order="7" place="-1" resultid="4574" />
                    <RANKING order="8" place="-1" resultid="4593" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2367" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4829" />
                    <RANKING order="2" place="2" resultid="5049" />
                    <RANKING order="3" place="3" resultid="4756" />
                    <RANKING order="4" place="4" resultid="3124" />
                    <RANKING order="5" place="5" resultid="4166" />
                    <RANKING order="6" place="6" resultid="4504" />
                    <RANKING order="7" place="7" resultid="2906" />
                    <RANKING order="8" place="8" resultid="5216" />
                    <RANKING order="9" place="9" resultid="4138" />
                    <RANKING order="10" place="10" resultid="4178" />
                    <RANKING order="11" place="11" resultid="5314" />
                    <RANKING order="12" place="12" resultid="2865" />
                    <RANKING order="13" place="13" resultid="2819" />
                    <RANKING order="14" place="14" resultid="2971" />
                    <RANKING order="15" place="15" resultid="4153" />
                    <RANKING order="16" place="16" resultid="3917" />
                    <RANKING order="17" place="17" resultid="3038" />
                    <RANKING order="18" place="18" resultid="4101" />
                    <RANKING order="19" place="-1" resultid="3857" />
                    <RANKING order="20" place="-1" resultid="6433" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2368" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4232" />
                    <RANKING order="2" place="2" resultid="6419" />
                    <RANKING order="3" place="3" resultid="3137" />
                    <RANKING order="4" place="4" resultid="4922" />
                    <RANKING order="5" place="5" resultid="4749" />
                    <RANKING order="6" place="6" resultid="4744" />
                    <RANKING order="7" place="7" resultid="4248" />
                    <RANKING order="8" place="8" resultid="4382" />
                    <RANKING order="9" place="9" resultid="4395" />
                    <RANKING order="10" place="10" resultid="4888" />
                    <RANKING order="11" place="11" resultid="3371" />
                    <RANKING order="12" place="12" resultid="2146" />
                    <RANKING order="13" place="13" resultid="3321" />
                    <RANKING order="14" place="14" resultid="3076" />
                    <RANKING order="15" place="15" resultid="4655" />
                    <RANKING order="16" place="16" resultid="4028" />
                    <RANKING order="17" place="17" resultid="3802" />
                    <RANKING order="18" place="18" resultid="4471" />
                    <RANKING order="19" place="-1" resultid="3130" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2369" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2779" />
                    <RANKING order="2" place="2" resultid="4525" />
                    <RANKING order="3" place="3" resultid="3282" />
                    <RANKING order="4" place="4" resultid="4985" />
                    <RANKING order="5" place="5" resultid="4062" />
                    <RANKING order="6" place="6" resultid="5184" />
                    <RANKING order="7" place="7" resultid="3843" />
                    <RANKING order="8" place="8" resultid="5441" />
                    <RANKING order="9" place="9" resultid="4941" />
                    <RANKING order="10" place="10" resultid="6415" />
                    <RANKING order="11" place="11" resultid="4901" />
                    <RANKING order="12" place="12" resultid="4418" />
                    <RANKING order="13" place="13" resultid="3515" />
                    <RANKING order="14" place="14" resultid="3328" />
                    <RANKING order="15" place="15" resultid="3612" />
                    <RANKING order="16" place="-1" resultid="4517" />
                    <RANKING order="17" place="-1" resultid="5448" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2370" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3699" />
                    <RANKING order="2" place="2" resultid="3782" />
                    <RANKING order="3" place="3" resultid="4850" />
                    <RANKING order="4" place="4" resultid="5479" />
                    <RANKING order="5" place="5" resultid="4725" />
                    <RANKING order="6" place="6" resultid="6424" />
                    <RANKING order="7" place="7" resultid="3574" />
                    <RANKING order="8" place="8" resultid="3810" />
                    <RANKING order="9" place="-1" resultid="5435" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2371" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2764" />
                    <RANKING order="2" place="2" resultid="4491" />
                    <RANKING order="3" place="3" resultid="4256" />
                    <RANKING order="4" place="4" resultid="4838" />
                    <RANKING order="5" place="5" resultid="2157" />
                    <RANKING order="6" place="6" resultid="5765" />
                    <RANKING order="7" place="7" resultid="5302" />
                    <RANKING order="8" place="8" resultid="3204" />
                    <RANKING order="9" place="9" resultid="2913" />
                    <RANKING order="10" place="10" resultid="5424" />
                    <RANKING order="11" place="-1" resultid="4964" />
                    <RANKING order="12" place="-1" resultid="5057" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2372" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4477" />
                    <RANKING order="2" place="2" resultid="3498" />
                    <RANKING order="3" place="3" resultid="4808" />
                    <RANKING order="4" place="4" resultid="3484" />
                    <RANKING order="5" place="5" resultid="3311" />
                    <RANKING order="6" place="6" resultid="4736" />
                    <RANKING order="7" place="7" resultid="3212" />
                    <RANKING order="8" place="8" resultid="4119" />
                    <RANKING order="9" place="-1" resultid="5323" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2373" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3901" />
                    <RANKING order="2" place="2" resultid="5116" />
                    <RANKING order="3" place="3" resultid="5016" />
                    <RANKING order="4" place="4" resultid="6439" />
                    <RANKING order="5" place="5" resultid="3387" />
                    <RANKING order="6" place="6" resultid="2798" />
                    <RANKING order="7" place="7" resultid="6019" />
                    <RANKING order="8" place="8" resultid="4799" />
                    <RANKING order="9" place="-1" resultid="3638" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2374" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2118" />
                    <RANKING order="2" place="2" resultid="2108" />
                    <RANKING order="3" place="3" resultid="3893" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2375" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2100" />
                    <RANKING order="2" place="2" resultid="4843" />
                    <RANKING order="3" place="3" resultid="3928" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2376" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4016" />
                    <RANKING order="2" place="2" resultid="3179" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2377" agemax="89" agemin="85" name="Kat. M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4086" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2378" agemax="94" agemin="90" name="Kat. N">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5076" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7980" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7981" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7982" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7983" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7984" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7985" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7986" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7987" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7988" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7989" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7990" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7991" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7992" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7993" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1243" daytime="10:28" gender="F" number="13" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2409" agemax="24" agemin="20" name="Kat. 0" />
                <AGEGROUP agegroupid="2410" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3104" />
                    <RANKING order="2" place="2" resultid="4634" />
                    <RANKING order="3" place="3" resultid="3059" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2411" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3968" />
                    <RANKING order="2" place="2" resultid="4821" />
                    <RANKING order="3" place="3" resultid="3471" />
                    <RANKING order="4" place="4" resultid="3093" />
                    <RANKING order="5" place="5" resultid="3887" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2412" agemax="39" agemin="35" name="Kat. C" />
                <AGEGROUP agegroupid="2413" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4996" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2414" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4263" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2415" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5095" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2416" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3448" />
                    <RANKING order="2" place="2" resultid="4447" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2417" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3416" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2418" agemax="69" agemin="65" name="Kat. I" />
                <AGEGROUP agegroupid="2419" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="2420" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="2421" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="2422" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2423" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8011" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8012" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1303" daytime="12:02" gender="F" number="17" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1304" agemax="119" agemin="100" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2977" />
                    <RANKING order="2" place="2" resultid="3989" />
                    <RANKING order="3" place="3" resultid="6101" />
                    <RANKING order="4" place="4" resultid="2976" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1305" agemax="159" agemin="120" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3158" />
                    <RANKING order="2" place="2" resultid="5228" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1306" agemax="199" agemin="160" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5462" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1307" agemax="239" agemin="200" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="5461" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1308" agemax="279" agemin="240" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3453" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1310" agemax="-1" agemin="280" name="Kat. F" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8029" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2015-06-27" daytime="15:00" name="III Blok" number="3" warmupfrom="14:00">
          <EVENTS>
            <EVENT eventid="1372" daytime="15:49" gender="M" number="22" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2514" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3772" />
                    <RANKING order="2" place="2" resultid="4209" />
                    <RANKING order="3" place="3" resultid="3145" />
                    <RANKING order="4" place="4" resultid="4440" />
                    <RANKING order="5" place="5" resultid="3797" />
                    <RANKING order="6" place="-1" resultid="3585" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2515" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4377" />
                    <RANKING order="2" place="2" resultid="2883" />
                    <RANKING order="3" place="3" resultid="4223" />
                    <RANKING order="4" place="4" resultid="4220" />
                    <RANKING order="5" place="5" resultid="5029" />
                    <RANKING order="6" place="6" resultid="4081" />
                    <RANKING order="7" place="7" resultid="2823" />
                    <RANKING order="8" place="8" resultid="4274" />
                    <RANKING order="9" place="9" resultid="5341" />
                    <RANKING order="10" place="10" resultid="3359" />
                    <RANKING order="11" place="11" resultid="4628" />
                    <RANKING order="12" place="12" resultid="5255" />
                    <RANKING order="13" place="13" resultid="4650" />
                    <RANKING order="14" place="14" resultid="3341" />
                    <RANKING order="15" place="15" resultid="3352" />
                    <RANKING order="16" place="-1" resultid="3305" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2516" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2138" />
                    <RANKING order="2" place="2" resultid="4642" />
                    <RANKING order="3" place="3" resultid="4285" />
                    <RANKING order="4" place="3" resultid="4298" />
                    <RANKING order="5" place="5" resultid="4935" />
                    <RANKING order="6" place="6" resultid="4291" />
                    <RANKING order="7" place="7" resultid="5225" />
                    <RANKING order="8" place="8" resultid="2843" />
                    <RANKING order="9" place="9" resultid="3150" />
                    <RANKING order="10" place="-1" resultid="2126" />
                    <RANKING order="11" place="-1" resultid="4575" />
                    <RANKING order="12" place="-1" resultid="4594" />
                    <RANKING order="13" place="-1" resultid="6000" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2517" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5051" />
                    <RANKING order="2" place="2" resultid="4139" />
                    <RANKING order="3" place="3" resultid="3125" />
                    <RANKING order="4" place="4" resultid="3565" />
                    <RANKING order="5" place="5" resultid="4579" />
                    <RANKING order="6" place="6" resultid="4168" />
                    <RANKING order="7" place="7" resultid="5316" />
                    <RANKING order="8" place="8" resultid="2907" />
                    <RANKING order="9" place="9" resultid="4759" />
                    <RANKING order="10" place="10" resultid="5217" />
                    <RANKING order="11" place="11" resultid="4179" />
                    <RANKING order="12" place="12" resultid="3860" />
                    <RANKING order="13" place="13" resultid="4160" />
                    <RANKING order="14" place="14" resultid="4150" />
                    <RANKING order="15" place="15" resultid="2972" />
                    <RANKING order="16" place="16" resultid="3919" />
                    <RANKING order="17" place="17" resultid="3039" />
                    <RANKING order="18" place="18" resultid="4133" />
                    <RANKING order="19" place="-1" resultid="4155" />
                    <RANKING order="20" place="-1" resultid="3030" />
                    <RANKING order="21" place="-1" resultid="6434" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2518" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4234" />
                    <RANKING order="2" place="2" resultid="6420" />
                    <RANKING order="3" place="3" resultid="3138" />
                    <RANKING order="4" place="4" resultid="4924" />
                    <RANKING order="5" place="5" resultid="2215" />
                    <RANKING order="6" place="6" resultid="3299" />
                    <RANKING order="7" place="7" resultid="2803" />
                    <RANKING order="8" place="8" resultid="4745" />
                    <RANKING order="9" place="9" resultid="4750" />
                    <RANKING order="10" place="10" resultid="4396" />
                    <RANKING order="11" place="11" resultid="4383" />
                    <RANKING order="12" place="12" resultid="3373" />
                    <RANKING order="13" place="12" resultid="4896" />
                    <RANKING order="14" place="14" resultid="2877" />
                    <RANKING order="15" place="15" resultid="4889" />
                    <RANKING order="16" place="16" resultid="4656" />
                    <RANKING order="17" place="17" resultid="4916" />
                    <RANKING order="18" place="18" resultid="2147" />
                    <RANKING order="19" place="19" resultid="3804" />
                    <RANKING order="20" place="20" resultid="3322" />
                    <RANKING order="21" place="21" resultid="4030" />
                    <RANKING order="22" place="22" resultid="4472" />
                    <RANKING order="23" place="-1" resultid="3026" />
                    <RANKING order="24" place="-1" resultid="3131" />
                    <RANKING order="25" place="-1" resultid="4214" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2519" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2780" />
                    <RANKING order="2" place="2" resultid="4526" />
                    <RANKING order="3" place="3" resultid="3283" />
                    <RANKING order="4" place="4" resultid="4520" />
                    <RANKING order="5" place="5" resultid="2743" />
                    <RANKING order="6" place="6" resultid="4988" />
                    <RANKING order="7" place="7" resultid="4064" />
                    <RANKING order="8" place="8" resultid="5443" />
                    <RANKING order="9" place="9" resultid="3844" />
                    <RANKING order="10" place="10" resultid="4943" />
                    <RANKING order="11" place="11" resultid="4420" />
                    <RANKING order="12" place="12" resultid="3516" />
                    <RANKING order="13" place="13" resultid="3329" />
                    <RANKING order="14" place="14" resultid="3614" />
                    <RANKING order="15" place="-1" resultid="3850" />
                    <RANKING order="16" place="-1" resultid="4903" />
                    <RANKING order="17" place="-1" resultid="5450" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2520" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3785" />
                    <RANKING order="2" place="2" resultid="4853" />
                    <RANKING order="3" place="3" resultid="5480" />
                    <RANKING order="4" place="4" resultid="5083" />
                    <RANKING order="5" place="5" resultid="4316" />
                    <RANKING order="6" place="6" resultid="3812" />
                    <RANKING order="7" place="-1" resultid="5436" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2521" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4493" />
                    <RANKING order="2" place="2" resultid="4840" />
                    <RANKING order="3" place="3" resultid="2160" />
                    <RANKING order="4" place="4" resultid="3293" />
                    <RANKING order="5" place="5" resultid="5305" />
                    <RANKING order="6" place="6" resultid="5766" />
                    <RANKING order="7" place="7" resultid="5419" />
                    <RANKING order="8" place="8" resultid="3206" />
                    <RANKING order="9" place="9" resultid="5425" />
                    <RANKING order="10" place="10" resultid="2915" />
                    <RANKING order="11" place="-1" resultid="4965" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2522" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2967" />
                    <RANKING order="2" place="2" resultid="4478" />
                    <RANKING order="3" place="3" resultid="4809" />
                    <RANKING order="4" place="4" resultid="3275" />
                    <RANKING order="5" place="5" resultid="3486" />
                    <RANKING order="6" place="6" resultid="3313" />
                    <RANKING order="7" place="7" resultid="3213" />
                    <RANKING order="8" place="8" resultid="4738" />
                    <RANKING order="9" place="9" resultid="4120" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2523" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5117" />
                    <RANKING order="2" place="2" resultid="5018" />
                    <RANKING order="3" place="3" resultid="3903" />
                    <RANKING order="4" place="4" resultid="3388" />
                    <RANKING order="5" place="5" resultid="2799" />
                    <RANKING order="6" place="6" resultid="6022" />
                    <RANKING order="7" place="7" resultid="5112" />
                    <RANKING order="8" place="-1" resultid="3641" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2524" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2110" />
                    <RANKING order="2" place="2" resultid="3895" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2525" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4846" />
                    <RANKING order="2" place="2" resultid="2101" />
                    <RANKING order="3" place="3" resultid="3930" />
                    <RANKING order="4" place="4" resultid="4025" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2526" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="2527" agemax="89" agemin="85" name="Kat. M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4088" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2528" agemax="94" agemin="90" name="Kat. N">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5078" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8051" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8052" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8053" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8054" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8055" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8056" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8057" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="8058" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="8059" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="8060" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="8061" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="8062" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="8063" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="8064" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="8065" number="15" order="15" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1402" daytime="16:42" gender="M" number="24" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2544" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4583" />
                    <RANKING order="2" place="2" resultid="3197" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2545" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3547" />
                    <RANKING order="2" place="2" resultid="5342" />
                    <RANKING order="3" place="3" resultid="3074" />
                    <RANKING order="4" place="4" resultid="2874" />
                    <RANKING order="5" place="5" resultid="5247" />
                    <RANKING order="6" place="6" resultid="3360" />
                    <RANKING order="7" place="7" resultid="3342" />
                    <RANKING order="8" place="8" resultid="3608" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2546" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2792" />
                    <RANKING order="2" place="2" resultid="5260" />
                    <RANKING order="3" place="3" resultid="2844" />
                    <RANKING order="4" place="-1" resultid="4145" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2547" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4831" />
                    <RANKING order="2" place="2" resultid="3126" />
                    <RANKING order="3" place="3" resultid="5317" />
                    <RANKING order="4" place="4" resultid="4161" />
                    <RANKING order="5" place="5" resultid="3920" />
                    <RANKING order="6" place="6" resultid="3068" />
                    <RANKING order="7" place="7" resultid="4104" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2548" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6412" />
                    <RANKING order="2" place="2" resultid="5348" />
                    <RANKING order="3" place="3" resultid="4917" />
                    <RANKING order="4" place="4" resultid="3961" />
                    <RANKING order="5" place="5" resultid="2152" />
                    <RANKING order="6" place="6" resultid="3079" />
                    <RANKING order="7" place="7" resultid="4052" />
                    <RANKING order="8" place="8" resultid="3805" />
                    <RANKING order="9" place="-1" resultid="3392" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2549" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5310" />
                    <RANKING order="2" place="2" resultid="6416" />
                    <RANKING order="3" place="3" resultid="5444" />
                    <RANKING order="4" place="4" resultid="4904" />
                    <RANKING order="5" place="5" resultid="4038" />
                    <RANKING order="6" place="6" resultid="2856" />
                    <RANKING order="7" place="7" resultid="3615" />
                    <RANKING order="8" place="-1" resultid="3633" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2550" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3682" />
                    <RANKING order="2" place="2" resultid="4713" />
                    <RANKING order="3" place="3" resultid="3154" />
                    <RANKING order="4" place="4" resultid="5431" />
                    <RANKING order="5" place="5" resultid="2838" />
                    <RANKING order="6" place="6" resultid="3576" />
                    <RANKING order="7" place="-1" resultid="3942" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2551" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4950" />
                    <RANKING order="2" place="2" resultid="2758" />
                    <RANKING order="3" place="3" resultid="3294" />
                    <RANKING order="4" place="4" resultid="5033" />
                    <RANKING order="5" place="5" resultid="4191" />
                    <RANKING order="6" place="6" resultid="2174" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2552" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3403" />
                    <RANKING order="2" place="2" resultid="3570" />
                    <RANKING order="3" place="3" resultid="3005" />
                    <RANKING order="4" place="4" resultid="4403" />
                    <RANKING order="5" place="5" resultid="4764" />
                    <RANKING order="6" place="6" resultid="3755" />
                    <RANKING order="7" place="7" resultid="4739" />
                    <RANKING order="8" place="8" resultid="4070" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2553" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4992" />
                    <RANKING order="2" place="2" resultid="5024" />
                    <RANKING order="3" place="3" resultid="3409" />
                    <RANKING order="4" place="4" resultid="3650" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2554" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2186" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2555" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5126" />
                    <RANKING order="2" place="2" resultid="3427" />
                    <RANKING order="3" place="3" resultid="4429" />
                    <RANKING order="4" place="4" resultid="2774" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2556" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3382" />
                    <RANKING order="2" place="2" resultid="3181" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2557" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2558" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8071" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8072" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8073" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8074" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8075" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8076" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8077" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1432" daytime="17:58" gender="M" number="26" order="8" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2574" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3708" />
                    <RANKING order="2" place="2" resultid="4312" />
                    <RANKING order="3" place="3" resultid="3798" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2575" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3010" />
                    <RANKING order="2" place="2" resultid="2201" />
                    <RANKING order="3" place="3" resultid="5248" />
                    <RANKING order="4" place="4" resultid="4184" />
                    <RANKING order="5" place="5" resultid="5256" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2576" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2793" />
                    <RANKING order="2" place="2" resultid="4643" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2577" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3659" />
                    <RANKING order="2" place="2" resultid="8292" />
                    <RANKING order="3" place="3" resultid="4507" />
                    <RANKING order="4" place="4" resultid="2866" />
                    <RANKING order="5" place="5" resultid="4169" />
                    <RANKING order="6" place="6" resultid="2973" />
                    <RANKING order="7" place="-1" resultid="4134" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2578" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8291" />
                    <RANKING order="2" place="2" resultid="3139" />
                    <RANKING order="3" place="3" resultid="3015" />
                    <RANKING order="4" place="4" resultid="6421" />
                    <RANKING order="5" place="5" resultid="4925" />
                    <RANKING order="6" place="6" resultid="4251" />
                    <RANKING order="7" place="7" resultid="4890" />
                    <RANKING order="8" place="8" resultid="2148" />
                    <RANKING order="9" place="9" resultid="8290" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2579" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4527" />
                    <RANKING order="2" place="2" resultid="8326" />
                    <RANKING order="3" place="3" resultid="3719" />
                    <RANKING order="4" place="4" resultid="4944" />
                    <RANKING order="5" place="5" resultid="3845" />
                    <RANKING order="6" place="6" resultid="4421" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2580" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8289" />
                    <RANKING order="2" place="2" resultid="6425" />
                    <RANKING order="3" place="3" resultid="4727" />
                    <RANKING order="4" place="4" resultid="3155" />
                    <RANKING order="5" place="5" resultid="5154" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2581" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3087" />
                    <RANKING order="2" place="2" resultid="4694" />
                    <RANKING order="3" place="3" resultid="4558" />
                    <RANKING order="4" place="4" resultid="5426" />
                    <RANKING order="5" place="5" resultid="2916" />
                    <RANKING order="6" place="6" resultid="3735" />
                    <RANKING order="7" place="7" resultid="3207" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2582" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3500" />
                    <RANKING order="2" place="2" resultid="3521" />
                    <RANKING order="3" place="3" resultid="8327" />
                    <RANKING order="4" place="4" resultid="5296" />
                    <RANKING order="5" place="5" resultid="4404" />
                    <RANKING order="6" place="6" resultid="3314" />
                    <RANKING order="7" place="7" resultid="3214" />
                    <RANKING order="8" place="-1" resultid="5326" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2583" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4242" />
                    <RANKING order="2" place="2" resultid="3792" />
                    <RANKING order="3" place="3" resultid="3904" />
                    <RANKING order="4" place="4" resultid="6440" />
                    <RANKING order="5" place="5" resultid="4801" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2584" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2120" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2585" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2102" />
                    <RANKING order="2" place="2" resultid="3931" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2586" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4019" />
                    <RANKING order="2" place="2" resultid="8336" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2587" agemax="89" agemin="85" name="Kat. M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4089" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2588" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8151" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8152" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8153" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8154" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8155" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8156" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8325" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1326" daytime="15:00" gender="F" number="19" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2469" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4669" />
                    <RANKING order="2" place="2" resultid="4057" />
                    <RANKING order="3" place="-1" resultid="3593" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2470" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3765" />
                    <RANKING order="2" place="2" resultid="2959" />
                    <RANKING order="3" place="3" resultid="3986" />
                    <RANKING order="4" place="4" resultid="4534" />
                    <RANKING order="5" place="5" resultid="2926" />
                    <RANKING order="6" place="6" resultid="5239" />
                    <RANKING order="7" place="-1" resultid="4329" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2471" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4075" />
                    <RANKING order="2" place="2" resultid="3318" />
                    <RANKING order="3" place="3" resultid="5193" />
                    <RANKING order="4" place="4" resultid="3510" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2472" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4872" />
                    <RANKING order="2" place="2" resultid="2132" />
                    <RANKING order="3" place="3" resultid="3119" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2473" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5002" />
                    <RANKING order="2" place="2" resultid="4686" />
                    <RANKING order="3" place="3" resultid="5395" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2474" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3876" />
                    <RANKING order="2" place="2" resultid="5172" />
                    <RANKING order="3" place="3" resultid="4680" />
                    <RANKING order="4" place="4" resultid="4045" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2475" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5011" />
                    <RANKING order="2" place="2" resultid="3693" />
                    <RANKING order="3" place="3" resultid="3672" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2476" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4550" />
                    <RANKING order="2" place="2" resultid="2747" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2477" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3418" />
                    <RANKING order="2" place="2" resultid="5104" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2478" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2806" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2479" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3441" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2480" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4958" />
                    <RANKING order="2" place="2" resultid="2229" />
                    <RANKING order="3" place="3" resultid="4003" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2481" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="2482" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2483" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8032" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8033" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8034" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8035" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1417" daytime="17:22" gender="F" number="25" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2559" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4622" />
                    <RANKING order="2" place="2" resultid="2851" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2560" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2960" />
                    <RANKING order="2" place="2" resultid="4771" />
                    <RANKING order="3" place="3" resultid="3060" />
                    <RANKING order="4" place="4" resultid="5090" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2561" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3099" />
                    <RANKING order="2" place="2" resultid="4541" />
                    <RANKING order="3" place="3" resultid="3094" />
                    <RANKING order="4" place="4" resultid="4589" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2562" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5760" />
                    <RANKING order="2" place="2" resultid="4873" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2563" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5142" />
                    <RANKING order="2" place="2" resultid="5403" />
                    <RANKING order="3" place="3" resultid="4687" />
                    <RANKING order="4" place="4" resultid="4116" />
                    <RANKING order="5" place="5" resultid="3949" />
                    <RANKING order="6" place="6" resultid="3741" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2564" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3665" />
                    <RANKING order="2" place="2" resultid="3023" />
                    <RANKING order="3" place="3" resultid="4865" />
                    <RANKING order="4" place="4" resultid="3112" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2565" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3289" />
                    <RANKING order="2" place="2" resultid="3694" />
                    <RANKING order="3" place="3" resultid="3398" />
                    <RANKING order="4" place="4" resultid="5096" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2566" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4500" />
                    <RANKING order="2" place="2" resultid="3052" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2567" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3626" />
                    <RANKING order="2" place="2" resultid="5105" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2568" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5274" />
                    <RANKING order="2" place="2" resultid="2892" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2569" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="2570" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4959" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2571" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="2572" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2573" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8147" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8148" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8149" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8150" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1342" daytime="15:13" gender="M" number="20" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2484" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4208" />
                    <RANKING order="2" place="2" resultid="4311" />
                    <RANKING order="3" place="3" resultid="4439" />
                    <RANKING order="4" place="4" resultid="3196" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2485" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4273" />
                    <RANKING order="2" place="2" resultid="2897" />
                    <RANKING order="3" place="3" resultid="3607" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2486" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6029" />
                    <RANKING order="2" place="2" resultid="3346" />
                    <RANKING order="3" place="3" resultid="4278" />
                    <RANKING order="4" place="4" resultid="3677" />
                    <RANKING order="5" place="5" resultid="4284" />
                    <RANKING order="6" place="-1" resultid="4144" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2487" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5202" />
                    <RANKING order="2" place="2" resultid="3466" />
                    <RANKING order="3" place="3" resultid="4758" />
                    <RANKING order="4" place="4" resultid="3172" />
                    <RANKING order="5" place="5" resultid="4571" />
                    <RANKING order="6" place="6" resultid="3859" />
                    <RANKING order="7" place="7" resultid="4795" />
                    <RANKING order="8" place="8" resultid="3366" />
                    <RANKING order="9" place="9" resultid="4103" />
                    <RANKING order="10" place="-1" resultid="4506" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2488" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4719" />
                    <RANKING order="2" place="2" resultid="5189" />
                    <RANKING order="3" place="3" resultid="6429" />
                    <RANKING order="4" place="4" resultid="3325" />
                    <RANKING order="5" place="5" resultid="3960" />
                    <RANKING order="6" place="6" resultid="4250" />
                    <RANKING order="7" place="7" resultid="3391" />
                    <RANKING order="8" place="-1" resultid="4213" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2489" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5160" />
                    <RANKING order="2" place="2" resultid="4519" />
                    <RANKING order="3" place="3" resultid="2813" />
                    <RANKING order="4" place="4" resultid="4987" />
                    <RANKING order="5" place="5" resultid="3849" />
                    <RANKING order="6" place="6" resultid="3718" />
                    <RANKING order="7" place="7" resultid="5166" />
                    <RANKING order="8" place="8" resultid="3632" />
                    <RANKING order="9" place="-1" resultid="5449" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2490" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4852" />
                    <RANKING order="2" place="2" resultid="4712" />
                    <RANKING order="3" place="3" resultid="3784" />
                    <RANKING order="4" place="4" resultid="5748" />
                    <RANKING order="5" place="5" resultid="2837" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2491" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6034" />
                    <RANKING order="2" place="2" resultid="4258" />
                    <RANKING order="3" place="3" resultid="4492" />
                    <RANKING order="4" place="4" resultid="3730" />
                    <RANKING order="5" place="5" resultid="4190" />
                    <RANKING order="6" place="6" resultid="4839" />
                    <RANKING order="7" place="7" resultid="5304" />
                    <RANKING order="8" place="8" resultid="2159" />
                    <RANKING order="9" place="-1" resultid="2167" />
                    <RANKING order="10" place="-1" resultid="2757" />
                    <RANKING order="11" place="-1" resultid="5059" />
                    <RANKING order="12" place="-1" resultid="5418" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2492" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2966" />
                    <RANKING order="2" place="2" resultid="5295" />
                    <RANKING order="3" place="3" resultid="4411" />
                    <RANKING order="4" place="4" resultid="5289" />
                    <RANKING order="5" place="5" resultid="5325" />
                    <RANKING order="6" place="6" resultid="4815" />
                    <RANKING order="7" place="7" resultid="4069" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2493" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4241" />
                    <RANKING order="2" place="2" resultid="4973" />
                    <RANKING order="3" place="3" resultid="3649" />
                    <RANKING order="4" place="4" resultid="4370" />
                    <RANKING order="5" place="5" resultid="5111" />
                    <RANKING order="6" place="6" resultid="3924" />
                    <RANKING order="7" place="-1" resultid="6021" />
                    <RANKING order="8" place="-1" resultid="3640" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2494" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3894" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2495" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3426" />
                    <RANKING order="2" place="2" resultid="4845" />
                    <RANKING order="3" place="3" resultid="2773" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2496" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4018" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2497" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2498" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8036" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8037" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8038" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8039" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8040" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8041" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8042" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="8043" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1357" daytime="15:36" gender="F" number="21" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2499" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4110" />
                    <RANKING order="2" place="2" resultid="5266" />
                    <RANKING order="3" place="3" resultid="4621" />
                    <RANKING order="4" place="4" resultid="3600" />
                    <RANKING order="5" place="5" resultid="2850" />
                    <RANKING order="6" place="6" resultid="3552" />
                    <RANKING order="7" place="7" resultid="4616" />
                    <RANKING order="8" place="8" resultid="4670" />
                    <RANKING order="9" place="-1" resultid="3594" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2500" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5413" />
                    <RANKING order="2" place="2" resultid="3766" />
                    <RANKING order="3" place="3" resultid="5038" />
                    <RANKING order="4" place="4" resultid="4663" />
                    <RANKING order="5" place="5" resultid="3987" />
                    <RANKING order="6" place="6" resultid="4599" />
                    <RANKING order="7" place="7" resultid="5211" />
                    <RANKING order="8" place="8" resultid="4535" />
                    <RANKING order="9" place="9" resultid="5240" />
                    <RANKING order="10" place="10" resultid="3105" />
                    <RANKING order="11" place="11" resultid="2902" />
                    <RANKING order="12" place="12" resultid="2938" />
                    <RANKING order="13" place="13" resultid="5089" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2501" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2870" />
                    <RANKING order="2" place="2" resultid="3969" />
                    <RANKING order="3" place="3" resultid="4588" />
                    <RANKING order="4" place="4" resultid="3491" />
                    <RANKING order="5" place="5" resultid="4540" />
                    <RANKING order="6" place="6" resultid="3888" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2502" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4909" />
                    <RANKING order="2" place="2" resultid="3120" />
                    <RANKING order="3" place="3" resultid="5198" />
                    <RANKING order="4" place="4" resultid="4881" />
                    <RANKING order="5" place="5" resultid="2133" />
                    <RANKING order="6" place="6" resultid="4779" />
                    <RANKING order="7" place="7" resultid="4095" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2503" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5003" />
                    <RANKING order="2" place="2" resultid="5396" />
                    <RANKING order="3" place="3" resultid="2948" />
                    <RANKING order="4" place="4" resultid="5402" />
                    <RANKING order="5" place="5" resultid="3948" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2504" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3664" />
                    <RANKING order="2" place="2" resultid="3877" />
                    <RANKING order="3" place="3" resultid="5178" />
                    <RANKING order="4" place="4" resultid="4681" />
                    <RANKING order="5" place="5" resultid="5173" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2505" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5067" />
                    <RANKING order="2" place="2" resultid="5379" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2506" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5374" />
                    <RANKING order="2" place="2" resultid="3883" />
                    <RANKING order="3" place="3" resultid="4499" />
                    <RANKING order="4" place="4" resultid="3051" />
                    <RANKING order="5" place="5" resultid="3747" />
                    <RANKING order="6" place="6" resultid="5755" />
                    <RANKING order="7" place="7" resultid="4457" />
                    <RANKING order="8" place="8" resultid="5285" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2507" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5367" />
                    <RANKING order="2" place="2" resultid="3435" />
                    <RANKING order="3" place="3" resultid="3625" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2508" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5273" />
                    <RANKING order="2" place="2" resultid="2807" />
                    <RANKING order="3" place="3" resultid="5148" />
                    <RANKING order="4" place="4" resultid="2891" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2509" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3442" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2510" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5356" />
                    <RANKING order="2" place="2" resultid="4004" />
                    <RANKING order="3" place="3" resultid="2230" />
                    <RANKING order="4" place="4" resultid="4011" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2511" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="2512" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2513" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8044" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8045" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8046" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8047" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8048" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8049" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8050" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1447" daytime="19:01" gender="F" number="27" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2589" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2590" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5212" />
                    <RANKING order="2" place="2" resultid="3106" />
                    <RANKING order="3" place="3" resultid="2786" />
                    <RANKING order="4" place="4" resultid="3980" />
                    <RANKING order="5" place="5" resultid="2927" />
                    <RANKING order="6" place="6" resultid="4635" />
                    <RANKING order="7" place="7" resultid="3061" />
                    <RANKING order="8" place="-1" resultid="4330" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2591" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2871" />
                    <RANKING order="2" place="2" resultid="3970" />
                    <RANKING order="3" place="3" resultid="3472" />
                    <RANKING order="4" place="4" resultid="4823" />
                    <RANKING order="5" place="5" resultid="3095" />
                    <RANKING order="6" place="6" resultid="2943" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2592" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4882" />
                    <RANKING order="2" place="2" resultid="5199" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2593" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4997" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2594" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4701" />
                    <RANKING order="2" place="2" resultid="4265" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2595" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5012" />
                    <RANKING order="2" place="2" resultid="3290" />
                    <RANKING order="3" place="3" resultid="5097" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2596" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5375" />
                    <RANKING order="2" place="2" resultid="4551" />
                    <RANKING order="3" place="3" resultid="3748" />
                    <RANKING order="4" place="4" resultid="4449" />
                    <RANKING order="5" place="-1" resultid="3450" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2597" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3419" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2598" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3913" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2599" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="2600" agemax="79" agemin="75" name="Kat. K" />
                <AGEGROUP agegroupid="2601" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="2602" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2603" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8078" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8079" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8080" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1387" daytime="16:13" gender="F" number="23" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2529" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4111" />
                    <RANKING order="2" place="2" resultid="3601" />
                    <RANKING order="3" place="3" resultid="3553" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2530" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2932" />
                    <RANKING order="2" place="2" resultid="2785" />
                    <RANKING order="3" place="3" resultid="4609" />
                    <RANKING order="4" place="4" resultid="4770" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2531" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4822" />
                    <RANKING order="2" place="2" resultid="5206" />
                    <RANKING order="3" place="3" resultid="3975" />
                    <RANKING order="4" place="4" resultid="2922" />
                    <RANKING order="5" place="5" resultid="3511" />
                    <RANKING order="6" place="6" resultid="3492" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2532" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5408" />
                    <RANKING order="2" place="2" resultid="4512" />
                    <RANKING order="3" place="3" resultid="4780" />
                    <RANKING order="4" place="4" resultid="4096" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2533" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5141" />
                    <RANKING order="2" place="2" resultid="2949" />
                    <RANKING order="3" place="3" resultid="4201" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2534" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3111" />
                    <RANKING order="2" place="2" resultid="2751" />
                    <RANKING order="3" place="3" resultid="4264" />
                    <RANKING order="4" place="4" resultid="3044" />
                    <RANKING order="5" place="5" resultid="4046" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2535" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5390" />
                    <RANKING order="2" place="2" resultid="2861" />
                    <RANKING order="3" place="3" resultid="4566" />
                    <RANKING order="4" place="4" resultid="3673" />
                    <RANKING order="5" place="-1" resultid="5068" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2536" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3936" />
                    <RANKING order="2" place="2" resultid="5280" />
                    <RANKING order="3" place="3" resultid="4458" />
                    <RANKING order="4" place="4" resultid="4448" />
                    <RANKING order="5" place="5" resultid="3449" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2537" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5361" />
                    <RANKING order="2" place="2" resultid="5368" />
                    <RANKING order="3" place="3" resultid="4197" />
                    <RANKING order="4" place="4" resultid="3436" />
                    <RANKING order="5" place="5" resultid="2829" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2538" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3912" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2539" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5136" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2540" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4012" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2541" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3018" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2542" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2543" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8066" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8067" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8068" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8069" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8070" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1462" daytime="19:13" gender="M" number="28" order="10" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2604" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4387" />
                    <RANKING order="2" place="2" resultid="3709" />
                    <RANKING order="3" place="3" resultid="4322" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2605" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5044" />
                    <RANKING order="2" place="2" resultid="2884" />
                    <RANKING order="3" place="3" resultid="2898" />
                    <RANKING order="4" place="4" resultid="4651" />
                    <RANKING order="5" place="5" resultid="4629" />
                    <RANKING order="6" place="6" resultid="2824" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2606" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4299" />
                    <RANKING order="2" place="2" resultid="4788" />
                    <RANKING order="3" place="-1" resultid="4595" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2607" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4832" />
                    <RANKING order="2" place="2" resultid="3467" />
                    <RANKING order="3" place="3" resultid="3660" />
                    <RANKING order="4" place="4" resultid="5052" />
                    <RANKING order="5" place="5" resultid="3367" />
                    <RANKING order="6" place="6" resultid="4796" />
                    <RANKING order="7" place="7" resultid="3069" />
                    <RANKING order="8" place="-1" resultid="3173" />
                    <RANKING order="9" place="-1" resultid="4180" />
                    <RANKING order="10" place="-1" resultid="6435" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2608" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4235" />
                    <RANKING order="2" place="2" resultid="3300" />
                    <RANKING order="3" place="3" resultid="4897" />
                    <RANKING order="4" place="4" resultid="4657" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2609" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2954" />
                    <RANKING order="2" place="2" resultid="5167" />
                    <RANKING order="3" place="3" resultid="4039" />
                    <RANKING order="4" place="4" resultid="3330" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2610" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5481" />
                    <RANKING order="2" place="2" resultid="3687" />
                    <RANKING order="3" place="3" resultid="4728" />
                    <RANKING order="4" place="4" resultid="5749" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2611" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5060" />
                    <RANKING order="2" place="2" resultid="4695" />
                    <RANKING order="3" place="3" resultid="2168" />
                    <RANKING order="4" place="-1" resultid="4559" />
                    <RANKING order="5" place="-1" resultid="4966" />
                    <RANKING order="6" place="-1" resultid="5767" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2612" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3501" />
                    <RANKING order="2" place="2" resultid="4412" />
                    <RANKING order="3" place="3" resultid="3522" />
                    <RANKING order="4" place="4" resultid="4810" />
                    <RANKING order="5" place="5" resultid="3756" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2613" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5019" />
                    <RANKING order="2" place="2" resultid="3410" />
                    <RANKING order="3" place="3" resultid="4974" />
                    <RANKING order="4" place="4" resultid="4371" />
                    <RANKING order="5" place="5" resultid="4802" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2614" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2111" />
                    <RANKING order="2" place="2" resultid="2187" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2615" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4430" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2616" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="2617" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2618" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8081" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8082" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8083" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8084" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8085" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8086" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2015-06-28" daytime="09:00" name="IV Blok" number="4" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="1509" daytime="09:28" gender="M" number="30" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2634" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3710" />
                    <RANKING order="2" place="2" resultid="4313" />
                    <RANKING order="3" place="3" resultid="4441" />
                    <RANKING order="4" place="-1" resultid="3198" />
                    <RANKING order="5" place="-1" resultid="3587" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2635" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2202" />
                    <RANKING order="2" place="2" resultid="2825" />
                    <RANKING order="3" place="3" resultid="5249" />
                    <RANKING order="4" place="4" resultid="4082" />
                    <RANKING order="5" place="5" resultid="3361" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2636" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4644" />
                    <RANKING order="2" place="2" resultid="4936" />
                    <RANKING order="3" place="3" resultid="3151" />
                    <RANKING order="4" place="4" resultid="4789" />
                    <RANKING order="5" place="-1" resultid="4576" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2637" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4833" />
                    <RANKING order="2" place="2" resultid="3661" />
                    <RANKING order="3" place="3" resultid="2909" />
                    <RANKING order="4" place="4" resultid="4170" />
                    <RANKING order="5" place="5" resultid="4508" />
                    <RANKING order="6" place="6" resultid="2867" />
                    <RANKING order="7" place="7" resultid="3070" />
                    <RANKING order="8" place="8" resultid="2974" />
                    <RANKING order="9" place="9" resultid="4140" />
                    <RANKING order="10" place="10" resultid="3040" />
                    <RANKING order="11" place="-1" resultid="3032" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2638" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4236" />
                    <RANKING order="2" place="2" resultid="3140" />
                    <RANKING order="3" place="3" resultid="6422" />
                    <RANKING order="4" place="4" resultid="4926" />
                    <RANKING order="5" place="5" resultid="3133" />
                    <RANKING order="6" place="6" resultid="4891" />
                    <RANKING order="7" place="7" resultid="4752" />
                    <RANKING order="8" place="8" resultid="4252" />
                    <RANKING order="9" place="9" resultid="2878" />
                    <RANKING order="10" place="10" resultid="4746" />
                    <RANKING order="11" place="11" resultid="2149" />
                    <RANKING order="12" place="12" resultid="4658" />
                    <RANKING order="13" place="13" resultid="4032" />
                    <RANKING order="14" place="14" resultid="4473" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2639" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2781" />
                    <RANKING order="2" place="2" resultid="4528" />
                    <RANKING order="3" place="3" resultid="2955" />
                    <RANKING order="4" place="4" resultid="5455" />
                    <RANKING order="5" place="5" resultid="2814" />
                    <RANKING order="6" place="6" resultid="5445" />
                    <RANKING order="7" place="7" resultid="3846" />
                    <RANKING order="8" place="8" resultid="4945" />
                    <RANKING order="9" place="9" resultid="4422" />
                    <RANKING order="10" place="10" resultid="3331" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2640" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3701" />
                    <RANKING order="2" place="2" resultid="5482" />
                    <RANKING order="3" place="3" resultid="6426" />
                    <RANKING order="4" place="4" resultid="4729" />
                    <RANKING order="5" place="5" resultid="5155" />
                    <RANKING order="6" place="6" resultid="3688" />
                    <RANKING order="7" place="7" resultid="3577" />
                    <RANKING order="8" place="-1" resultid="3156" />
                    <RANKING order="9" place="-1" resultid="4337" />
                    <RANKING order="10" place="-1" resultid="5438" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2641" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2766" />
                    <RANKING order="2" place="2" resultid="5061" />
                    <RANKING order="3" place="3" resultid="4951" />
                    <RANKING order="4" place="4" resultid="4560" />
                    <RANKING order="5" place="5" resultid="5768" />
                    <RANKING order="6" place="6" resultid="3731" />
                    <RANKING order="7" place="7" resultid="5427" />
                    <RANKING order="8" place="8" resultid="3208" />
                    <RANKING order="9" place="9" resultid="3736" />
                    <RANKING order="10" place="10" resultid="2917" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2642" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2968" />
                    <RANKING order="2" place="2" resultid="3502" />
                    <RANKING order="3" place="3" resultid="4479" />
                    <RANKING order="4" place="4" resultid="4811" />
                    <RANKING order="5" place="5" resultid="3854" />
                    <RANKING order="6" place="6" resultid="3315" />
                    <RANKING order="7" place="7" resultid="3215" />
                    <RANKING order="8" place="8" resultid="4740" />
                    <RANKING order="9" place="9" resultid="4121" />
                    <RANKING order="10" place="-1" resultid="3523" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2643" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3905" />
                    <RANKING order="2" place="2" resultid="6441" />
                    <RANKING order="3" place="3" resultid="4803" />
                    <RANKING order="4" place="4" resultid="4372" />
                    <RANKING order="5" place="-1" resultid="3642" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2644" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2121" />
                    <RANKING order="2" place="2" resultid="2112" />
                    <RANKING order="3" place="3" resultid="2188" />
                    <RANKING order="4" place="4" resultid="3896" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2645" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2103" />
                    <RANKING order="2" place="2" resultid="3932" />
                    <RANKING order="3" place="3" resultid="4847" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2646" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4020" />
                    <RANKING order="2" place="2" resultid="3183" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2647" agemax="89" agemin="85" name="Kat. M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4090" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2648" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8093" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8094" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8095" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8096" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8097" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8098" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8099" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="8100" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="8101" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="8102" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1539" daytime="10:26" gender="M" number="32" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2664" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3773" />
                    <RANKING order="2" place="2" resultid="4210" />
                    <RANKING order="3" place="3" resultid="4442" />
                    <RANKING order="4" place="-1" resultid="3199" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2665" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4378" />
                    <RANKING order="2" place="2" resultid="2899" />
                    <RANKING order="3" place="3" resultid="4275" />
                    <RANKING order="4" place="4" resultid="2826" />
                    <RANKING order="5" place="5" resultid="2885" />
                    <RANKING order="6" place="-1" resultid="3353" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2666" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4300" />
                    <RANKING order="2" place="2" resultid="6030" />
                    <RANKING order="3" place="3" resultid="4279" />
                    <RANKING order="4" place="4" resultid="4286" />
                    <RANKING order="5" place="5" resultid="3678" />
                    <RANKING order="6" place="6" resultid="4146" />
                    <RANKING order="7" place="-1" resultid="3347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2667" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3468" />
                    <RANKING order="2" place="2" resultid="5203" />
                    <RANKING order="3" place="3" resultid="5053" />
                    <RANKING order="4" place="4" resultid="4760" />
                    <RANKING order="5" place="5" resultid="3861" />
                    <RANKING order="6" place="6" resultid="3368" />
                    <RANKING order="7" place="7" resultid="4135" />
                    <RANKING order="8" place="8" resultid="4797" />
                    <RANKING order="9" place="9" resultid="3174" />
                    <RANKING order="10" place="10" resultid="4156" />
                    <RANKING order="11" place="11" resultid="2975" />
                    <RANKING order="12" place="12" resultid="4105" />
                    <RANKING order="13" place="-1" resultid="3566" />
                    <RANKING order="14" place="-1" resultid="4572" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2668" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4720" />
                    <RANKING order="2" place="2" resultid="5190" />
                    <RANKING order="3" place="3" resultid="3326" />
                    <RANKING order="4" place="4" resultid="6430" />
                    <RANKING order="5" place="5" resultid="4898" />
                    <RANKING order="6" place="6" resultid="3393" />
                    <RANKING order="7" place="7" resultid="4033" />
                    <RANKING order="8" place="-1" resultid="3806" />
                    <RANKING order="9" place="-1" resultid="4215" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2669" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5161" />
                    <RANKING order="2" place="2" resultid="4521" />
                    <RANKING order="3" place="3" resultid="2744" />
                    <RANKING order="4" place="4" resultid="3284" />
                    <RANKING order="5" place="5" resultid="2815" />
                    <RANKING order="6" place="6" resultid="3720" />
                    <RANKING order="7" place="7" resultid="5168" />
                    <RANKING order="8" place="8" resultid="4946" />
                    <RANKING order="9" place="9" resultid="3634" />
                    <RANKING order="10" place="-1" resultid="3851" />
                    <RANKING order="11" place="-1" resultid="5451" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2670" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4854" />
                    <RANKING order="2" place="2" resultid="4714" />
                    <RANKING order="3" place="3" resultid="3786" />
                    <RANKING order="4" place="4" resultid="5084" />
                    <RANKING order="5" place="5" resultid="3702" />
                    <RANKING order="6" place="6" resultid="5750" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2671" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6035" />
                    <RANKING order="2" place="2" resultid="3088" />
                    <RANKING order="3" place="3" resultid="4494" />
                    <RANKING order="4" place="4" resultid="2759" />
                    <RANKING order="5" place="5" resultid="2161" />
                    <RANKING order="6" place="6" resultid="4841" />
                    <RANKING order="7" place="7" resultid="5306" />
                    <RANKING order="8" place="8" resultid="3732" />
                    <RANKING order="9" place="9" resultid="4192" />
                    <RANKING order="10" place="10" resultid="3209" />
                    <RANKING order="11" place="11" resultid="2918" />
                    <RANKING order="12" place="-1" resultid="5062" />
                    <RANKING order="13" place="-1" resultid="5420" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2672" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3277" />
                    <RANKING order="2" place="2" resultid="5328" />
                    <RANKING order="3" place="3" resultid="5290" />
                    <RANKING order="4" place="4" resultid="4413" />
                    <RANKING order="5" place="5" resultid="5297" />
                    <RANKING order="6" place="6" resultid="4816" />
                    <RANKING order="7" place="7" resultid="3216" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2673" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4243" />
                    <RANKING order="2" place="2" resultid="5118" />
                    <RANKING order="3" place="3" resultid="5020" />
                    <RANKING order="4" place="4" resultid="4975" />
                    <RANKING order="5" place="5" resultid="3651" />
                    <RANKING order="6" place="6" resultid="5113" />
                    <RANKING order="7" place="7" resultid="2800" />
                    <RANKING order="8" place="8" resultid="3925" />
                    <RANKING order="9" place="9" resultid="6023" />
                    <RANKING order="10" place="-1" resultid="3643" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2674" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3897" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2675" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3428" />
                    <RANKING order="2" place="2" resultid="4848" />
                    <RANKING order="3" place="3" resultid="2775" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2676" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3383" />
                    <RANKING order="2" place="2" resultid="4021" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2677" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2678" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8108" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8109" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8110" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8111" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8112" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8113" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8114" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="8115" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="8116" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="8117" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1584" daytime="11:29" gender="F" number="35" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2709" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4624" />
                    <RANKING order="2" place="2" resultid="4618" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2710" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2962" />
                    <RANKING order="2" place="2" resultid="3107" />
                    <RANKING order="3" place="3" resultid="4636" />
                    <RANKING order="4" place="4" resultid="3981" />
                    <RANKING order="5" place="5" resultid="4773" />
                    <RANKING order="6" place="-1" resultid="4332" />
                    <RANKING order="7" place="-1" resultid="4611" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2711" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3971" />
                    <RANKING order="2" place="2" resultid="4825" />
                    <RANKING order="3" place="3" resultid="4077" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2712" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5762" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2713" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5005" />
                    <RANKING order="2" place="2" resultid="4734" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2714" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3667" />
                    <RANKING order="2" place="2" resultid="3114" />
                    <RANKING order="3" place="3" resultid="4702" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2715" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5392" />
                    <RANKING order="2" place="2" resultid="5099" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2716" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4553" />
                    <RANKING order="2" place="2" resultid="3452" />
                    <RANKING order="3" place="3" resultid="4451" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2717" agemax="64" agemin="60" name="Kat. H" />
                <AGEGROUP agegroupid="2718" agemax="69" agemin="65" name="Kat. I" />
                <AGEGROUP agegroupid="2719" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="2720" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4961" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2721" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="2722" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2723" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8159" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8160" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8161" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1569" daytime="11:04" gender="M" number="34" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2694" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4584" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2695" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3548" />
                    <RANKING order="2" place="2" resultid="5343" />
                    <RANKING order="3" place="3" resultid="2875" />
                    <RANKING order="4" place="4" resultid="5045" />
                    <RANKING order="5" place="5" resultid="5250" />
                    <RANKING order="6" place="6" resultid="3362" />
                    <RANKING order="7" place="7" resultid="3343" />
                    <RANKING order="8" place="8" resultid="3609" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2696" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5261" />
                    <RANKING order="2" place="2" resultid="2794" />
                    <RANKING order="3" place="3" resultid="2845" />
                    <RANKING order="4" place="4" resultid="4292" />
                    <RANKING order="5" place="5" resultid="4147" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2697" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4834" />
                    <RANKING order="2" place="2" resultid="3127" />
                    <RANKING order="3" place="3" resultid="5318" />
                    <RANKING order="4" place="4" resultid="3175" />
                    <RANKING order="5" place="5" resultid="4162" />
                    <RANKING order="6" place="6" resultid="4151" />
                    <RANKING order="7" place="7" resultid="4106" />
                    <RANKING order="8" place="-1" resultid="3921" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2698" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6413" />
                    <RANKING order="2" place="2" resultid="5350" />
                    <RANKING order="3" place="3" resultid="2216" />
                    <RANKING order="4" place="4" resultid="4918" />
                    <RANKING order="5" place="5" resultid="4927" />
                    <RANKING order="6" place="6" resultid="3962" />
                    <RANKING order="7" place="7" resultid="5221" />
                    <RANKING order="8" place="8" resultid="2153" />
                    <RANKING order="9" place="9" resultid="3309" />
                    <RANKING order="10" place="10" resultid="3081" />
                    <RANKING order="11" place="11" resultid="4053" />
                    <RANKING order="12" place="-1" resultid="3374" />
                    <RANKING order="13" place="-1" resultid="3394" />
                    <RANKING order="14" place="-1" resultid="3807" />
                    <RANKING order="15" place="-1" resultid="4747" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2699" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6417" />
                    <RANKING order="2" place="2" resultid="5311" />
                    <RANKING order="3" place="3" resultid="5446" />
                    <RANKING order="4" place="4" resultid="4905" />
                    <RANKING order="5" place="5" resultid="3635" />
                    <RANKING order="6" place="6" resultid="4040" />
                    <RANKING order="7" place="7" resultid="2857" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2700" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3943" />
                    <RANKING order="2" place="2" resultid="4715" />
                    <RANKING order="3" place="3" resultid="5483" />
                    <RANKING order="4" place="4" resultid="3787" />
                    <RANKING order="5" place="5" resultid="3683" />
                    <RANKING order="6" place="6" resultid="2839" />
                    <RANKING order="7" place="7" resultid="3578" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2701" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2767" />
                    <RANKING order="2" place="2" resultid="6036" />
                    <RANKING order="3" place="3" resultid="4952" />
                    <RANKING order="4" place="4" resultid="2760" />
                    <RANKING order="5" place="5" resultid="5307" />
                    <RANKING order="6" place="6" resultid="4857" />
                    <RANKING order="7" place="7" resultid="5034" />
                    <RANKING order="8" place="8" resultid="5421" />
                    <RANKING order="9" place="9" resultid="4193" />
                    <RANKING order="10" place="10" resultid="2175" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2702" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3571" />
                    <RANKING order="2" place="2" resultid="3404" />
                    <RANKING order="3" place="3" resultid="3006" />
                    <RANKING order="4" place="4" resultid="3487" />
                    <RANKING order="5" place="5" resultid="3757" />
                    <RANKING order="6" place="6" resultid="4741" />
                    <RANKING order="7" place="7" resultid="4405" />
                    <RANKING order="8" place="8" resultid="3855" />
                    <RANKING order="9" place="9" resultid="4817" />
                    <RANKING order="10" place="10" resultid="4071" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2703" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4993" />
                    <RANKING order="2" place="2" resultid="5025" />
                    <RANKING order="3" place="3" resultid="3411" />
                    <RANKING order="4" place="4" resultid="3652" />
                    <RANKING order="5" place="5" resultid="6024" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2704" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2113" />
                    <RANKING order="2" place="2" resultid="2189" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2705" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5127" />
                    <RANKING order="2" place="2" resultid="3429" />
                    <RANKING order="3" place="3" resultid="4431" />
                    <RANKING order="4" place="4" resultid="2776" />
                    <RANKING order="5" place="5" resultid="3933" />
                    <RANKING order="6" place="6" resultid="4026" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2706" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3384" />
                    <RANKING order="2" place="2" resultid="3184" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2707" agemax="89" agemin="85" name="Kat. M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4091" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2708" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8124" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8125" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8126" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8127" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8128" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8129" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="8130" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="8131" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="8132" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1554" daytime="10:45" gender="F" number="33" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2679" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4113" />
                    <RANKING order="2" place="2" resultid="3602" />
                    <RANKING order="3" place="3" resultid="3555" />
                    <RANKING order="4" place="-1" resultid="3595" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2680" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2934" />
                    <RANKING order="2" place="2" resultid="2787" />
                    <RANKING order="3" place="3" resultid="4610" />
                    <RANKING order="4" place="4" resultid="4772" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2681" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4824" />
                    <RANKING order="2" place="2" resultid="3976" />
                    <RANKING order="3" place="3" resultid="2923" />
                    <RANKING order="4" place="4" resultid="3493" />
                    <RANKING order="5" place="5" resultid="3513" />
                    <RANKING order="6" place="6" resultid="4543" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2682" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5409" />
                    <RANKING order="2" place="2" resultid="4513" />
                    <RANKING order="3" place="3" resultid="4875" />
                    <RANKING order="4" place="4" resultid="4884" />
                    <RANKING order="5" place="5" resultid="4782" />
                    <RANKING order="6" place="6" resultid="4098" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2683" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5143" />
                    <RANKING order="2" place="2" resultid="4998" />
                    <RANKING order="3" place="3" resultid="2950" />
                    <RANKING order="4" place="4" resultid="4733" />
                    <RANKING order="5" place="5" resultid="4202" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2684" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3879" />
                    <RANKING order="2" place="2" resultid="2752" />
                    <RANKING order="3" place="3" resultid="4267" />
                    <RANKING order="4" place="4" resultid="4683" />
                    <RANKING order="5" place="5" resultid="5180" />
                    <RANKING order="6" place="6" resultid="4048" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2685" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5391" />
                    <RANKING order="2" place="2" resultid="5069" />
                    <RANKING order="3" place="3" resultid="2862" />
                    <RANKING order="4" place="4" resultid="4567" />
                    <RANKING order="5" place="5" resultid="3674" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2686" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5281" />
                    <RANKING order="2" place="2" resultid="3937" />
                    <RANKING order="3" place="3" resultid="3054" />
                    <RANKING order="4" place="4" resultid="4460" />
                    <RANKING order="5" place="5" resultid="4450" />
                    <RANKING order="6" place="-1" resultid="3451" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2687" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5362" />
                    <RANKING order="2" place="2" resultid="5369" />
                    <RANKING order="3" place="3" resultid="4198" />
                    <RANKING order="4" place="4" resultid="3438" />
                    <RANKING order="5" place="5" resultid="2831" />
                    <RANKING order="6" place="6" resultid="5107" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2688" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3915" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2689" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5137" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2690" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5357" />
                    <RANKING order="2" place="2" resultid="4013" />
                    <RANKING order="3" place="3" resultid="2232" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2691" agemax="84" agemin="80" name="Kat. L">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3019" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2692" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2693" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8118" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8119" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8120" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8121" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8122" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8123" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1614" daytime="13:06" gender="X" number="37" order="9" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1629" agemax="119" agemin="100" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6005" />
                    <RANKING order="2" place="2" resultid="6007" />
                    <RANKING order="3" place="3" resultid="6099" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1630" agemax="159" agemin="120" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5071" />
                    <RANKING order="2" place="2" resultid="5229" />
                    <RANKING order="3" place="3" resultid="3160" />
                    <RANKING order="4" place="4" resultid="6006" />
                    <RANKING order="5" place="5" resultid="5226" />
                    <RANKING order="6" place="6" resultid="6100" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1631" agemax="199" agemin="160" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5466" />
                    <RANKING order="2" place="2" resultid="6004" />
                    <RANKING order="3" place="3" resultid="6170" />
                    <RANKING order="4" place="4" resultid="5181" />
                    <RANKING order="5" place="5" resultid="3721" />
                    <RANKING order="6" place="6" resultid="4835" />
                    <RANKING order="7" place="7" resultid="3161" />
                    <RANKING order="8" place="8" resultid="8169" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1632" agemax="239" agemin="200" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3951" />
                    <RANKING order="2" place="2" resultid="5465" />
                    <RANKING order="3" place="3" resultid="2761" />
                    <RANKING order="4" place="4" resultid="5319" />
                    <RANKING order="5" place="5" resultid="3759" />
                    <RANKING order="6" place="-1" resultid="4474" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1633" agemax="279" agemin="240" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5072" />
                    <RANKING order="2" place="2" resultid="5464" />
                    <RANKING order="3" place="3" resultid="3952" />
                    <RANKING order="4" place="-1" resultid="3455" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1634" agemax="-1" agemin="280" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3454" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8133" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8134" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8135" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1524" daytime="10:16" gender="F" number="31" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2649" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4623" />
                    <RANKING order="2" place="2" resultid="4671" />
                    <RANKING order="3" place="3" resultid="4058" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2650" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5040" />
                    <RANKING order="2" place="2" resultid="3768" />
                    <RANKING order="3" place="3" resultid="4665" />
                    <RANKING order="4" place="4" resultid="3988" />
                    <RANKING order="5" place="5" resultid="4536" />
                    <RANKING order="6" place="6" resultid="2928" />
                    <RANKING order="7" place="7" resultid="5242" />
                    <RANKING order="8" place="-1" resultid="2939" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2651" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4076" />
                    <RANKING order="2" place="2" resultid="3319" />
                    <RANKING order="3" place="3" resultid="5194" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2652" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4874" />
                    <RANKING order="2" place="2" resultid="3121" />
                    <RANKING order="3" place="3" resultid="2134" />
                    <RANKING order="4" place="4" resultid="4911" />
                    <RANKING order="5" place="5" resultid="4883" />
                    <RANKING order="6" place="6" resultid="4781" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2653" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5004" />
                    <RANKING order="2" place="2" resultid="4688" />
                    <RANKING order="3" place="3" resultid="5397" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2654" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5174" />
                    <RANKING order="2" place="2" resultid="3878" />
                    <RANKING order="3" place="3" resultid="4866" />
                    <RANKING order="4" place="4" resultid="4047" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2655" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5013" />
                    <RANKING order="2" place="2" resultid="3400" />
                    <RANKING order="3" place="3" resultid="3696" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2656" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4552" />
                    <RANKING order="2" place="2" resultid="2748" />
                    <RANKING order="3" place="3" resultid="5286" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2657" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3420" />
                    <RANKING order="2" place="2" resultid="3628" />
                    <RANKING order="3" place="3" resultid="5106" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2658" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2808" />
                    <RANKING order="2" place="2" resultid="5276" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2659" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2660" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4960" />
                    <RANKING order="2" place="2" resultid="2231" />
                    <RANKING order="3" place="3" resultid="4006" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2661" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="2662" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2663" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8103" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8104" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8105" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8106" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8107" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1599" daytime="12:03" gender="M" number="36" order="8" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2724" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3711" />
                    <RANKING order="2" place="2" resultid="4314" />
                    <RANKING order="3" place="3" resultid="3146" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2725" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3011" />
                    <RANKING order="2" place="2" resultid="4185" />
                    <RANKING order="3" place="3" resultid="5344" />
                    <RANKING order="4" place="4" resultid="4652" />
                    <RANKING order="5" place="5" resultid="3610" />
                    <RANKING order="6" place="-1" resultid="2886" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2726" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4645" />
                    <RANKING order="2" place="2" resultid="2795" />
                    <RANKING order="3" place="3" resultid="4790" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2727" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3662" />
                    <RANKING order="2" place="2" resultid="3777" />
                    <RANKING order="3" place="3" resultid="3071" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2728" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4237" />
                    <RANKING order="2" place="2" resultid="5351" />
                    <RANKING order="3" place="3" resultid="3141" />
                    <RANKING order="4" place="4" resultid="3963" />
                    <RANKING order="5" place="5" resultid="3866" />
                    <RANKING order="6" place="6" resultid="4253" />
                    <RANKING order="7" place="7" resultid="4892" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2729" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4529" />
                    <RANKING order="2" place="2" resultid="4066" />
                    <RANKING order="3" place="3" resultid="4041" />
                    <RANKING order="4" place="4" resultid="4423" />
                    <RANKING order="5" place="5" resultid="2858" />
                    <RANKING order="6" place="-1" resultid="4522" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2730" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5085" />
                    <RANKING order="2" place="2" resultid="5432" />
                    <RANKING order="3" place="3" resultid="3157" />
                    <RANKING order="4" place="4" resultid="4730" />
                    <RANKING order="5" place="5" resultid="5751" />
                    <RANKING order="6" place="6" resultid="3689" />
                    <RANKING order="7" place="7" resultid="2840" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2731" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3089" />
                    <RANKING order="2" place="2" resultid="4259" />
                    <RANKING order="3" place="3" resultid="4696" />
                    <RANKING order="4" place="4" resultid="3737" />
                    <RANKING order="5" place="5" resultid="2169" />
                    <RANKING order="6" place="-1" resultid="2162" />
                    <RANKING order="7" place="-1" resultid="4561" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2732" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3503" />
                    <RANKING order="2" place="2" resultid="5298" />
                    <RANKING order="3" place="3" resultid="4414" />
                    <RANKING order="4" place="4" resultid="3278" />
                    <RANKING order="5" place="5" resultid="3758" />
                    <RANKING order="6" place="6" resultid="4765" />
                    <RANKING order="7" place="7" resultid="4406" />
                    <RANKING order="8" place="8" resultid="3316" />
                    <RANKING order="9" place="-1" resultid="3524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2733" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4244" />
                    <RANKING order="2" place="2" resultid="3793" />
                    <RANKING order="3" place="3" resultid="3412" />
                    <RANKING order="4" place="4" resultid="4976" />
                    <RANKING order="5" place="5" resultid="3906" />
                    <RANKING order="6" place="6" resultid="4373" />
                    <RANKING order="7" place="7" resultid="4804" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2734" agemax="74" agemin="70" name="Kat. J">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2122" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2735" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4432" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2736" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="2737" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2738" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8162" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8163" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8164" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8165" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8166" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8167" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1493" daytime="09:00" gender="F" number="29" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2619" agemax="24" agemin="20" name="Kat. 0">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4112" />
                    <RANKING order="2" place="2" resultid="5267" />
                    <RANKING order="3" place="3" resultid="2852" />
                    <RANKING order="4" place="4" resultid="3554" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2620" agemax="29" agemin="25" name="Kat. A">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3767" />
                    <RANKING order="2" place="2" resultid="2961" />
                    <RANKING order="3" place="3" resultid="2933" />
                    <RANKING order="4" place="4" resultid="5213" />
                    <RANKING order="5" place="5" resultid="4600" />
                    <RANKING order="6" place="6" resultid="5241" />
                    <RANKING order="7" place="7" resultid="5091" />
                    <RANKING order="8" place="8" resultid="3062" />
                    <RANKING order="9" place="-1" resultid="4331" />
                    <RANKING order="10" place="-1" resultid="4664" />
                    <RANKING order="11" place="-1" resultid="5039" />
                    <RANKING order="12" place="-1" resultid="5414" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2621" agemax="34" agemin="30" name="Kat. B">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3100" />
                    <RANKING order="2" place="2" resultid="3096" />
                    <RANKING order="3" place="3" resultid="3512" />
                    <RANKING order="4" place="4" resultid="4542" />
                    <RANKING order="5" place="5" resultid="2944" />
                    <RANKING order="6" place="6" resultid="3889" />
                    <RANKING order="7" place="-1" resultid="4590" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2622" agemax="39" agemin="35" name="Kat. C">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5761" />
                    <RANKING order="2" place="2" resultid="4910" />
                    <RANKING order="3" place="3" resultid="4097" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2623" agemax="44" agemin="40" name="Kat. D">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5404" />
                    <RANKING order="2" place="2" resultid="4117" />
                    <RANKING order="3" place="3" resultid="3742" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2624" agemax="49" agemin="45" name="Kat. E">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3666" />
                    <RANKING order="2" place="2" resultid="3113" />
                    <RANKING order="3" place="3" resultid="4682" />
                    <RANKING order="4" place="4" resultid="5179" />
                    <RANKING order="5" place="5" resultid="4266" />
                    <RANKING order="6" place="6" resultid="3045" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2625" agemax="54" agemin="50" name="Kat. F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5380" />
                    <RANKING order="2" place="2" resultid="3291" />
                    <RANKING order="3" place="3" resultid="3695" />
                    <RANKING order="4" place="4" resultid="3399" />
                    <RANKING order="5" place="5" resultid="5098" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2626" agemax="59" agemin="55" name="Kat. G">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5376" />
                    <RANKING order="2" place="2" resultid="4501" />
                    <RANKING order="3" place="3" resultid="3884" />
                    <RANKING order="4" place="4" resultid="4459" />
                    <RANKING order="5" place="5" resultid="5756" />
                    <RANKING order="6" place="6" resultid="3749" />
                    <RANKING order="7" place="-1" resultid="3053" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2627" agemax="64" agemin="60" name="Kat. H">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3437" />
                    <RANKING order="2" place="2" resultid="3627" />
                    <RANKING order="3" place="3" resultid="2830" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2628" agemax="69" agemin="65" name="Kat. I">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5275" />
                    <RANKING order="2" place="2" resultid="5149" />
                    <RANKING order="3" place="3" resultid="2893" />
                    <RANKING order="4" place="4" resultid="3914" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2629" agemax="74" agemin="70" name="Kat. J" />
                <AGEGROUP agegroupid="2630" agemax="79" agemin="75" name="Kat. K">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4005" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2631" agemax="84" agemin="80" name="Kat. L" />
                <AGEGROUP agegroupid="2632" agemax="89" agemin="85" name="Kat. M" />
                <AGEGROUP agegroupid="2633" agemax="94" agemin="90" name="Kat. N" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="8087" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="8088" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="8089" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="8090" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="8091" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="8092" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" nation="POL" clubid="2135" name="Andrzej Waszkewicz Sports Project" shortname="Andrzej Waszkewicz Sports Proj">
          <CONTACT email="info@swim.by" internet="www.swim.by" name="Swim Academy" />
          <ATHLETES>
            <ATHLETE birthdate="1983-05-01" firstname="Andrzej" gender="M" lastname="Waszkewicz" nation="POL" athleteid="2136">
              <RESULTS>
                <RESULT eventid="1105" points="884" reactiontime="+91" swimtime="00:00:26.07" resultid="2137" heatid="7972" lane="5" entrytime="00:00:25.20" entrycourse="LCM" />
                <RESULT eventid="1372" points="823" reactiontime="+90" swimtime="00:00:24.81" resultid="2138" heatid="8065" lane="3" entrytime="00:00:24.20" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3033" name="Aquapark Wrocław">
          <CONTACT name="Stasiaczek" phone="792883772" />
          <ATHLETES>
            <ATHLETE birthdate="1960-05-11" firstname="Joanna" gender="F" lastname="Krowicka" nation="POL" athleteid="3046">
              <RESULTS>
                <RESULT eventid="1058" points="464" reactiontime="+75" swimtime="00:03:44.25" resultid="3047" heatid="7942" lane="8" entrytime="00:03:52.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.18" />
                    <SPLIT distance="100" swimtime="00:01:53.97" />
                    <SPLIT distance="150" swimtime="00:02:53.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="385" reactiontime="+81" swimtime="00:00:47.59" resultid="3048" heatid="7956" lane="7" entrytime="00:00:46.02" />
                <RESULT eventid="1181" points="473" reactiontime="+82" swimtime="00:01:28.75" resultid="3049" heatid="7975" lane="6" entrytime="00:01:24.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="517" reactiontime="+76" swimtime="00:00:47.75" resultid="3050" heatid="7996" lane="3" entrytime="00:00:46.38" />
                <RESULT eventid="1357" points="563" reactiontime="+66" swimtime="00:00:37.38" resultid="3051" heatid="8046" lane="8" entrytime="00:00:37.73" />
                <RESULT eventid="1417" points="504" reactiontime="+69" swimtime="00:07:13.75" resultid="3052" heatid="8149" lane="2" entrytime="00:07:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.29" />
                    <SPLIT distance="100" swimtime="00:01:37.97" />
                    <SPLIT distance="150" swimtime="00:02:34.42" />
                    <SPLIT distance="200" swimtime="00:03:30.87" />
                    <SPLIT distance="250" swimtime="00:04:28.51" />
                    <SPLIT distance="300" swimtime="00:05:26.21" />
                    <SPLIT distance="350" swimtime="00:06:23.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" status="DNS" swimtime="00:00:00.00" resultid="3053" heatid="8088" lane="4" entrytime="00:03:24.00" />
                <RESULT eventid="1554" points="596" swimtime="00:01:41.48" resultid="3054" heatid="8121" lane="9" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-07-24" firstname="Tomasz" gender="M" lastname="Olas" nation="POL" athleteid="3037">
              <RESULTS>
                <RESULT eventid="1198" points="311" reactiontime="+76" swimtime="00:01:16.69" resultid="3038" heatid="7984" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="360" reactiontime="+73" swimtime="00:00:33.07" resultid="3039" heatid="8054" lane="0" entrytime="00:00:37.00" />
                <RESULT eventid="1509" points="281" reactiontime="+96" swimtime="00:02:56.51" resultid="3040" heatid="8098" lane="1" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.72" />
                    <SPLIT distance="100" swimtime="00:01:22.52" />
                    <SPLIT distance="150" swimtime="00:02:09.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-04-23" firstname="Agata" gender="F" lastname="Sobczak" nation="POL" athleteid="3055">
              <RESULTS>
                <RESULT eventid="1090" points="213" reactiontime="+106" swimtime="00:00:47.36" resultid="3056" heatid="7957" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1150" points="289" reactiontime="+98" swimtime="00:28:12.89" resultid="3057" heatid="8142" lane="5" entrytime="00:22:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.56" />
                    <SPLIT distance="100" swimtime="00:01:39.00" />
                    <SPLIT distance="150" swimtime="00:02:33.87" />
                    <SPLIT distance="200" swimtime="00:03:28.63" />
                    <SPLIT distance="250" swimtime="00:04:24.88" />
                    <SPLIT distance="300" swimtime="00:05:21.39" />
                    <SPLIT distance="350" swimtime="00:06:18.34" />
                    <SPLIT distance="400" swimtime="00:07:14.94" />
                    <SPLIT distance="450" swimtime="00:08:11.17" />
                    <SPLIT distance="500" swimtime="00:09:07.82" />
                    <SPLIT distance="550" swimtime="00:10:04.21" />
                    <SPLIT distance="600" swimtime="00:11:01.48" />
                    <SPLIT distance="650" swimtime="00:11:58.47" />
                    <SPLIT distance="700" swimtime="00:12:55.04" />
                    <SPLIT distance="750" swimtime="00:13:51.93" />
                    <SPLIT distance="800" swimtime="00:14:48.72" />
                    <SPLIT distance="850" swimtime="00:15:47.32" />
                    <SPLIT distance="900" swimtime="00:16:45.63" />
                    <SPLIT distance="950" swimtime="00:17:43.84" />
                    <SPLIT distance="1000" swimtime="00:18:39.17" />
                    <SPLIT distance="1050" swimtime="00:19:37.30" />
                    <SPLIT distance="1100" swimtime="00:20:35.81" />
                    <SPLIT distance="1150" swimtime="00:21:32.98" />
                    <SPLIT distance="1200" swimtime="00:22:30.33" />
                    <SPLIT distance="1250" swimtime="00:23:27.88" />
                    <SPLIT distance="1300" swimtime="00:24:25.05" />
                    <SPLIT distance="1350" swimtime="00:25:22.98" />
                    <SPLIT distance="1400" swimtime="00:26:20.15" />
                    <SPLIT distance="1450" swimtime="00:27:17.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="243" reactiontime="+102" swimtime="00:01:34.04" resultid="3058" heatid="7975" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1243" points="194" reactiontime="+106" swimtime="00:04:12.96" resultid="3059" heatid="8012" lane="6" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.33" />
                    <SPLIT distance="100" swimtime="00:01:58.80" />
                    <SPLIT distance="150" swimtime="00:03:05.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="262" reactiontime="+101" swimtime="00:07:06.49" resultid="3060" heatid="8147" lane="0" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.10" />
                    <SPLIT distance="100" swimtime="00:01:40.04" />
                    <SPLIT distance="150" swimtime="00:02:34.22" />
                    <SPLIT distance="200" swimtime="00:03:29.37" />
                    <SPLIT distance="250" swimtime="00:04:24.63" />
                    <SPLIT distance="300" swimtime="00:05:19.01" />
                    <SPLIT distance="350" swimtime="00:06:13.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="178" reactiontime="+100" swimtime="00:01:53.91" resultid="3061" heatid="8078" lane="6" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="243" reactiontime="+100" swimtime="00:03:26.51" resultid="3062" heatid="8090" lane="0" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.82" />
                    <SPLIT distance="100" swimtime="00:01:40.61" />
                    <SPLIT distance="150" swimtime="00:02:34.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-12-31" firstname="Agata" gender="F" lastname="Szydło" nation="POL" athleteid="3041">
              <RESULTS>
                <RESULT eventid="1120" points="284" reactiontime="+101" swimtime="00:14:42.44" resultid="3042" heatid="8137" lane="1" entrytime="00:14:44.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.46" />
                    <SPLIT distance="100" swimtime="00:01:43.20" />
                    <SPLIT distance="150" swimtime="00:02:38.91" />
                    <SPLIT distance="200" swimtime="00:03:35.45" />
                    <SPLIT distance="250" swimtime="00:04:31.73" />
                    <SPLIT distance="300" swimtime="00:05:27.67" />
                    <SPLIT distance="350" swimtime="00:06:24.21" />
                    <SPLIT distance="400" swimtime="00:07:20.52" />
                    <SPLIT distance="450" swimtime="00:08:16.44" />
                    <SPLIT distance="500" swimtime="00:09:12.13" />
                    <SPLIT distance="550" swimtime="00:10:08.19" />
                    <SPLIT distance="600" swimtime="00:11:04.12" />
                    <SPLIT distance="650" swimtime="00:11:59.79" />
                    <SPLIT distance="700" swimtime="00:12:55.33" />
                    <SPLIT distance="750" swimtime="00:13:50.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="329" reactiontime="+80" swimtime="00:00:52.99" resultid="3043" heatid="7995" lane="6" entrytime="00:00:55.76" />
                <RESULT eventid="1387" points="360" swimtime="00:04:00.11" resultid="3044" heatid="8068" lane="9" entrytime="00:03:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.26" />
                    <SPLIT distance="100" swimtime="00:01:55.06" />
                    <SPLIT distance="150" swimtime="00:02:57.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="271" reactiontime="+85" swimtime="00:03:29.76" resultid="3045" heatid="8089" lane="9" entrytime="00:03:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.97" />
                    <SPLIT distance="100" swimtime="00:01:39.71" />
                    <SPLIT distance="150" swimtime="00:02:35.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-07" firstname="Radosław" gender="M" lastname="Stefurak" nation="POL" athleteid="3075">
              <RESULTS>
                <RESULT eventid="1198" points="367" reactiontime="+80" swimtime="00:01:15.83" resultid="3076" heatid="7983" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="470" reactiontime="+85" swimtime="00:00:39.24" resultid="3077" heatid="8005" lane="2" entrytime="00:00:39.00" />
                <RESULT eventid="1402" points="473" reactiontime="+91" swimtime="00:03:13.58" resultid="3079" heatid="8075" lane="6" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.37" />
                    <SPLIT distance="100" swimtime="00:01:32.22" />
                    <SPLIT distance="150" swimtime="00:02:22.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="455" reactiontime="+84" swimtime="00:01:29.35" resultid="3081" heatid="8128" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-02-15" firstname="Wojciech" gender="M" lastname="Sobczak" nation="POL" athleteid="3063">
              <RESULTS>
                <RESULT eventid="1075" points="303" reactiontime="+111" swimtime="00:03:21.12" resultid="3064" heatid="7949" lane="0" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.58" />
                    <SPLIT distance="100" swimtime="00:01:37.84" />
                    <SPLIT distance="150" swimtime="00:02:38.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="341" reactiontime="+111" swimtime="00:12:45.99" resultid="3065" heatid="8140" lane="3" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.13" />
                    <SPLIT distance="100" swimtime="00:01:26.07" />
                    <SPLIT distance="150" swimtime="00:02:13.89" />
                    <SPLIT distance="200" swimtime="00:03:01.39" />
                    <SPLIT distance="250" swimtime="00:03:49.45" />
                    <SPLIT distance="300" swimtime="00:04:39.56" />
                    <SPLIT distance="350" swimtime="00:05:28.03" />
                    <SPLIT distance="400" swimtime="00:06:17.14" />
                    <SPLIT distance="450" swimtime="00:07:05.80" />
                    <SPLIT distance="500" swimtime="00:07:55.35" />
                    <SPLIT distance="550" swimtime="00:08:45.11" />
                    <SPLIT distance="600" swimtime="00:09:35.23" />
                    <SPLIT distance="650" swimtime="00:10:24.52" />
                    <SPLIT distance="700" swimtime="00:11:13.68" />
                    <SPLIT distance="750" swimtime="00:12:00.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="194" reactiontime="+109" swimtime="00:03:52.18" resultid="3066" heatid="8016" lane="9" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.49" />
                    <SPLIT distance="100" swimtime="00:01:47.24" />
                    <SPLIT distance="150" swimtime="00:02:49.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="268" reactiontime="+84" swimtime="00:03:27.08" resultid="3067" heatid="8025" lane="7" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.18" />
                    <SPLIT distance="100" swimtime="00:01:41.28" />
                    <SPLIT distance="150" swimtime="00:02:35.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="320" reactiontime="+101" swimtime="00:03:41.18" resultid="3068" heatid="8074" lane="1" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.82" />
                    <SPLIT distance="100" swimtime="00:01:46.82" />
                    <SPLIT distance="150" swimtime="00:02:46.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="183" reactiontime="+105" swimtime="00:01:42.43" resultid="3069" heatid="8082" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="354" reactiontime="+105" swimtime="00:02:43.39" resultid="3070" heatid="8098" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.34" />
                    <SPLIT distance="100" swimtime="00:01:15.72" />
                    <SPLIT distance="150" swimtime="00:01:59.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="314" reactiontime="+117" swimtime="00:07:09.53" resultid="3071" heatid="8165" lane="9" entrytime="00:07:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.60" />
                    <SPLIT distance="100" swimtime="00:01:51.54" />
                    <SPLIT distance="150" swimtime="00:02:46.34" />
                    <SPLIT distance="200" swimtime="00:03:41.00" />
                    <SPLIT distance="250" swimtime="00:04:44.17" />
                    <SPLIT distance="300" swimtime="00:05:46.31" />
                    <SPLIT distance="350" swimtime="00:06:27.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-07-21" firstname="Mateusz" gender="M" lastname="Dudek" nation="POL" athleteid="3072">
              <RESULTS>
                <RESULT eventid="1228" points="759" reactiontime="+75" swimtime="00:00:32.12" resultid="3073" heatid="8010" lane="2" entrytime="00:00:31.50" />
                <RESULT eventid="1402" points="725" reactiontime="+75" swimtime="00:02:42.86" resultid="3074" heatid="8077" lane="2" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                    <SPLIT distance="100" swimtime="00:01:17.92" />
                    <SPLIT distance="150" swimtime="00:01:59.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3082" name="Aquasfera Masters Olsztyn">
          <CONTACT email="gozdzik@uwm.edu.pl" name="Goździejewska Anna" />
          <ATHLETES>
            <ATHLETE birthdate="1992-08-16" firstname="Paweł" gender="M" lastname="Szczuka" nation="POL" athleteid="3142">
              <RESULTS>
                <RESULT eventid="1075" points="682" reactiontime="+71" swimtime="00:02:27.22" resultid="3143" heatid="7952" lane="4" entrytime="00:02:30.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.69" />
                    <SPLIT distance="100" swimtime="00:01:08.95" />
                    <SPLIT distance="150" swimtime="00:01:51.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="704" reactiontime="+72" swimtime="00:00:32.81" resultid="3144" heatid="8010" lane="9" entrytime="00:00:32.80" />
                <RESULT eventid="1372" points="683" reactiontime="+75" swimtime="00:00:26.14" resultid="3145" heatid="8064" lane="8" entrytime="00:00:26.10" />
                <RESULT eventid="1599" points="646" reactiontime="+78" swimtime="00:05:23.54" resultid="3146" heatid="8162" lane="2" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                    <SPLIT distance="100" swimtime="00:01:09.75" />
                    <SPLIT distance="150" swimtime="00:01:52.81" />
                    <SPLIT distance="200" swimtime="00:02:36.85" />
                    <SPLIT distance="250" swimtime="00:03:22.02" />
                    <SPLIT distance="300" swimtime="00:04:08.86" />
                    <SPLIT distance="350" swimtime="00:04:46.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-04-24" firstname="Przemysław" gender="M" lastname="Bielski" nation="POL" athleteid="3128">
              <RESULTS>
                <RESULT eventid="1105" points="479" reactiontime="+76" swimtime="00:00:33.08" resultid="3129" heatid="7966" lane="8" entrytime="00:00:34.50" />
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="3130" heatid="7987" lane="7" entrytime="00:01:06.89" />
                <RESULT eventid="1372" status="DNS" swimtime="00:00:00.00" resultid="3131" heatid="8056" lane="4" entrytime="00:00:30.67" />
                <RESULT eventid="1509" points="474" reactiontime="+92" swimtime="00:02:31.92" resultid="3133" heatid="8099" lane="0" entrytime="00:02:33.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                    <SPLIT distance="100" swimtime="00:01:11.62" />
                    <SPLIT distance="150" swimtime="00:01:51.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-02-15" firstname="Jowita" gender="F" lastname="Kucharska" nation="POL" athleteid="3115">
              <RESULTS>
                <RESULT eventid="1058" points="572" reactiontime="+93" swimtime="00:02:59.64" resultid="3116" heatid="7943" lane="7" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.61" />
                    <SPLIT distance="100" swimtime="00:01:25.14" />
                    <SPLIT distance="150" swimtime="00:02:20.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="588" reactiontime="+86" swimtime="00:00:35.46" resultid="3117" heatid="7958" lane="5" entrytime="00:00:36.00" />
                <RESULT eventid="1273" points="507" reactiontime="+76" swimtime="00:03:06.70" resultid="3118" heatid="8020" lane="8" entrytime="00:03:07.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.77" />
                    <SPLIT distance="100" swimtime="00:01:31.89" />
                    <SPLIT distance="150" swimtime="00:02:20.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="572" reactiontime="+76" swimtime="00:01:24.14" resultid="3119" heatid="8034" lane="2" entrytime="00:01:24.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="615" reactiontime="+81" swimtime="00:00:32.27" resultid="3120" heatid="8048" lane="8" entrytime="00:00:33.00" />
                <RESULT eventid="1524" points="553" reactiontime="+76" swimtime="00:00:39.10" resultid="3121" heatid="8105" lane="5" entrytime="00:00:39.71" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-17" firstname="Anna" gender="F" lastname="Piekut" nation="POL" athleteid="3101">
              <RESULTS>
                <RESULT eventid="1058" points="523" reactiontime="+69" swimtime="00:03:00.32" resultid="3102" heatid="7944" lane="8" entrytime="00:02:55.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                    <SPLIT distance="100" swimtime="00:01:22.84" />
                    <SPLIT distance="150" swimtime="00:02:17.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="547" reactiontime="+77" swimtime="00:00:34.59" resultid="3103" heatid="7959" lane="3" entrytime="00:00:34.40" />
                <RESULT eventid="1243" points="635" reactiontime="+79" swimtime="00:02:50.49" resultid="3104" heatid="8012" lane="5" entrytime="00:02:46.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.42" />
                    <SPLIT distance="100" swimtime="00:01:20.61" />
                    <SPLIT distance="150" swimtime="00:02:05.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="502" reactiontime="+76" swimtime="00:00:34.02" resultid="3105" heatid="8047" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="1447" points="566" reactiontime="+82" swimtime="00:01:17.55" resultid="3106" heatid="8080" lane="7" entrytime="00:01:16.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1584" points="559" reactiontime="+85" swimtime="00:06:18.50" resultid="3107" heatid="8159" lane="7" entrytime="00:06:10.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.87" />
                    <SPLIT distance="100" swimtime="00:01:21.93" />
                    <SPLIT distance="150" swimtime="00:02:12.57" />
                    <SPLIT distance="200" swimtime="00:03:01.30" />
                    <SPLIT distance="250" swimtime="00:03:55.32" />
                    <SPLIT distance="300" swimtime="00:04:50.12" />
                    <SPLIT distance="350" swimtime="00:05:34.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-13" firstname="Michał" gender="M" lastname="Kozikowski" nation="POL" athleteid="3122">
              <RESULTS>
                <RESULT eventid="1075" points="683" reactiontime="+73" swimtime="00:02:33.40" resultid="3123" heatid="7952" lane="7" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.13" />
                    <SPLIT distance="100" swimtime="00:01:12.36" />
                    <SPLIT distance="150" swimtime="00:01:55.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="599" reactiontime="+78" swimtime="00:01:01.65" resultid="3124" heatid="7988" lane="7" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="651" reactiontime="+76" swimtime="00:00:27.14" resultid="3125" heatid="8051" lane="3" />
                <RESULT eventid="1402" points="761" reactiontime="+75" swimtime="00:02:45.77" resultid="3126" heatid="8077" lane="7" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.50" />
                    <SPLIT distance="100" swimtime="00:01:20.38" />
                    <SPLIT distance="150" swimtime="00:02:03.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="694" reactiontime="+70" swimtime="00:01:15.04" resultid="3127" heatid="8131" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-03-18" firstname="Anna" gender="F" lastname="Goździejewska" nation="POL" athleteid="3108">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1150" points="759" reactiontime="+91" swimtime="00:22:34.77" resultid="3109" heatid="8142" lane="3" entrytime="00:23:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.71" />
                    <SPLIT distance="100" swimtime="00:01:25.95" />
                    <SPLIT distance="150" swimtime="00:02:11.20" />
                    <SPLIT distance="200" swimtime="00:02:57.10" />
                    <SPLIT distance="250" swimtime="00:03:42.62" />
                    <SPLIT distance="300" swimtime="00:04:28.55" />
                    <SPLIT distance="350" swimtime="00:05:13.44" />
                    <SPLIT distance="400" swimtime="00:05:58.71" />
                    <SPLIT distance="450" swimtime="00:06:43.70" />
                    <SPLIT distance="500" swimtime="00:07:28.70" />
                    <SPLIT distance="550" swimtime="00:08:13.89" />
                    <SPLIT distance="600" swimtime="00:08:59.29" />
                    <SPLIT distance="650" swimtime="00:09:44.80" />
                    <SPLIT distance="700" swimtime="00:10:30.00" />
                    <SPLIT distance="750" swimtime="00:11:15.48" />
                    <SPLIT distance="800" swimtime="00:12:01.16" />
                    <SPLIT distance="850" swimtime="00:12:46.56" />
                    <SPLIT distance="900" swimtime="00:13:32.10" />
                    <SPLIT distance="950" swimtime="00:14:17.11" />
                    <SPLIT distance="1000" swimtime="00:15:02.94" />
                    <SPLIT distance="1050" swimtime="00:15:48.16" />
                    <SPLIT distance="1100" swimtime="00:16:33.51" />
                    <SPLIT distance="1150" swimtime="00:17:18.80" />
                    <SPLIT distance="1200" swimtime="00:18:04.58" />
                    <SPLIT distance="1250" swimtime="00:18:50.61" />
                    <SPLIT distance="1300" swimtime="00:19:36.08" />
                    <SPLIT distance="1350" swimtime="00:20:21.37" />
                    <SPLIT distance="1400" swimtime="00:21:06.64" />
                    <SPLIT distance="1450" swimtime="00:21:51.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="604" reactiontime="+77" swimtime="00:01:14.17" resultid="3110" heatid="7977" lane="9" entrytime="00:01:16.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1387" points="510" reactiontime="+86" swimtime="00:03:33.84" resultid="3111" heatid="8068" lane="7" entrytime="00:03:40.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.94" />
                    <SPLIT distance="100" swimtime="00:01:44.47" />
                    <SPLIT distance="150" swimtime="00:02:38.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="515" reactiontime="+88" swimtime="00:05:54.65" resultid="3112" heatid="8148" lane="3" entrytime="00:06:00.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.94" />
                    <SPLIT distance="100" swimtime="00:01:24.61" />
                    <SPLIT distance="150" swimtime="00:02:09.97" />
                    <SPLIT distance="200" swimtime="00:02:55.19" />
                    <SPLIT distance="250" swimtime="00:03:40.03" />
                    <SPLIT distance="300" swimtime="00:04:25.36" />
                    <SPLIT distance="350" swimtime="00:05:10.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="587" reactiontime="+89" swimtime="00:02:42.29" resultid="3113" heatid="8090" lane="3" entrytime="00:02:48.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.20" />
                    <SPLIT distance="100" swimtime="00:01:18.95" />
                    <SPLIT distance="150" swimtime="00:02:01.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1584" points="487" reactiontime="+92" swimtime="00:07:02.64" resultid="3114" heatid="8160" lane="8" entrytime="00:07:05.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.87" />
                    <SPLIT distance="100" swimtime="00:01:44.30" />
                    <SPLIT distance="150" swimtime="00:02:39.37" />
                    <SPLIT distance="200" swimtime="00:03:34.15" />
                    <SPLIT distance="250" swimtime="00:04:31.66" />
                    <SPLIT distance="300" swimtime="00:05:28.96" />
                    <SPLIT distance="350" swimtime="00:06:16.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-01-29" firstname="Mariusz" gender="M" lastname="Gabiec" nation="POL" athleteid="3083">
              <RESULTS>
                <RESULT eventid="1075" points="817" reactiontime="+82" swimtime="00:02:45.79" resultid="3084" heatid="7947" lane="1" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.96" />
                    <SPLIT distance="100" swimtime="00:01:17.13" />
                    <SPLIT distance="150" swimtime="00:02:07.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="783" reactiontime="+78" swimtime="00:00:30.95" resultid="3085" heatid="7968" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="1258" points="686" reactiontime="+83" swimtime="00:02:55.86" resultid="3086" heatid="8016" lane="2" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                    <SPLIT distance="100" swimtime="00:01:16.14" />
                    <SPLIT distance="150" swimtime="00:02:02.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="826" reactiontime="+77" swimtime="00:05:14.40" resultid="3087" heatid="8152" lane="0" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                    <SPLIT distance="100" swimtime="00:01:17.82" />
                    <SPLIT distance="150" swimtime="00:01:57.79" />
                    <SPLIT distance="200" swimtime="00:02:37.82" />
                    <SPLIT distance="250" swimtime="00:03:17.75" />
                    <SPLIT distance="300" swimtime="00:03:57.63" />
                    <SPLIT distance="350" swimtime="00:04:37.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="840" reactiontime="+84" swimtime="00:00:34.43" resultid="3088" heatid="8110" lane="7" entrytime="00:00:48.00" />
                <RESULT comment="Rekord Polski Masters" eventid="1599" points="732" reactiontime="+78" swimtime="00:06:09.16" resultid="3089" heatid="8163" lane="8" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.90" />
                    <SPLIT distance="100" swimtime="00:01:23.99" />
                    <SPLIT distance="150" swimtime="00:02:10.93" />
                    <SPLIT distance="200" swimtime="00:02:56.97" />
                    <SPLIT distance="250" swimtime="00:03:52.97" />
                    <SPLIT distance="300" swimtime="00:04:49.90" />
                    <SPLIT distance="350" swimtime="00:05:30.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-26" firstname="Aleksandra" gender="F" lastname="Przybysz" nation="POL" athleteid="3090">
              <RESULTS>
                <RESULT eventid="1120" points="414" reactiontime="+76" swimtime="00:12:49.40" resultid="3091" heatid="8136" lane="9" entrytime="00:12:21.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.89" />
                    <SPLIT distance="100" swimtime="00:01:25.36" />
                    <SPLIT distance="150" swimtime="00:02:11.64" />
                    <SPLIT distance="200" swimtime="00:02:58.22" />
                    <SPLIT distance="250" swimtime="00:03:45.64" />
                    <SPLIT distance="300" swimtime="00:04:32.90" />
                    <SPLIT distance="350" swimtime="00:05:20.96" />
                    <SPLIT distance="400" swimtime="00:06:09.69" />
                    <SPLIT distance="450" swimtime="00:06:58.55" />
                    <SPLIT distance="500" swimtime="00:07:47.92" />
                    <SPLIT distance="550" swimtime="00:08:38.41" />
                    <SPLIT distance="600" swimtime="00:09:28.88" />
                    <SPLIT distance="650" swimtime="00:10:19.98" />
                    <SPLIT distance="700" swimtime="00:11:10.40" />
                    <SPLIT distance="750" swimtime="00:12:00.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="443" reactiontime="+77" swimtime="00:01:17.30" resultid="3092" heatid="7976" lane="3" entrytime="00:01:17.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1243" points="374" reactiontime="+94" swimtime="00:03:23.54" resultid="3093" heatid="8012" lane="7" entrytime="00:03:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.26" />
                    <SPLIT distance="100" swimtime="00:01:35.37" />
                    <SPLIT distance="150" swimtime="00:02:29.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="405" reactiontime="+84" swimtime="00:06:10.18" resultid="3094" heatid="8148" lane="6" entrytime="00:06:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.41" />
                    <SPLIT distance="100" swimtime="00:01:26.87" />
                    <SPLIT distance="150" swimtime="00:02:14.04" />
                    <SPLIT distance="200" swimtime="00:03:01.56" />
                    <SPLIT distance="250" swimtime="00:03:49.39" />
                    <SPLIT distance="300" swimtime="00:04:36.64" />
                    <SPLIT distance="350" swimtime="00:05:24.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="334" reactiontime="+70" swimtime="00:01:34.36" resultid="3095" heatid="8079" lane="9" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="434" reactiontime="+81" swimtime="00:02:48.77" resultid="3096" heatid="8090" lane="7" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.71" />
                    <SPLIT distance="100" swimtime="00:01:21.05" />
                    <SPLIT distance="150" swimtime="00:02:05.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-08-01" firstname="Małgorzata" gender="F" lastname="Polito" nation="POL" athleteid="3097">
              <RESULTS>
                <RESULT eventid="1120" points="514" reactiontime="+80" swimtime="00:11:55.76" resultid="3098" heatid="8136" lane="8" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.88" />
                    <SPLIT distance="100" swimtime="00:01:22.16" />
                    <SPLIT distance="150" swimtime="00:02:06.72" />
                    <SPLIT distance="200" swimtime="00:02:51.79" />
                    <SPLIT distance="250" swimtime="00:03:37.02" />
                    <SPLIT distance="300" swimtime="00:04:22.49" />
                    <SPLIT distance="350" swimtime="00:05:08.02" />
                    <SPLIT distance="400" swimtime="00:05:53.50" />
                    <SPLIT distance="450" swimtime="00:06:39.21" />
                    <SPLIT distance="500" swimtime="00:07:25.02" />
                    <SPLIT distance="550" swimtime="00:08:10.87" />
                    <SPLIT distance="600" swimtime="00:08:56.51" />
                    <SPLIT distance="650" swimtime="00:09:42.16" />
                    <SPLIT distance="700" swimtime="00:10:27.85" />
                    <SPLIT distance="750" swimtime="00:11:13.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="492" reactiontime="+72" swimtime="00:05:46.92" resultid="3099" heatid="8148" lane="4" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.65" />
                    <SPLIT distance="100" swimtime="00:01:23.01" />
                    <SPLIT distance="150" swimtime="00:02:07.25" />
                    <SPLIT distance="200" swimtime="00:02:51.69" />
                    <SPLIT distance="250" swimtime="00:03:35.34" />
                    <SPLIT distance="300" swimtime="00:04:19.93" />
                    <SPLIT distance="350" swimtime="00:05:04.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="475" swimtime="00:02:43.82" resultid="3100" heatid="8091" lane="9" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.76" />
                    <SPLIT distance="100" swimtime="00:01:19.32" />
                    <SPLIT distance="150" swimtime="00:02:01.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-09-29" firstname="Jakub" gender="M" lastname="Stępień" nation="POL" athleteid="3147">
              <RESULTS>
                <RESULT eventid="1105" points="356" reactiontime="+82" swimtime="00:00:35.28" resultid="3148" heatid="7965" lane="8" entrytime="00:00:35.20" />
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="3149" heatid="7987" lane="5" entrytime="00:01:05.80" />
                <RESULT eventid="1372" points="464" reactiontime="+80" swimtime="00:00:30.03" resultid="3150" heatid="8058" lane="5" entrytime="00:00:29.10" />
                <RESULT eventid="1509" points="442" reactiontime="+84" swimtime="00:02:31.85" resultid="3151" heatid="8099" lane="1" entrytime="00:02:30.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                    <SPLIT distance="100" swimtime="00:01:10.20" />
                    <SPLIT distance="150" swimtime="00:01:50.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-30" firstname="Paweł" gender="M" lastname="Gregorowicz" nation="POL" athleteid="3134">
              <RESULTS>
                <RESULT eventid="1075" points="675" reactiontime="+80" swimtime="00:02:30.93" resultid="3135" heatid="7948" lane="1" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.05" />
                    <SPLIT distance="100" swimtime="00:01:12.10" />
                    <SPLIT distance="150" swimtime="00:01:55.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="716" reactiontime="+76" swimtime="00:00:28.94" resultid="3136" heatid="7970" lane="7" entrytime="00:00:29.10" />
                <RESULT eventid="1198" points="799" reactiontime="+76" swimtime="00:00:58.53" resultid="3137" heatid="7992" lane="1" entrytime="00:00:58.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="768" reactiontime="+71" swimtime="00:00:26.84" resultid="3138" heatid="8058" lane="4" entrytime="00:00:29.10" />
                <RESULT eventid="1432" points="700" reactiontime="+81" swimtime="00:04:46.44" resultid="3139" heatid="8151" lane="0" entrytime="00:04:59.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                    <SPLIT distance="100" swimtime="00:01:07.58" />
                    <SPLIT distance="150" swimtime="00:01:43.56" />
                    <SPLIT distance="200" swimtime="00:02:20.47" />
                    <SPLIT distance="250" swimtime="00:02:56.81" />
                    <SPLIT distance="300" swimtime="00:03:33.63" />
                    <SPLIT distance="350" swimtime="00:04:10.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="759" reactiontime="+76" swimtime="00:02:09.89" resultid="3140" heatid="8101" lane="4" entrytime="00:02:12.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.95" />
                    <SPLIT distance="100" swimtime="00:01:02.71" />
                    <SPLIT distance="150" swimtime="00:01:35.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="620" reactiontime="+80" swimtime="00:05:31.75" resultid="3141" heatid="8163" lane="5" entrytime="00:05:50.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                    <SPLIT distance="100" swimtime="00:01:11.96" />
                    <SPLIT distance="150" swimtime="00:01:58.33" />
                    <SPLIT distance="200" swimtime="00:02:42.76" />
                    <SPLIT distance="250" swimtime="00:03:30.58" />
                    <SPLIT distance="300" swimtime="00:04:18.30" />
                    <SPLIT distance="350" swimtime="00:04:56.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-09-01" firstname="Marek" gender="M" lastname="Koźlikowski" nation="POL" athleteid="3152">
              <RESULTS>
                <RESULT eventid="1075" points="468" reactiontime="+94" swimtime="00:03:05.74" resultid="3153" heatid="7948" lane="2" entrytime="00:03:17.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                    <SPLIT distance="100" swimtime="00:01:35.38" />
                    <SPLIT distance="150" swimtime="00:02:26.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="493" reactiontime="+95" swimtime="00:03:22.53" resultid="3154" heatid="8073" lane="1" entrytime="00:03:35.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.41" />
                    <SPLIT distance="100" swimtime="00:01:38.29" />
                    <SPLIT distance="150" swimtime="00:02:31.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="429" reactiontime="+95" swimtime="00:06:01.35" resultid="3155" heatid="8154" lane="2" entrytime="00:06:10.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.77" />
                    <SPLIT distance="100" swimtime="00:01:25.79" />
                    <SPLIT distance="150" swimtime="00:02:12.99" />
                    <SPLIT distance="200" swimtime="00:03:00.97" />
                    <SPLIT distance="250" swimtime="00:03:48.50" />
                    <SPLIT distance="300" swimtime="00:04:35.62" />
                    <SPLIT distance="350" swimtime="00:05:19.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" status="DNS" swimtime="00:00:00.00" resultid="3156" heatid="8097" lane="1" entrytime="00:02:47.24" />
                <RESULT eventid="1599" points="468" reactiontime="+77" swimtime="00:06:50.38" resultid="3157" heatid="8165" lane="8" entrytime="00:07:05.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.52" />
                    <SPLIT distance="100" swimtime="00:01:44.87" />
                    <SPLIT distance="150" swimtime="00:02:41.80" />
                    <SPLIT distance="200" swimtime="00:03:36.96" />
                    <SPLIT distance="250" swimtime="00:04:30.60" />
                    <SPLIT distance="300" swimtime="00:05:24.65" />
                    <SPLIT distance="350" swimtime="00:06:08.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1318" reactiontime="+77" swimtime="00:04:16.26" resultid="3159" heatid="8031" lane="8" entrytime="00:04:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                    <SPLIT distance="100" swimtime="00:01:07.88" />
                    <SPLIT distance="150" swimtime="00:01:39.50" />
                    <SPLIT distance="200" swimtime="00:02:15.37" />
                    <SPLIT distance="250" swimtime="00:02:43.65" />
                    <SPLIT distance="300" swimtime="00:03:16.28" />
                    <SPLIT distance="350" swimtime="00:03:45.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3083" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="3128" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="3122" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="3134" number="4" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1303" reactiontime="+81" swimtime="00:04:55.44" resultid="3158" heatid="8029" lane="7" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.35" />
                    <SPLIT distance="100" swimtime="00:01:11.24" />
                    <SPLIT distance="150" swimtime="00:01:45.50" />
                    <SPLIT distance="200" swimtime="00:02:24.54" />
                    <SPLIT distance="250" swimtime="00:03:00.73" />
                    <SPLIT distance="300" swimtime="00:03:39.44" />
                    <SPLIT distance="350" swimtime="00:04:15.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3115" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="3101" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="3097" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="3108" number="4" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1614" reactiontime="+79" swimtime="00:02:15.79" resultid="3160" heatid="8135" lane="0" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.46" />
                    <SPLIT distance="100" swimtime="00:01:14.17" />
                    <SPLIT distance="150" swimtime="00:01:48.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3115" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="3122" number="2" />
                    <RELAYPOSITION athleteid="3101" number="3" reactiontime="+13" />
                    <RELAYPOSITION athleteid="3134" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1614" reactiontime="+93" swimtime="00:02:31.38" resultid="3161" heatid="8134" lane="9" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.73" />
                    <SPLIT distance="100" swimtime="00:01:18.92" />
                    <SPLIT distance="150" swimtime="00:01:59.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3083" number="1" reactiontime="+93" />
                    <RELAYPOSITION athleteid="3097" number="2" />
                    <RELAYPOSITION athleteid="3090" number="3" reactiontime="+10" />
                    <RELAYPOSITION athleteid="3152" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3162" name="AquaStars Gdynia">
          <CONTACT name="GOLON MARIUSZ" />
          <ATHLETES>
            <ATHLETE birthdate="1978-01-01" firstname="Mariusz" gender="M" lastname="Golon" nation="POL" athleteid="3168">
              <RESULTS>
                <RESULT eventid="1105" points="685" reactiontime="+84" swimtime="00:00:28.95" resultid="3169" heatid="7965" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1228" points="588" reactiontime="+81" swimtime="00:00:34.86" resultid="3170" heatid="8003" lane="5" entrytime="00:00:42.00" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="3171" heatid="8025" lane="0" entrytime="00:03:05.00" />
                <RESULT eventid="1342" points="601" reactiontime="+79" swimtime="00:01:13.50" resultid="3172" heatid="8039" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" status="DNS" swimtime="00:00:00.00" resultid="3173" heatid="8084" lane="9" entrytime="00:01:25.00" />
                <RESULT eventid="1539" points="368" reactiontime="+80" swimtime="00:00:39.33" resultid="3174" heatid="8112" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1569" points="536" reactiontime="+91" swimtime="00:01:21.79" resultid="3175" heatid="8128" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AWBIA" nation="POL" region="LBL" clubid="5329" name="AZS AWF Biała Podlaska">
          <CONTACT email="zielakko@gmail.com" name="Zieliński Kamil" phone="781529483" />
          <ATHLETES>
            <ATHLETE birthdate="1989-04-27" firstname="Kamil" gender="M" lastname="Zieliński" nation="POL" license="S02203200002" athleteid="5337">
              <RESULTS>
                <RESULT eventid="1228" points="757" reactiontime="+65" swimtime="00:00:32.14" resultid="5340" heatid="8010" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1372" points="624" reactiontime="+66" swimtime="00:00:27.08" resultid="5341" heatid="8052" lane="2" entrytime="00:00:48.00" />
                <RESULT eventid="1402" points="773" reactiontime="+71" swimtime="00:02:39.42" resultid="5342" heatid="8077" lane="4" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                    <SPLIT distance="100" swimtime="00:01:17.64" />
                    <SPLIT distance="150" swimtime="00:01:58.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="721" reactiontime="+66" swimtime="00:01:12.11" resultid="5343" heatid="8132" lane="3" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="565" reactiontime="+72" swimtime="00:05:45.07" resultid="5344" heatid="8164" lane="7" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                    <SPLIT distance="100" swimtime="00:01:16.99" />
                    <SPLIT distance="150" swimtime="00:02:05.48" />
                    <SPLIT distance="200" swimtime="00:02:53.49" />
                    <SPLIT distance="250" swimtime="00:03:36.66" />
                    <SPLIT distance="300" swimtime="00:04:20.69" />
                    <SPLIT distance="350" swimtime="00:05:03.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00611" nation="POL" region="SLA" clubid="3176" name="AZS AWF Katowice">
          <CONTACT city="Katowice" email="m.skora@awf.katowice.pl" name="Michał Skóra" phone="501 370 222" state="ŚLĄSK" street="Mikołowska 72a" zip="40-065" />
          <ATHLETES>
            <ATHLETE birthdate="1931-04-27" firstname="Jan" gender="M" lastname="Ślężyński" nation="POL" athleteid="3177">
              <RESULTS>
                <RESULT eventid="1165" points="186" reactiontime="+104" swimtime="00:47:39.65" resultid="3178" heatid="8146" lane="3" entrytime="00:44:50.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.06" />
                    <SPLIT distance="100" swimtime="00:02:42.82" />
                    <SPLIT distance="150" swimtime="00:04:21.97" />
                    <SPLIT distance="200" swimtime="00:05:59.34" />
                    <SPLIT distance="250" swimtime="00:07:28.45" />
                    <SPLIT distance="300" swimtime="00:09:00.26" />
                    <SPLIT distance="350" swimtime="00:10:40.38" />
                    <SPLIT distance="400" swimtime="00:12:21.65" />
                    <SPLIT distance="450" swimtime="00:13:52.72" />
                    <SPLIT distance="500" swimtime="00:15:24.73" />
                    <SPLIT distance="550" swimtime="00:17:07.36" />
                    <SPLIT distance="600" swimtime="00:18:48.80" />
                    <SPLIT distance="650" swimtime="00:20:20.38" />
                    <SPLIT distance="700" swimtime="00:21:54.75" />
                    <SPLIT distance="750" swimtime="00:23:36.87" />
                    <SPLIT distance="800" swimtime="00:25:17.08" />
                    <SPLIT distance="850" swimtime="00:26:47.85" />
                    <SPLIT distance="900" swimtime="00:28:21.18" />
                    <SPLIT distance="950" swimtime="00:30:03.49" />
                    <SPLIT distance="1000" swimtime="00:31:44.37" />
                    <SPLIT distance="1050" swimtime="00:33:16.81" />
                    <SPLIT distance="1100" swimtime="00:34:51.90" />
                    <SPLIT distance="1150" swimtime="00:36:33.53" />
                    <SPLIT distance="1200" swimtime="00:38:13.31" />
                    <SPLIT distance="1250" swimtime="00:39:45.58" />
                    <SPLIT distance="1300" swimtime="00:41:21.57" />
                    <SPLIT distance="1350" swimtime="00:43:02.20" />
                    <SPLIT distance="1400" swimtime="00:44:44.72" />
                    <SPLIT distance="1450" swimtime="00:46:12.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="131" swimtime="00:02:47.13" resultid="3179" heatid="7981" lane="8" entrytime="00:02:21.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="283" reactiontime="+95" swimtime="00:01:08.08" resultid="3180" heatid="8000" lane="8" />
                <RESULT eventid="1402" points="262" reactiontime="+90" swimtime="00:05:56.24" resultid="3181" heatid="8071" lane="2" entrytime="00:05:32.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.20" />
                    <SPLIT distance="100" swimtime="00:02:54.14" />
                    <SPLIT distance="150" swimtime="00:04:28.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="159" reactiontime="+104" swimtime="00:05:46.06" resultid="3183" heatid="8093" lane="5" entrytime="00:05:03.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.43" />
                    <SPLIT distance="100" swimtime="00:02:44.61" />
                    <SPLIT distance="150" swimtime="00:04:22.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="261" reactiontime="+106" swimtime="00:02:42.45" resultid="3184" heatid="8125" lane="9" entrytime="00:02:38.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="189" swimtime="00:11:49.51" resultid="8336" heatid="8325" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.55" />
                    <SPLIT distance="100" swimtime="00:02:46.33" />
                    <SPLIT distance="150" swimtime="00:04:19.19" />
                    <SPLIT distance="200" swimtime="00:05:50.90" />
                    <SPLIT distance="250" swimtime="00:07:22.76" />
                    <SPLIT distance="300" swimtime="00:08:54.66" />
                    <SPLIT distance="350" swimtime="00:10:25.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3185" name="AZS WSB Dąbrowa Górnicza">
          <CONTACT name="Kaproń Kacper" />
          <ATHLETES>
            <ATHLETE birthdate="1993-02-05" firstname="Kacper" gender="M" lastname="Kaproń" nation="POL" athleteid="3193">
              <RESULTS>
                <RESULT eventid="1228" status="DNS" swimtime="00:00:00.00" resultid="3194" heatid="8009" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="1288" points="370" reactiontime="+80" swimtime="00:02:56.96" resultid="3195" heatid="8026" lane="1" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.20" />
                    <SPLIT distance="100" swimtime="00:01:22.29" />
                    <SPLIT distance="150" swimtime="00:02:08.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="436" reactiontime="+67" swimtime="00:01:16.93" resultid="3196" heatid="8040" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="418" reactiontime="+79" swimtime="00:03:12.82" resultid="3197" heatid="8076" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.33" />
                    <SPLIT distance="100" swimtime="00:01:34.32" />
                    <SPLIT distance="150" swimtime="00:02:25.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" status="DNS" swimtime="00:00:00.00" resultid="3198" heatid="8100" lane="3" entrytime="00:02:22.00" />
                <RESULT eventid="1539" status="DNS" swimtime="00:00:00.00" resultid="3199" heatid="8115" lane="2" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="BASTA" nation="POL" region="ZAC" clubid="3200" name="BARAKUDA Stargard">
          <CONTACT city="Stargard Szczec." email="jerzychelstowski@gmail.com" name="Chełstowski" phone="601914514" street="Pl.Majdanek 11" zip="73-110" />
          <ATHLETES>
            <ATHLETE birthdate="1956-10-16" firstname="Jerzy" gender="M" lastname="Chełstowski" nation="POL" athleteid="3201">
              <RESULTS>
                <RESULT eventid="1105" points="298" reactiontime="+86" swimtime="00:00:42.69" resultid="3202" heatid="7963" lane="7" entrytime="00:00:44.50" />
                <RESULT eventid="1165" points="362" reactiontime="+66" swimtime="00:27:39.71" resultid="3203" heatid="8145" lane="8" entrytime="00:29:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.25" />
                    <SPLIT distance="100" swimtime="00:01:41.63" />
                    <SPLIT distance="150" swimtime="00:02:38.33" />
                    <SPLIT distance="200" swimtime="00:03:34.87" />
                    <SPLIT distance="250" swimtime="00:04:31.16" />
                    <SPLIT distance="300" swimtime="00:05:27.47" />
                    <SPLIT distance="350" swimtime="00:06:23.55" />
                    <SPLIT distance="400" swimtime="00:07:19.90" />
                    <SPLIT distance="450" swimtime="00:08:16.94" />
                    <SPLIT distance="500" swimtime="00:09:11.87" />
                    <SPLIT distance="550" swimtime="00:10:08.35" />
                    <SPLIT distance="600" swimtime="00:11:03.90" />
                    <SPLIT distance="650" swimtime="00:12:00.66" />
                    <SPLIT distance="700" swimtime="00:12:57.02" />
                    <SPLIT distance="750" swimtime="00:13:52.00" />
                    <SPLIT distance="800" swimtime="00:14:47.88" />
                    <SPLIT distance="850" swimtime="00:15:44.26" />
                    <SPLIT distance="900" swimtime="00:16:40.28" />
                    <SPLIT distance="950" swimtime="00:17:35.80" />
                    <SPLIT distance="1000" swimtime="00:18:32.06" />
                    <SPLIT distance="1050" swimtime="00:19:28.25" />
                    <SPLIT distance="1100" swimtime="00:20:25.19" />
                    <SPLIT distance="1150" swimtime="00:23:14.18" />
                    <SPLIT distance="1200" swimtime="00:22:18.30" />
                    <SPLIT distance="1250" swimtime="00:25:03.99" />
                    <SPLIT distance="1300" swimtime="00:24:09.72" />
                    <SPLIT distance="1400" swimtime="00:25:59.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="386" reactiontime="+73" swimtime="00:01:23.44" resultid="3204" heatid="7983" lane="0" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="256" reactiontime="+71" swimtime="00:00:48.89" resultid="3205" heatid="8001" lane="4" entrytime="00:00:48.00" />
                <RESULT eventid="1372" points="450" reactiontime="+70" swimtime="00:00:34.70" resultid="3206" heatid="8053" lane="6" entrytime="00:00:38.00" />
                <RESULT eventid="1432" points="332" reactiontime="+77" swimtime="00:07:05.95" resultid="3207" heatid="8155" lane="2" entrytime="00:06:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.74" />
                    <SPLIT distance="100" swimtime="00:01:39.41" />
                    <SPLIT distance="150" swimtime="00:02:35.13" />
                    <SPLIT distance="200" swimtime="00:03:30.32" />
                    <SPLIT distance="250" swimtime="00:04:26.36" />
                    <SPLIT distance="300" swimtime="00:05:22.15" />
                    <SPLIT distance="350" swimtime="00:06:16.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="356" reactiontime="+68" swimtime="00:03:11.91" resultid="3208" heatid="8095" lane="2" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.03" />
                    <SPLIT distance="100" swimtime="00:01:34.75" />
                    <SPLIT distance="150" swimtime="00:02:26.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="266" reactiontime="+125" swimtime="00:00:50.46" resultid="3209" heatid="8111" lane="0" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-02" firstname="Jerzy" gender="M" lastname="Grzesiak" nation="POL" athleteid="3210">
              <RESULTS>
                <RESULT eventid="1165" points="226" reactiontime="+123" swimtime="00:33:36.27" resultid="3211" heatid="8145" lane="9" entrytime="00:34:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.55" />
                    <SPLIT distance="100" swimtime="00:01:59.60" />
                    <SPLIT distance="150" swimtime="00:03:06.39" />
                    <SPLIT distance="200" swimtime="00:04:12.57" />
                    <SPLIT distance="250" swimtime="00:05:19.24" />
                    <SPLIT distance="300" swimtime="00:06:26.11" />
                    <SPLIT distance="350" swimtime="00:07:33.11" />
                    <SPLIT distance="400" swimtime="00:08:40.38" />
                    <SPLIT distance="450" swimtime="00:09:47.47" />
                    <SPLIT distance="500" swimtime="00:10:54.18" />
                    <SPLIT distance="550" swimtime="00:12:01.28" />
                    <SPLIT distance="600" swimtime="00:13:08.70" />
                    <SPLIT distance="650" swimtime="00:14:17.69" />
                    <SPLIT distance="700" swimtime="00:15:25.26" />
                    <SPLIT distance="750" swimtime="00:16:33.10" />
                    <SPLIT distance="800" swimtime="00:17:39.08" />
                    <SPLIT distance="850" swimtime="00:18:46.84" />
                    <SPLIT distance="900" swimtime="00:19:53.33" />
                    <SPLIT distance="950" swimtime="00:21:01.39" />
                    <SPLIT distance="1000" swimtime="00:22:09.90" />
                    <SPLIT distance="1050" swimtime="00:23:20.31" />
                    <SPLIT distance="1100" swimtime="00:24:30.02" />
                    <SPLIT distance="1150" swimtime="00:25:40.58" />
                    <SPLIT distance="1200" swimtime="00:26:50.67" />
                    <SPLIT distance="1250" swimtime="00:28:00.78" />
                    <SPLIT distance="1300" swimtime="00:29:10.49" />
                    <SPLIT distance="1350" swimtime="00:30:19.12" />
                    <SPLIT distance="1400" swimtime="00:31:27.79" />
                    <SPLIT distance="1450" swimtime="00:32:36.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="206" reactiontime="+120" swimtime="00:01:43.19" resultid="3212" heatid="7982" lane="9" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="325" reactiontime="+117" swimtime="00:00:39.74" resultid="3213" heatid="8052" lane="4" entrytime="00:00:44.90" />
                <RESULT eventid="1432" points="199" reactiontime="+111" swimtime="00:08:49.97" resultid="3214" heatid="8156" lane="4" entrytime="00:07:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.33" />
                    <SPLIT distance="100" swimtime="00:02:05.78" />
                    <SPLIT distance="150" swimtime="00:03:14.80" />
                    <SPLIT distance="200" swimtime="00:04:24.52" />
                    <SPLIT distance="250" swimtime="00:05:33.88" />
                    <SPLIT distance="300" swimtime="00:06:43.57" />
                    <SPLIT distance="350" swimtime="00:07:50.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="228" reactiontime="+102" swimtime="00:03:51.83" resultid="3215" heatid="8094" lane="7" entrytime="00:03:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.96" />
                    <SPLIT distance="100" swimtime="00:01:53.13" />
                    <SPLIT distance="150" swimtime="00:02:55.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="108" reactiontime="+159" swimtime="00:01:10.42" resultid="3216" heatid="8109" lane="0" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="8168" name="Biegacze Szczecin">
          <ATHLETES>
            <ATHLETE birthdate="1978-05-31" firstname="Magdalena" gender="F" lastname="Miśkiewicz" nation="POL" athleteid="8170" />
            <ATHLETE birthdate="1959-07-15" firstname="Dariusz" gender="M" lastname="Kochanowicz" nation="POL" athleteid="3292">
              <RESULTS>
                <RESULT eventid="1372" points="536" reactiontime="+77" swimtime="00:00:32.74" resultid="3293" heatid="8055" lane="6" entrytime="00:00:32.70" />
                <RESULT eventid="1402" points="419" reactiontime="+83" swimtime="00:03:41.22" resultid="3294" heatid="8073" lane="6" entrytime="00:03:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.10" />
                    <SPLIT distance="100" swimtime="00:01:46.82" />
                    <SPLIT distance="150" swimtime="00:02:45.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-11-04" firstname="Kamil" gender="M" lastname="Zieliński" nation="POL" athleteid="8171" />
            <ATHLETE birthdate="1980-12-12" firstname="Dominika" gender="F" lastname="Zielińska" nation="POL" athleteid="2128">
              <RESULTS>
                <RESULT eventid="1058" points="498" reactiontime="+79" swimtime="00:03:08.19" resultid="2129" heatid="7942" lane="7" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.26" />
                    <SPLIT distance="100" swimtime="00:01:25.83" />
                    <SPLIT distance="150" swimtime="00:02:22.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="522" reactiontime="+78" swimtime="00:00:36.89" resultid="2130" heatid="7957" lane="9" entrytime="00:00:41.00" />
                <RESULT eventid="1273" points="555" reactiontime="+88" swimtime="00:03:01.20" resultid="2131" heatid="8019" lane="2" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.14" />
                    <SPLIT distance="100" swimtime="00:01:27.40" />
                    <SPLIT distance="150" swimtime="00:02:14.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="575" reactiontime="+77" swimtime="00:01:24.00" resultid="2132" heatid="8033" lane="3" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="535" reactiontime="+80" swimtime="00:00:33.81" resultid="2133" heatid="8047" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="1524" points="543" reactiontime="+79" swimtime="00:00:39.35" resultid="2134" heatid="8105" lane="3" entrytime="00:00:41.00" />
                <RESULT eventid="1493" points="471" reactiontime="+86" status="EXH" swimtime="00:02:50.16" resultid="8347" heatid="8087" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.16" />
                    <SPLIT distance="100" swimtime="00:01:19.53" />
                    <SPLIT distance="150" swimtime="00:02:05.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X">
              <RESULTS>
                <RESULT eventid="1614" reactiontime="+83" swimtime="00:03:05.89" resultid="8169" heatid="8133" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.69" />
                    <SPLIT distance="100" swimtime="00:01:54.33" />
                    <SPLIT distance="150" swimtime="00:02:31.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3292" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="8170" number="2" />
                    <RELAYPOSITION athleteid="2128" number="3" reactiontime="+64" />
                    <RELAYPOSITION athleteid="8171" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" clubid="6677" name="Bąbel Sport">
          <ATHLETES>
            <ATHLETE birthdate="1978-09-01" firstname="Andrzej" gender="M" lastname="Lemański" athleteid="3774">
              <RESULTS>
                <RESULT eventid="1075" points="547" reactiontime="+82" swimtime="00:02:45.14" resultid="3775" heatid="7951" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                    <SPLIT distance="100" swimtime="00:01:15.55" />
                    <SPLIT distance="150" swimtime="00:02:03.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="538" reactiontime="+79" swimtime="00:00:35.91" resultid="3776" heatid="8008" lane="0" entrytime="00:00:35.00" />
                <RESULT eventid="1599" points="546" reactiontime="+72" swimtime="00:05:57.09" resultid="3777" heatid="8163" lane="9" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                    <SPLIT distance="100" swimtime="00:01:17.73" />
                    <SPLIT distance="150" swimtime="00:02:06.18" />
                    <SPLIT distance="200" swimtime="00:02:53.52" />
                    <SPLIT distance="250" swimtime="00:03:42.63" />
                    <SPLIT distance="300" swimtime="00:04:32.97" />
                    <SPLIT distance="350" swimtime="00:05:15.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CKS SZCZEC" nation="POL" region="SZ" clubid="5262" name="CKS-SMS Szczecin">
          <CONTACT city="Szczecin" email="s.juszkiewicz@cks.szczecin.pl" internet="www.cks.szczecin.pl" name="Juszkiewicz" street="rydla 49" zip="70-783" />
          <ATHLETES>
            <ATHLETE birthdate="1995-05-16" firstname="Nikola" gender="F" lastname="Vacek" nation="POL" athleteid="5263">
              <RESULTS>
                <RESULT eventid="1090" points="721" reactiontime="+69" swimtime="00:00:31.09" resultid="5264" heatid="7960" lane="6" entrytime="00:00:31.68" />
                <RESULT eventid="1181" points="826" reactiontime="+69" swimtime="00:01:02.52" resultid="5265" heatid="7979" lane="2" entrytime="00:01:02.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="803" reactiontime="+70" swimtime="00:00:28.63" resultid="5266" heatid="8050" lane="2" entrytime="00:00:28.78" />
                <RESULT eventid="1493" points="718" reactiontime="+73" swimtime="00:02:23.11" resultid="5267" heatid="8091" lane="1" entrytime="00:02:40.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                    <SPLIT distance="100" swimtime="00:01:09.74" />
                    <SPLIT distance="150" swimtime="00:01:47.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="MAL" clubid="3279" name="Collegium Medicum UJ Masters Kraków" shortname="Collegium Medicum UJ Masters K">
          <CONTACT city="Kraków" email="MariuszBaranik@gmail.com" name="Mariusz Baranik" phone="698128222" street="Białoprądnicka 32c/3" zip="31-221" />
          <ATHLETES>
            <ATHLETE birthdate="1969-06-29" firstname="Mariusz" gender="M" lastname="Baranik" nation="POL" athleteid="3280">
              <RESULTS>
                <RESULT eventid="1105" points="801" reactiontime="+74" swimtime="00:00:29.32" resultid="3281" heatid="7970" lane="1" entrytime="00:00:29.20" />
                <RESULT eventid="1198" points="756" reactiontime="+75" swimtime="00:01:01.29" resultid="3282" heatid="7990" lane="5" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="796" reactiontime="+75" swimtime="00:00:27.14" resultid="3283" heatid="8062" lane="4" entrytime="00:00:27.00" />
                <RESULT eventid="1539" points="666" reactiontime="+72" swimtime="00:00:33.47" resultid="3284" heatid="8115" lane="3" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DELOD" nation="POL" region="LOD" clubid="3301" name="DELFIN MASTERS Łódź">
          <CONTACT city="Łódź" email="jblasiak@biol.uni.lodz.pl" name="Błasiak" phone="696033013" street="Podchorążych 35 m 20" zip="94-234" />
          <ATHLETES>
            <ATHLETE birthdate="1974-01-24" firstname="Piotr" gender="M" lastname="Gaede" nation="POL" athleteid="3307">
              <RESULTS>
                <RESULT eventid="1228" points="459" reactiontime="+81" swimtime="00:00:39.55" resultid="3308" heatid="8005" lane="6" entrytime="00:00:38.87" />
                <RESULT eventid="1569" points="483" reactiontime="+87" swimtime="00:01:27.55" resultid="3309" heatid="8130" lane="0" entrytime="00:01:22.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-04-11" firstname="Rafał" gender="M" lastname="Maciejewski" nation="POL" athleteid="3320">
              <RESULTS>
                <RESULT eventid="1198" points="372" reactiontime="+97" swimtime="00:01:15.49" resultid="3321" heatid="7984" lane="2" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="393" reactiontime="+96" swimtime="00:00:33.53" resultid="3322" heatid="8056" lane="9" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-05-26" firstname="Ewa" gender="F" lastname="Cieplucha" nation="POL" athleteid="3317">
              <RESULTS>
                <RESULT eventid="1326" points="698" reactiontime="+68" swimtime="00:01:17.97" resultid="3318" heatid="8034" lane="5" entrytime="00:01:20.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="701" reactiontime="+67" swimtime="00:00:35.92" resultid="3319" heatid="8106" lane="3" entrytime="00:00:36.31" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-06-03" firstname="Tomasz" gender="M" lastname="Wiaderny" nation="POL" athleteid="3327">
              <RESULTS>
                <RESULT eventid="1198" points="347" reactiontime="+91" swimtime="00:01:19.42" resultid="3328" heatid="7984" lane="6" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="391" reactiontime="+92" swimtime="00:00:34.38" resultid="3329" heatid="8056" lane="0" entrytime="00:00:32.00" />
                <RESULT eventid="1462" points="189" reactiontime="+110" swimtime="00:01:45.86" resultid="3330" heatid="8082" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="268" reactiontime="+98" swimtime="00:03:05.04" resultid="3331" heatid="8096" lane="7" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                    <SPLIT distance="100" swimtime="00:01:27.63" />
                    <SPLIT distance="150" swimtime="00:02:18.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-05-03" firstname="Adam" gender="M" lastname="Jerzykowski" nation="POL" athleteid="3302">
              <RESULTS>
                <RESULT eventid="1165" points="359" reactiontime="+117" swimtime="00:23:10.16" resultid="3303" heatid="8143" lane="1" entrytime="00:21:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.43" />
                    <SPLIT distance="100" swimtime="00:01:20.81" />
                    <SPLIT distance="150" swimtime="00:02:04.32" />
                    <SPLIT distance="200" swimtime="00:02:48.11" />
                    <SPLIT distance="250" swimtime="00:03:33.17" />
                    <SPLIT distance="300" swimtime="00:04:18.90" />
                    <SPLIT distance="350" swimtime="00:05:04.99" />
                    <SPLIT distance="400" swimtime="00:05:52.25" />
                    <SPLIT distance="450" swimtime="00:06:38.56" />
                    <SPLIT distance="500" swimtime="00:07:26.74" />
                    <SPLIT distance="550" swimtime="00:08:13.73" />
                    <SPLIT distance="600" swimtime="00:09:01.44" />
                    <SPLIT distance="650" swimtime="00:09:49.43" />
                    <SPLIT distance="700" swimtime="00:10:36.33" />
                    <SPLIT distance="750" swimtime="00:11:24.21" />
                    <SPLIT distance="800" swimtime="00:12:12.68" />
                    <SPLIT distance="850" swimtime="00:13:00.29" />
                    <SPLIT distance="900" swimtime="00:13:48.15" />
                    <SPLIT distance="950" swimtime="00:14:35.72" />
                    <SPLIT distance="1000" swimtime="00:15:24.52" />
                    <SPLIT distance="1050" swimtime="00:16:11.33" />
                    <SPLIT distance="1100" swimtime="00:16:59.14" />
                    <SPLIT distance="1150" swimtime="00:19:20.99" />
                    <SPLIT distance="1200" swimtime="00:18:33.85" />
                    <SPLIT distance="1250" swimtime="00:20:54.48" />
                    <SPLIT distance="1300" swimtime="00:20:07.33" />
                    <SPLIT distance="1400" swimtime="00:21:39.89" />
                    <SPLIT distance="1450" swimtime="00:22:27.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="3304" heatid="7985" lane="4" entrytime="00:01:10.00" />
                <RESULT eventid="1372" status="DNS" swimtime="00:00:00.00" resultid="3305" heatid="8059" lane="2" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-11" firstname="Arkadiusz" gender="M" lastname="Piecyk" nation="POL" athleteid="3323">
              <RESULTS>
                <RESULT eventid="1288" points="498" reactiontime="+89" swimtime="00:02:51.04" resultid="3324" heatid="8026" lane="3" entrytime="00:02:45.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                    <SPLIT distance="100" swimtime="00:01:15.43" />
                    <SPLIT distance="150" swimtime="00:02:00.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="627" reactiontime="+84" swimtime="00:01:13.53" resultid="3325" heatid="8040" lane="5" entrytime="00:01:18.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="610" reactiontime="+76" swimtime="00:00:33.59" resultid="3326" heatid="8112" lane="5" entrytime="00:00:37.45" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-03-16" firstname="Janusz" gender="M" lastname="Błasiak" nation="POL" athleteid="3310">
              <RESULTS>
                <RESULT eventid="1198" points="310" reactiontime="+77" swimtime="00:01:30.12" resultid="3311" heatid="7982" lane="4" entrytime="00:01:27.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="191" swimtime="00:04:54.46" resultid="3312" heatid="8014" lane="9" entrytime="00:05:04.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.37" />
                    <SPLIT distance="100" swimtime="00:02:21.94" />
                    <SPLIT distance="150" swimtime="00:03:40.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="356" reactiontime="+80" swimtime="00:00:38.56" resultid="3313" heatid="8053" lane="4" entrytime="00:00:37.43" />
                <RESULT eventid="1432" points="291" reactiontime="+91" swimtime="00:07:46.91" resultid="3314" heatid="8156" lane="5" entrytime="00:08:03.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.25" />
                    <SPLIT distance="100" swimtime="00:01:47.67" />
                    <SPLIT distance="150" swimtime="00:02:51.02" />
                    <SPLIT distance="200" swimtime="00:03:52.12" />
                    <SPLIT distance="250" swimtime="00:04:52.70" />
                    <SPLIT distance="300" swimtime="00:05:54.46" />
                    <SPLIT distance="350" swimtime="00:06:54.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="290" swimtime="00:03:34.03" resultid="3315" heatid="8095" lane="9" entrytime="00:03:26.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.89" />
                    <SPLIT distance="100" swimtime="00:01:37.61" />
                    <SPLIT distance="150" swimtime="00:02:39.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="244" reactiontime="+102" swimtime="00:09:24.35" resultid="3316" heatid="8167" lane="7" entrytime="00:09:57.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.53" />
                    <SPLIT distance="100" swimtime="00:02:20.53" />
                    <SPLIT distance="150" swimtime="00:03:36.58" />
                    <SPLIT distance="200" swimtime="00:04:49.70" />
                    <SPLIT distance="250" swimtime="00:06:09.66" />
                    <SPLIT distance="300" swimtime="00:07:30.05" />
                    <SPLIT distance="350" swimtime="00:08:29.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1318" swimtime="00:05:22.98" resultid="6038" heatid="8030" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.11" />
                    <SPLIT distance="100" swimtime="00:01:33.63" />
                    <SPLIT distance="150" swimtime="00:02:10.03" />
                    <SPLIT distance="200" swimtime="00:02:52.58" />
                    <SPLIT distance="250" swimtime="00:03:29.29" />
                    <SPLIT distance="300" swimtime="00:04:09.38" />
                    <SPLIT distance="350" swimtime="00:04:44.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3310" number="1" />
                    <RELAYPOSITION athleteid="3320" number="2" reactiontime="+89" />
                    <RELAYPOSITION athleteid="3327" number="3" reactiontime="+94" />
                    <RELAYPOSITION athleteid="3302" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="CZE" clubid="3333" name="Dr. Regele Károly Szenior Úszóklub (Hungary)" shortname="Dr. Regele Károly Szenior Úszó">
          <CONTACT name="Bagdi Ferenc" />
          <ATHLETES>
            <ATHLETE birthdate="1989-05-02" firstname="Ferenc" gender="M" lastname="Bagdi" nation="HUN" athleteid="3337">
              <RESULTS>
                <RESULT eventid="1075" points="417" reactiontime="+87" swimtime="00:02:48.50" resultid="3338" heatid="7949" lane="6" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                    <SPLIT distance="100" swimtime="00:01:14.79" />
                    <SPLIT distance="150" swimtime="00:02:04.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="507" reactiontime="+94" swimtime="00:01:04.81" resultid="3339" heatid="7988" lane="1" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="482" reactiontime="+83" swimtime="00:00:37.35" resultid="3340" heatid="8006" lane="0" entrytime="00:00:38.00" />
                <RESULT eventid="1372" points="512" reactiontime="+80" swimtime="00:00:28.92" resultid="3341" heatid="8057" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1402" points="481" reactiontime="+82" swimtime="00:03:06.81" resultid="3342" heatid="8075" lane="5" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.57" />
                    <SPLIT distance="100" swimtime="00:01:26.99" />
                    <SPLIT distance="150" swimtime="00:02:16.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="434" reactiontime="+83" swimtime="00:01:25.37" resultid="3343" heatid="8129" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="UKR" clubid="2114" name="Dynamo">
          <CONTACT city="Kharkiv" email="swimmer2003@ukr.net" name="Vadym Kutsenko" phone="+38 057 7204282" street="16 Novgorodska" zip="61145" />
          <ATHLETES>
            <ATHLETE birthdate="1945-05-05" firstname="Vadym" gender="M" lastname="Kutsenko" nation="UKR" license="001" athleteid="2115">
              <RESULTS>
                <RESULT eventid="1075" points="758" reactiontime="+129" swimtime="00:03:18.96" resultid="2116" heatid="7949" lane="2" entrytime="00:03:04.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.45" />
                    <SPLIT distance="100" swimtime="00:01:40.52" />
                    <SPLIT distance="150" swimtime="00:02:38.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="893" reactiontime="+123" swimtime="00:22:40.09" resultid="2117" heatid="8144" lane="4" entrytime="00:21:56.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.56" />
                    <SPLIT distance="100" swimtime="00:01:24.92" />
                    <SPLIT distance="150" swimtime="00:02:10.16" />
                    <SPLIT distance="200" swimtime="00:02:55.24" />
                    <SPLIT distance="250" swimtime="00:03:40.43" />
                    <SPLIT distance="300" swimtime="00:04:25.23" />
                    <SPLIT distance="350" swimtime="00:05:10.29" />
                    <SPLIT distance="400" swimtime="00:05:55.43" />
                    <SPLIT distance="450" swimtime="00:06:40.95" />
                    <SPLIT distance="500" swimtime="00:07:26.20" />
                    <SPLIT distance="550" swimtime="00:08:11.55" />
                    <SPLIT distance="600" swimtime="00:08:56.63" />
                    <SPLIT distance="650" swimtime="00:09:42.64" />
                    <SPLIT distance="700" swimtime="00:10:28.87" />
                    <SPLIT distance="750" swimtime="00:11:15.02" />
                    <SPLIT distance="800" swimtime="00:12:00.60" />
                    <SPLIT distance="850" swimtime="00:12:46.33" />
                    <SPLIT distance="900" swimtime="00:13:31.97" />
                    <SPLIT distance="950" swimtime="00:14:18.11" />
                    <SPLIT distance="1000" swimtime="00:15:03.75" />
                    <SPLIT distance="1050" swimtime="00:15:49.71" />
                    <SPLIT distance="1100" swimtime="00:16:35.60" />
                    <SPLIT distance="1150" swimtime="00:17:21.58" />
                    <SPLIT distance="1200" swimtime="00:18:07.18" />
                    <SPLIT distance="1250" swimtime="00:18:53.39" />
                    <SPLIT distance="1300" swimtime="00:19:39.29" />
                    <SPLIT distance="1350" swimtime="00:20:25.12" />
                    <SPLIT distance="1400" swimtime="00:21:10.87" />
                    <SPLIT distance="1450" swimtime="00:21:56.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="612" reactiontime="+125" swimtime="00:01:17.49" resultid="2118" heatid="7984" lane="7" entrytime="00:01:16.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="562" swimtime="00:03:43.34" resultid="2119" heatid="8015" lane="6" entrytime="00:03:23.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.71" />
                    <SPLIT distance="100" swimtime="00:01:46.76" />
                    <SPLIT distance="150" swimtime="00:02:46.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="835" reactiontime="+121" swimtime="00:05:45.81" resultid="2120" heatid="8153" lane="5" entrytime="00:05:29.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.52" />
                    <SPLIT distance="100" swimtime="00:01:23.98" />
                    <SPLIT distance="150" swimtime="00:02:08.77" />
                    <SPLIT distance="200" swimtime="00:02:52.87" />
                    <SPLIT distance="250" swimtime="00:03:37.40" />
                    <SPLIT distance="300" swimtime="00:04:21.06" />
                    <SPLIT distance="350" swimtime="00:05:04.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="834" reactiontime="+120" swimtime="00:02:42.43" resultid="2121" heatid="8098" lane="3" entrytime="00:02:37.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                    <SPLIT distance="100" swimtime="00:01:19.51" />
                    <SPLIT distance="150" swimtime="00:02:02.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="1009" reactiontime="+104" swimtime="00:06:55.05" resultid="2122" heatid="8164" lane="1" entrytime="00:06:34.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.65" />
                    <SPLIT distance="100" swimtime="00:01:44.72" />
                    <SPLIT distance="150" swimtime="00:02:40.31" />
                    <SPLIT distance="200" swimtime="00:03:32.12" />
                    <SPLIT distance="250" swimtime="00:04:32.38" />
                    <SPLIT distance="300" swimtime="00:05:31.68" />
                    <SPLIT distance="350" swimtime="00:06:14.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3348" name="GB Sport Rzeszów">
          <CONTACT name="Bartek Czarnota" />
          <ATHLETES>
            <ATHLETE birthdate="1977-02-01" firstname="Mariusz" gender="M" lastname="Wójcicki" nation="POL" athleteid="3363">
              <RESULTS>
                <RESULT eventid="1105" points="472" reactiontime="+77" swimtime="00:00:32.76" resultid="3364" heatid="7968" lane="1" entrytime="00:00:31.80" />
                <RESULT eventid="1288" points="446" reactiontime="+65" swimtime="00:02:54.75" resultid="3365" heatid="8022" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.04" />
                    <SPLIT distance="100" swimtime="00:01:21.59" />
                    <SPLIT distance="150" swimtime="00:02:08.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="449" reactiontime="+61" swimtime="00:01:20.96" resultid="3366" heatid="8041" lane="7" entrytime="00:01:15.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="494" reactiontime="+84" swimtime="00:01:13.64" resultid="3367" heatid="8084" lane="4" entrytime="00:01:13.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="482" reactiontime="+61" swimtime="00:00:35.95" resultid="3368" heatid="8114" lane="3" entrytime="00:00:33.61" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-04-18" firstname="Sergiej" gender="M" lastname="Wojciechowski" nation="POL" athleteid="3354">
              <RESULTS>
                <RESULT eventid="1105" points="479" reactiontime="+82" swimtime="00:00:32.04" resultid="3355" heatid="7971" lane="1" entrytime="00:00:28.56" />
                <RESULT eventid="1135" points="359" reactiontime="+78" swimtime="00:12:13.01" resultid="3356" heatid="8139" lane="5" entrytime="00:10:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                    <SPLIT distance="100" swimtime="00:01:15.31" />
                    <SPLIT distance="150" swimtime="00:01:57.78" />
                    <SPLIT distance="200" swimtime="00:02:42.25" />
                    <SPLIT distance="250" swimtime="00:03:29.09" />
                    <SPLIT distance="300" swimtime="00:04:16.06" />
                    <SPLIT distance="350" swimtime="00:05:03.81" />
                    <SPLIT distance="400" swimtime="00:05:51.98" />
                    <SPLIT distance="450" swimtime="00:06:39.64" />
                    <SPLIT distance="500" swimtime="00:07:27.48" />
                    <SPLIT distance="550" swimtime="00:08:15.01" />
                    <SPLIT distance="600" swimtime="00:09:02.24" />
                    <SPLIT distance="650" swimtime="00:09:50.94" />
                    <SPLIT distance="700" swimtime="00:10:39.44" />
                    <SPLIT distance="750" swimtime="00:11:27.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="588" reactiontime="+74" swimtime="00:01:01.70" resultid="3357" heatid="7991" lane="4" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="566" reactiontime="+85" swimtime="00:00:35.41" resultid="3358" heatid="8008" lane="5" entrytime="00:00:34.00" />
                <RESULT eventid="1372" points="600" reactiontime="+86" swimtime="00:00:27.44" resultid="3359" heatid="8063" lane="1" entrytime="00:00:26.90" />
                <RESULT eventid="1402" points="507" reactiontime="+80" swimtime="00:03:03.49" resultid="3360" heatid="8077" lane="0" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.16" />
                    <SPLIT distance="100" swimtime="00:01:25.36" />
                    <SPLIT distance="150" swimtime="00:02:14.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="474" reactiontime="+82" swimtime="00:02:27.64" resultid="3361" heatid="8101" lane="1" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.12" />
                    <SPLIT distance="100" swimtime="00:01:05.24" />
                    <SPLIT distance="150" swimtime="00:01:44.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="530" reactiontime="+78" swimtime="00:01:19.90" resultid="3362" heatid="8131" lane="8" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-07-15" firstname="Grzegorz" gender="M" lastname="Wójcicki" nation="POL" athleteid="3369">
              <RESULTS>
                <RESULT eventid="1105" points="432" reactiontime="+72" swimtime="00:00:34.25" resultid="3370" heatid="7966" lane="2" entrytime="00:00:33.40" />
                <RESULT eventid="1198" points="455" reactiontime="+71" swimtime="00:01:10.59" resultid="3371" heatid="7987" lane="8" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="400" reactiontime="+80" swimtime="00:00:41.39" resultid="3372" heatid="8006" lane="1" entrytime="00:00:37.78" />
                <RESULT eventid="1372" points="542" reactiontime="+75" swimtime="00:00:30.13" resultid="3373" heatid="8058" lane="0" entrytime="00:00:29.78" />
                <RESULT eventid="1569" status="DNS" swimtime="00:00:00.00" resultid="3374" heatid="8130" lane="5" entrytime="00:01:19.54" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-17" firstname="Tomasz" gender="M" lastname="Pustelak" nation="POL" athleteid="3349">
              <RESULTS>
                <RESULT eventid="1105" points="371" reactiontime="+79" swimtime="00:00:34.86" resultid="3350" heatid="7967" lane="4" entrytime="00:00:32.30" />
                <RESULT eventid="1198" points="446" reactiontime="+79" swimtime="00:01:07.67" resultid="3351" heatid="7987" lane="4" entrytime="00:01:05.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="500" reactiontime="+82" swimtime="00:00:29.16" resultid="3352" heatid="8062" lane="7" entrytime="00:00:27.76" />
                <RESULT eventid="1539" status="DNS" swimtime="00:00:00.00" resultid="3353" heatid="8115" lane="1" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1318" reactiontime="+89" swimtime="00:04:28.22" resultid="3375" heatid="8030" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.00" />
                    <SPLIT distance="100" swimtime="00:01:07.14" />
                    <SPLIT distance="150" swimtime="00:01:36.14" />
                    <SPLIT distance="200" swimtime="00:02:11.53" />
                    <SPLIT distance="250" swimtime="00:02:43.20" />
                    <SPLIT distance="300" swimtime="00:03:21.61" />
                    <SPLIT distance="350" swimtime="00:03:52.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3349" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="3354" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="3369" number="3" reactiontime="+7" />
                    <RELAYPOSITION athleteid="3363" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="RUS" clubid="4697" name="GCOLIFK-masters">
          <CONTACT name="Tabakova" />
          <ATHLETES>
            <ATHLETE birthdate="1967-04-14" firstname="Elena" gender="F" lastname="Tabakova" nation="RUS" athleteid="4698">
              <RESULTS>
                <RESULT eventid="1150" points="575" reactiontime="+114" swimtime="00:24:46.36" resultid="4699" heatid="8142" lane="6" entrytime="00:26:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.45" />
                    <SPLIT distance="100" swimtime="00:01:27.66" />
                    <SPLIT distance="150" swimtime="00:02:15.93" />
                    <SPLIT distance="200" swimtime="00:03:05.67" />
                    <SPLIT distance="250" swimtime="00:03:54.81" />
                    <SPLIT distance="300" swimtime="00:04:45.08" />
                    <SPLIT distance="350" swimtime="00:05:34.84" />
                    <SPLIT distance="400" swimtime="00:06:24.82" />
                    <SPLIT distance="450" swimtime="00:07:14.86" />
                    <SPLIT distance="500" swimtime="00:08:05.06" />
                    <SPLIT distance="550" swimtime="00:08:54.70" />
                    <SPLIT distance="600" swimtime="00:09:44.32" />
                    <SPLIT distance="650" swimtime="00:10:34.08" />
                    <SPLIT distance="700" swimtime="00:11:23.95" />
                    <SPLIT distance="750" swimtime="00:12:13.78" />
                    <SPLIT distance="800" swimtime="00:13:03.63" />
                    <SPLIT distance="850" swimtime="00:13:53.30" />
                    <SPLIT distance="900" swimtime="00:14:43.63" />
                    <SPLIT distance="950" swimtime="00:15:33.76" />
                    <SPLIT distance="1000" swimtime="00:16:24.29" />
                    <SPLIT distance="1050" swimtime="00:17:14.36" />
                    <SPLIT distance="1100" swimtime="00:18:05.40" />
                    <SPLIT distance="1150" swimtime="00:18:55.36" />
                    <SPLIT distance="1200" swimtime="00:19:45.83" />
                    <SPLIT distance="1250" swimtime="00:20:36.00" />
                    <SPLIT distance="1300" swimtime="00:21:27.01" />
                    <SPLIT distance="1350" swimtime="00:22:16.83" />
                    <SPLIT distance="1400" swimtime="00:23:08.04" />
                    <SPLIT distance="1450" swimtime="00:23:58.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="454" reactiontime="+102" swimtime="00:00:47.59" resultid="4700" heatid="7996" lane="1" entrytime="00:00:48.00" />
                <RESULT eventid="1447" points="376" reactiontime="+107" swimtime="00:01:36.47" resultid="4701" heatid="8078" lane="3" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1584" points="444" reactiontime="+112" swimtime="00:07:15.99" resultid="4702" heatid="8160" lane="0" entrytime="00:07:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.01" />
                    <SPLIT distance="100" swimtime="00:01:41.03" />
                    <SPLIT distance="150" swimtime="00:02:35.86" />
                    <SPLIT distance="200" swimtime="00:03:31.42" />
                    <SPLIT distance="250" swimtime="00:04:31.56" />
                    <SPLIT distance="300" swimtime="00:05:34.53" />
                    <SPLIT distance="350" swimtime="00:06:25.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3376" name="Gdynia masters">
          <CONTACT email="k.mysiak@wpit.am.gdynia.pl" name="Mysiak" />
          <ATHLETES>
            <ATHLETE birthdate="1953-01-01" firstname="Andrzej" gender="M" lastname="Jacaszek" nation="POL" athleteid="3401">
              <RESULTS>
                <RESULT eventid="1228" points="565" reactiontime="+102" swimtime="00:00:41.53" resultid="3402" heatid="8003" lane="6" entrytime="00:00:42.00" />
                <RESULT eventid="1402" points="646" reactiontime="+84" swimtime="00:03:26.98" resultid="3403" heatid="8073" lane="8" entrytime="00:03:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.43" />
                    <SPLIT distance="100" swimtime="00:01:41.38" />
                    <SPLIT distance="150" swimtime="00:02:36.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="640" reactiontime="+98" swimtime="00:01:32.03" resultid="3404" heatid="8127" lane="6" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-01" firstname="Barbara" gender="F" lastname="Chomicka" nation="POL" athleteid="3413">
              <RESULTS>
                <RESULT eventid="1058" points="231" reactiontime="+104" swimtime="00:04:49.94" resultid="3414" heatid="7941" lane="5" entrytime="00:04:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.23" />
                    <SPLIT distance="100" swimtime="00:02:23.38" />
                    <SPLIT distance="150" swimtime="00:03:43.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="166" reactiontime="+99" swimtime="00:01:03.71" resultid="3415" heatid="7955" lane="8" entrytime="00:01:00.00" />
                <RESULT eventid="1243" points="278" reactiontime="+104" swimtime="00:05:09.53" resultid="3416" heatid="8011" lane="3" entrytime="00:05:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.18" />
                    <SPLIT distance="100" swimtime="00:02:30.96" />
                    <SPLIT distance="150" swimtime="00:03:51.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="285" reactiontime="+78" swimtime="00:04:49.54" resultid="3417" heatid="8018" lane="6" entrytime="00:04:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.72" />
                    <SPLIT distance="100" swimtime="00:02:26.19" />
                    <SPLIT distance="150" swimtime="00:03:40.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="261" reactiontime="+74" swimtime="00:02:09.40" resultid="3418" heatid="8032" lane="4" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="163" reactiontime="+106" swimtime="00:02:28.51" resultid="3419" heatid="8078" lane="0" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="353" reactiontime="+73" swimtime="00:00:56.81" resultid="3420" heatid="8104" lane="7" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-01-01" firstname="Andrzej" gender="M" lastname="Skwarło" nation="POL" athleteid="3421">
              <RESULTS>
                <RESULT eventid="1075" points="487" reactiontime="+105" swimtime="00:03:58.00" resultid="3422" heatid="7947" lane="9" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.52" />
                    <SPLIT distance="100" swimtime="00:01:59.27" />
                    <SPLIT distance="150" swimtime="00:03:03.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="502" reactiontime="+107" swimtime="00:00:46.20" resultid="3423" heatid="7963" lane="1" entrytime="00:00:45.50" />
                <RESULT eventid="1228" points="636" reactiontime="+104" swimtime="00:00:46.00" resultid="3424" heatid="8002" lane="1" entrytime="00:00:45.50" />
                <RESULT eventid="1288" points="391" reactiontime="+90" swimtime="00:04:24.74" resultid="3425" heatid="8023" lane="4" entrytime="00:04:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.95" />
                    <SPLIT distance="100" swimtime="00:02:07.02" />
                    <SPLIT distance="150" swimtime="00:03:19.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="434" reactiontime="+88" swimtime="00:01:58.02" resultid="3426" heatid="8037" lane="4" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="500" reactiontime="+112" swimtime="00:04:17.12" resultid="3427" heatid="8072" lane="7" entrytime="00:03:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.63" />
                    <SPLIT distance="100" swimtime="00:02:03.13" />
                    <SPLIT distance="150" swimtime="00:03:12.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="536" reactiontime="+87" swimtime="00:00:49.50" resultid="3428" heatid="8109" lane="3" entrytime="00:00:49.50" />
                <RESULT eventid="1569" points="597" reactiontime="+105" swimtime="00:01:46.75" resultid="3429" heatid="8126" lane="1" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Czesław" gender="M" lastname="Mikołajczyk" nation="POL" athleteid="3405">
              <RESULTS>
                <RESULT eventid="1075" points="382" reactiontime="+98" swimtime="00:03:48.11" resultid="3406" heatid="7947" lane="7" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.18" />
                    <SPLIT distance="100" swimtime="00:01:57.71" />
                    <SPLIT distance="150" swimtime="00:02:57.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="408" reactiontime="+100" swimtime="00:00:48.84" resultid="3407" heatid="8002" lane="0" entrytime="00:00:48.00" />
                <RESULT eventid="1258" points="296" reactiontime="+98" swimtime="00:04:23.99" resultid="3408" heatid="8015" lane="1" entrytime="00:04:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.77" />
                    <SPLIT distance="100" swimtime="00:02:04.97" />
                    <SPLIT distance="150" swimtime="00:03:13.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="530" swimtime="00:03:54.21" resultid="3409" heatid="8072" lane="3" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.97" />
                    <SPLIT distance="100" swimtime="00:01:55.13" />
                    <SPLIT distance="150" swimtime="00:02:54.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="193" reactiontime="+98" swimtime="00:02:06.37" resultid="3410" heatid="8082" lane="0" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="421" reactiontime="+94" swimtime="00:01:49.90" resultid="3411" heatid="8126" lane="7" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="479" reactiontime="+95" swimtime="00:08:02.05" resultid="3412" heatid="8166" lane="7" entrytime="00:08:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.61" />
                    <SPLIT distance="100" swimtime="00:02:07.00" />
                    <SPLIT distance="150" swimtime="00:03:11.82" />
                    <SPLIT distance="200" swimtime="00:04:12.36" />
                    <SPLIT distance="250" swimtime="00:05:14.28" />
                    <SPLIT distance="300" swimtime="00:06:15.59" />
                    <SPLIT distance="350" swimtime="00:07:10.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-01-01" firstname="Anna" gender="F" lastname="Walczak" nation="POL" athleteid="3439">
              <RESULTS>
                <RESULT eventid="1181" points="299" swimtime="00:01:52.08" resultid="3440" heatid="7974" lane="9" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="524" reactiontime="+69" swimtime="00:01:54.10" resultid="3441" heatid="8033" lane="0" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="318" reactiontime="+98" swimtime="00:00:49.16" resultid="3442" heatid="8045" lane="9" entrytime="00:00:48.00" />
                <RESULT eventid="1524" points="506" reactiontime="+55" swimtime="00:00:53.08" resultid="3443" heatid="8104" lane="5" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="Jerzy" gender="M" lastname="Pluskota" nation="POL" athleteid="3385">
              <RESULTS>
                <RESULT eventid="1105" points="309" reactiontime="+102" swimtime="00:00:45.12" resultid="3386" heatid="7962" lane="4" entrytime="00:00:50.00" />
                <RESULT eventid="1198" points="394" reactiontime="+93" swimtime="00:01:30.00" resultid="3387" heatid="7982" lane="6" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="560" reactiontime="+96" swimtime="00:00:34.92" resultid="3388" heatid="8054" lane="7" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-01-01" firstname="Katarzyna" gender="F" lastname="Mysiak" nation="POL" athleteid="3395">
              <RESULTS>
                <RESULT eventid="1120" points="343" reactiontime="+100" swimtime="00:14:42.94" resultid="3396" heatid="8137" lane="8" entrytime="00:15:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.52" />
                    <SPLIT distance="100" swimtime="00:01:39.51" />
                    <SPLIT distance="150" swimtime="00:02:35.01" />
                    <SPLIT distance="200" swimtime="00:03:30.27" />
                    <SPLIT distance="250" swimtime="00:04:27.01" />
                    <SPLIT distance="300" swimtime="00:05:23.50" />
                    <SPLIT distance="350" swimtime="00:06:20.41" />
                    <SPLIT distance="400" swimtime="00:07:17.34" />
                    <SPLIT distance="450" swimtime="00:08:14.00" />
                    <SPLIT distance="500" swimtime="00:09:11.35" />
                    <SPLIT distance="550" swimtime="00:10:07.51" />
                    <SPLIT distance="600" swimtime="00:11:04.97" />
                    <SPLIT distance="650" swimtime="00:12:01.42" />
                    <SPLIT distance="700" swimtime="00:12:58.15" />
                    <SPLIT distance="750" swimtime="00:13:52.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="415" reactiontime="+99" swimtime="00:03:43.81" resultid="3397" heatid="8019" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.68" />
                    <SPLIT distance="100" swimtime="00:01:47.95" />
                    <SPLIT distance="150" swimtime="00:02:47.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="316" reactiontime="+102" swimtime="00:07:07.33" resultid="3398" heatid="8149" lane="5" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.19" />
                    <SPLIT distance="100" swimtime="00:01:37.56" />
                    <SPLIT distance="150" swimtime="00:02:32.11" />
                    <SPLIT distance="200" swimtime="00:03:27.43" />
                    <SPLIT distance="250" swimtime="00:04:23.02" />
                    <SPLIT distance="300" swimtime="00:05:19.61" />
                    <SPLIT distance="350" swimtime="00:06:15.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="323" reactiontime="+102" swimtime="00:03:21.17" resultid="3399" heatid="8088" lane="3" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.96" />
                    <SPLIT distance="100" swimtime="00:01:36.10" />
                    <SPLIT distance="150" swimtime="00:02:29.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="374" reactiontime="+88" swimtime="00:00:47.67" resultid="3400" heatid="8105" lane="7" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1934-01-01" firstname="Bogdan" gender="M" lastname="Ciundziewicki" nation="POL" athleteid="3380">
              <RESULTS>
                <RESULT eventid="1228" points="685" reactiontime="+89" swimtime="00:00:50.72" resultid="3381" heatid="8001" lane="3" entrytime="00:00:48.76" />
                <RESULT comment="Rekord Polski Masters" eventid="1402" points="760" reactiontime="+96" swimtime="00:04:09.80" resultid="3382" heatid="8071" lane="4" entrytime="00:04:11.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.67" />
                    <SPLIT distance="100" swimtime="00:01:58.95" />
                    <SPLIT distance="150" swimtime="00:03:05.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="739" reactiontime="+109" swimtime="00:00:49.54" resultid="3383" heatid="8110" lane="0" entrytime="00:00:48.76" />
                <RESULT eventid="1569" points="753" reactiontime="+95" swimtime="00:01:54.11" resultid="3384" heatid="8126" lane="8" entrytime="00:01:48.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-01" firstname="Maciej" gender="M" lastname="Piwowarczyk" nation="POL" athleteid="3389">
              <RESULTS>
                <RESULT eventid="1228" points="454" reactiontime="+93" swimtime="00:00:39.69" resultid="3390" heatid="8005" lane="7" entrytime="00:00:39.00" />
                <RESULT eventid="1342" points="380" reactiontime="+75" swimtime="00:01:26.84" resultid="3391" heatid="8039" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" status="DNS" swimtime="00:00:00.00" resultid="3392" heatid="8074" lane="2" entrytime="00:03:22.00" />
                <RESULT eventid="1539" points="437" reactiontime="+71" swimtime="00:00:37.54" resultid="3393" heatid="8112" lane="2" entrytime="00:00:38.00" />
                <RESULT eventid="1569" status="DNS" swimtime="00:00:00.00" resultid="3394" heatid="8129" lane="8" entrytime="00:01:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-01" firstname="Danuta" gender="F" lastname="Radkowiak" nation="POL" athleteid="3444">
              <RESULTS>
                <RESULT eventid="1058" points="376" reactiontime="+100" swimtime="00:04:00.48" resultid="3445" heatid="7942" lane="0" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.06" />
                    <SPLIT distance="100" swimtime="00:02:03.34" />
                    <SPLIT distance="150" swimtime="00:03:05.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="350" reactiontime="+95" swimtime="00:00:49.12" resultid="3446" heatid="7956" lane="6" entrytime="00:00:45.00" />
                <RESULT eventid="1213" points="404" reactiontime="+101" swimtime="00:00:51.86" resultid="3447" heatid="7996" lane="0" entrytime="00:00:50.00" />
                <RESULT eventid="1243" points="379" reactiontime="+94" swimtime="00:04:28.57" resultid="3448" heatid="8012" lane="9" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.37" />
                    <SPLIT distance="100" swimtime="00:02:05.50" />
                    <SPLIT distance="150" swimtime="00:03:15.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1387" points="431" reactiontime="+100" swimtime="00:04:14.13" resultid="3449" heatid="8068" lane="0" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.83" />
                    <SPLIT distance="100" swimtime="00:02:04.02" />
                    <SPLIT distance="150" swimtime="00:03:09.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" status="DNS" swimtime="00:00:00.00" resultid="3450" heatid="8078" lane="2" entrytime="00:01:50.00" />
                <RESULT eventid="1554" status="DNS" swimtime="00:00:00.00" resultid="3451" heatid="8120" lane="8" entrytime="00:01:50.00" />
                <RESULT eventid="1584" points="365" reactiontime="+97" swimtime="00:08:43.86" resultid="3452" heatid="8161" lane="4" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.78" />
                    <SPLIT distance="100" swimtime="00:02:02.50" />
                    <SPLIT distance="150" swimtime="00:03:19.45" />
                    <SPLIT distance="200" swimtime="00:04:33.42" />
                    <SPLIT distance="250" swimtime="00:05:43.55" />
                    <SPLIT distance="300" swimtime="00:06:52.68" />
                    <SPLIT distance="350" swimtime="00:07:50.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-01-01" firstname="Hanka" gender="F" lastname="Kania" nation="POL" athleteid="3430">
              <RESULTS>
                <RESULT eventid="1058" points="472" reactiontime="+118" swimtime="00:03:48.63" resultid="3431" heatid="7942" lane="1" entrytime="00:03:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.04" />
                    <SPLIT distance="100" swimtime="00:01:54.64" />
                    <SPLIT distance="150" swimtime="00:02:57.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="322" reactiontime="+106" swimtime="00:00:51.12" resultid="3432" heatid="7955" lane="3" entrytime="00:00:51.00" />
                <RESULT eventid="1181" points="427" reactiontime="+106" swimtime="00:01:33.30" resultid="3433" heatid="7974" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="399" reactiontime="+107" swimtime="00:00:52.23" resultid="3434" heatid="7995" lane="5" entrytime="00:00:52.00" />
                <RESULT eventid="1357" points="463" reactiontime="+108" swimtime="00:00:40.76" resultid="3435" heatid="8045" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1387" points="526" reactiontime="+109" swimtime="00:04:02.76" resultid="3436" heatid="8067" lane="6" entrytime="00:04:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.92" />
                    <SPLIT distance="100" swimtime="00:01:57.51" />
                    <SPLIT distance="150" swimtime="00:03:00.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="483" reactiontime="+116" swimtime="00:03:22.60" resultid="3437" heatid="8088" lane="5" entrytime="00:03:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.62" />
                    <SPLIT distance="100" swimtime="00:01:36.36" />
                    <SPLIT distance="150" swimtime="00:02:31.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="520" reactiontime="+114" swimtime="00:01:51.73" resultid="3438" heatid="8119" lane="4" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="280" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="3456" heatid="8031" lane="4" entrytime="00:03:40.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3380" number="1" />
                    <RELAYPOSITION athleteid="3401" number="2" />
                    <RELAYPOSITION athleteid="3385" number="3" />
                    <RELAYPOSITION athleteid="3421" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1303" status="DNS" swimtime="00:00:00.00" resultid="3453" heatid="8029" lane="4" entrytime="00:03:40.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3430" number="1" />
                    <RELAYPOSITION athleteid="3395" number="2" />
                    <RELAYPOSITION athleteid="3439" number="3" />
                    <RELAYPOSITION athleteid="3444" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="280" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1614" status="DNS" swimtime="00:00:00.00" resultid="3454" heatid="8133" lane="1" entrytime="00:03:40.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3439" number="1" />
                    <RELAYPOSITION athleteid="3380" number="2" />
                    <RELAYPOSITION athleteid="3430" number="3" />
                    <RELAYPOSITION athleteid="3421" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1614" status="DNS" swimtime="00:00:00.00" resultid="3455" heatid="8133" lane="0">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3395" number="1" />
                    <RELAYPOSITION athleteid="3405" number="2" />
                    <RELAYPOSITION athleteid="3444" number="3" />
                    <RELAYPOSITION athleteid="3385" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3488" name="Hasacze Szczecin">
          <CONTACT city="Szczecin" email="martahanczewska@yahoo.pl" name="Hanczewska Marta" phone="664935249" />
          <ATHLETES>
            <ATHLETE birthdate="1984-10-05" firstname="Marta" gender="F" lastname="Hanczewska" nation="POL" athleteid="3489">
              <RESULTS>
                <RESULT eventid="1213" points="448" swimtime="00:00:42.66" resultid="3490" heatid="7998" lane="5" entrytime="00:00:40.59" />
                <RESULT eventid="1357" points="516" reactiontime="+87" swimtime="00:00:33.85" resultid="3491" heatid="8048" lane="9" entrytime="00:00:33.09" />
                <RESULT eventid="1387" points="401" reactiontime="+89" swimtime="00:03:37.42" resultid="3492" heatid="8069" lane="8" entrytime="00:03:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.03" />
                    <SPLIT distance="100" swimtime="00:01:40.59" />
                    <SPLIT distance="150" swimtime="00:02:39.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="421" swimtime="00:01:37.51" resultid="3493" heatid="8122" lane="9" entrytime="00:01:32.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="AUS" clubid="3494" name="Hobart Aquatic Masters SC">
          <CONTACT name="Slugocki" />
          <ATHLETES>
            <ATHLETE birthdate="1952-12-13" firstname="Maciej" gender="M" lastname="Slugocki" nation="AUS" athleteid="3495">
              <RESULTS>
                <RESULT eventid="1075" points="813" reactiontime="+103" swimtime="00:02:53.90" resultid="3496" heatid="7950" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.99" />
                    <SPLIT distance="100" swimtime="00:01:24.92" />
                    <SPLIT distance="150" swimtime="00:02:15.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="976" swimtime="00:20:39.30" resultid="3497" heatid="8146" lane="9" entrytime="00:21:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.34" />
                    <SPLIT distance="100" swimtime="00:01:18.95" />
                    <SPLIT distance="150" swimtime="00:01:59.93" />
                    <SPLIT distance="200" swimtime="00:02:41.19" />
                    <SPLIT distance="250" swimtime="00:03:22.77" />
                    <SPLIT distance="300" swimtime="00:04:04.51" />
                    <SPLIT distance="350" swimtime="00:04:46.50" />
                    <SPLIT distance="400" swimtime="00:05:28.03" />
                    <SPLIT distance="450" swimtime="00:06:09.60" />
                    <SPLIT distance="500" swimtime="00:06:51.41" />
                    <SPLIT distance="550" swimtime="00:07:33.29" />
                    <SPLIT distance="600" swimtime="00:08:14.96" />
                    <SPLIT distance="650" swimtime="00:08:56.57" />
                    <SPLIT distance="700" swimtime="00:09:38.63" />
                    <SPLIT distance="750" swimtime="00:10:20.68" />
                    <SPLIT distance="800" swimtime="00:11:02.28" />
                    <SPLIT distance="850" swimtime="00:11:43.95" />
                    <SPLIT distance="900" swimtime="00:12:25.40" />
                    <SPLIT distance="950" swimtime="00:13:06.96" />
                    <SPLIT distance="1000" swimtime="00:13:48.23" />
                    <SPLIT distance="1050" swimtime="00:14:29.85" />
                    <SPLIT distance="1100" swimtime="00:15:11.28" />
                    <SPLIT distance="1150" swimtime="00:15:52.02" />
                    <SPLIT distance="1200" swimtime="00:16:33.09" />
                    <SPLIT distance="1250" swimtime="00:17:14.47" />
                    <SPLIT distance="1300" swimtime="00:17:56.17" />
                    <SPLIT distance="1350" swimtime="00:18:38.06" />
                    <SPLIT distance="1400" swimtime="00:19:19.89" />
                    <SPLIT distance="1450" swimtime="00:20:00.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="683" reactiontime="+98" swimtime="00:01:09.30" resultid="3498" heatid="7986" lane="7" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1258" points="705" reactiontime="+103" swimtime="00:03:10.67" resultid="3499" heatid="8016" lane="1" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.65" />
                    <SPLIT distance="100" swimtime="00:01:31.61" />
                    <SPLIT distance="150" swimtime="00:02:21.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="891" reactiontime="+97" swimtime="00:05:21.78" resultid="3500" heatid="8152" lane="1" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                    <SPLIT distance="100" swimtime="00:01:19.29" />
                    <SPLIT distance="150" swimtime="00:02:00.11" />
                    <SPLIT distance="200" swimtime="00:02:41.04" />
                    <SPLIT distance="250" swimtime="00:03:21.99" />
                    <SPLIT distance="300" swimtime="00:04:03.19" />
                    <SPLIT distance="350" swimtime="00:04:43.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="647" reactiontime="+78" swimtime="00:01:22.74" resultid="3501" heatid="8084" lane="8" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="863" reactiontime="+90" swimtime="00:02:28.87" resultid="3502" heatid="8099" lane="6" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.52" />
                    <SPLIT distance="100" swimtime="00:01:13.27" />
                    <SPLIT distance="150" swimtime="00:01:51.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="815" reactiontime="+96" swimtime="00:06:17.52" resultid="3503" heatid="8164" lane="5" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.44" />
                    <SPLIT distance="100" swimtime="00:01:30.67" />
                    <SPLIT distance="150" swimtime="00:02:22.37" />
                    <SPLIT distance="200" swimtime="00:03:11.71" />
                    <SPLIT distance="250" swimtime="00:04:05.67" />
                    <SPLIT distance="300" swimtime="00:04:59.67" />
                    <SPLIT distance="350" swimtime="00:05:39.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZWAW" nation="POL" region="WA" clubid="3723" name="K.S. niezrzeszeni.pl">
          <CONTACT name="K.S. niezrzeszeni.pl" />
          <ATHLETES>
            <ATHLETE birthdate="1960-07-16" firstname="Matylda" gender="F" lastname="Wawer" nation="POL" athleteid="3743">
              <RESULTS>
                <RESULT eventid="1058" points="348" reactiontime="+82" swimtime="00:04:06.82" resultid="3744" heatid="7941" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.10" />
                    <SPLIT distance="100" swimtime="00:01:58.80" />
                    <SPLIT distance="150" swimtime="00:03:14.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="380" swimtime="00:00:47.80" resultid="3745" heatid="7956" lane="9" entrytime="00:00:47.00" />
                <RESULT eventid="1181" points="480" reactiontime="+89" swimtime="00:01:28.27" resultid="3746" heatid="7975" lane="0" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="561" reactiontime="+86" swimtime="00:00:37.43" resultid="3747" heatid="8046" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="1447" points="303" reactiontime="+96" swimtime="00:01:58.02" resultid="3748" heatid="8078" lane="1" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="444" reactiontime="+90" swimtime="00:03:25.51" resultid="3749" heatid="8088" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.23" />
                    <SPLIT distance="100" swimtime="00:01:35.99" />
                    <SPLIT distance="150" swimtime="00:02:31.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-08-26" firstname="Małgorzata" gender="F" lastname="Piechura" nation="POL" athleteid="3738">
              <RESULTS>
                <RESULT eventid="1058" points="234" swimtime="00:04:05.62" resultid="3739" heatid="7942" lane="9" entrytime="00:04:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.61" />
                    <SPLIT distance="100" swimtime="00:02:08.19" />
                    <SPLIT distance="150" swimtime="00:03:14.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="141" reactiontime="+111" swimtime="00:00:57.11" resultid="3740" heatid="7955" lane="1" entrytime="00:00:58.00" />
                <RESULT eventid="1417" points="233" reactiontime="+101" swimtime="00:07:39.49" resultid="3741" heatid="8149" lane="1" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.07" />
                    <SPLIT distance="100" swimtime="00:01:43.01" />
                    <SPLIT distance="150" swimtime="00:02:41.05" />
                    <SPLIT distance="200" swimtime="00:03:39.58" />
                    <SPLIT distance="250" swimtime="00:04:39.50" />
                    <SPLIT distance="300" swimtime="00:05:41.39" />
                    <SPLIT distance="350" swimtime="00:06:41.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="229" reactiontime="+110" swimtime="00:03:37.58" resultid="3742" heatid="8088" lane="6" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.07" />
                    <SPLIT distance="100" swimtime="00:01:40.60" />
                    <SPLIT distance="150" swimtime="00:02:38.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-14" firstname="Andrzej" gender="M" lastname="Miński" nation="POL" athleteid="3733">
              <RESULTS>
                <RESULT eventid="1165" points="393" reactiontime="+134" swimtime="00:26:55.34" resultid="3734" heatid="8145" lane="5" entrytime="00:26:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.05" />
                    <SPLIT distance="100" swimtime="00:01:40.72" />
                    <SPLIT distance="150" swimtime="00:02:33.98" />
                    <SPLIT distance="200" swimtime="00:03:28.32" />
                    <SPLIT distance="250" swimtime="00:04:22.64" />
                    <SPLIT distance="300" swimtime="00:05:17.55" />
                    <SPLIT distance="350" swimtime="00:06:11.15" />
                    <SPLIT distance="400" swimtime="00:07:06.12" />
                    <SPLIT distance="450" swimtime="00:08:00.49" />
                    <SPLIT distance="500" swimtime="00:08:55.46" />
                    <SPLIT distance="550" swimtime="00:09:49.98" />
                    <SPLIT distance="600" swimtime="00:10:44.23" />
                    <SPLIT distance="650" swimtime="00:11:38.41" />
                    <SPLIT distance="700" swimtime="00:12:32.82" />
                    <SPLIT distance="750" swimtime="00:13:25.88" />
                    <SPLIT distance="800" swimtime="00:14:18.79" />
                    <SPLIT distance="850" swimtime="00:15:13.02" />
                    <SPLIT distance="900" swimtime="00:16:07.68" />
                    <SPLIT distance="950" swimtime="00:17:01.21" />
                    <SPLIT distance="1000" swimtime="00:17:55.12" />
                    <SPLIT distance="1050" swimtime="00:18:50.49" />
                    <SPLIT distance="1100" swimtime="00:19:45.18" />
                    <SPLIT distance="1150" swimtime="00:20:39.32" />
                    <SPLIT distance="1200" swimtime="00:21:33.81" />
                    <SPLIT distance="1250" swimtime="00:22:28.27" />
                    <SPLIT distance="1300" swimtime="00:23:22.75" />
                    <SPLIT distance="1350" swimtime="00:24:17.36" />
                    <SPLIT distance="1400" swimtime="00:25:12.66" />
                    <SPLIT distance="1450" swimtime="00:26:05.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="355" swimtime="00:06:56.34" resultid="3735" heatid="8154" lane="9" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.40" />
                    <SPLIT distance="100" swimtime="00:01:36.53" />
                    <SPLIT distance="150" swimtime="00:02:30.56" />
                    <SPLIT distance="200" swimtime="00:03:25.03" />
                    <SPLIT distance="250" swimtime="00:04:19.43" />
                    <SPLIT distance="300" swimtime="00:05:14.61" />
                    <SPLIT distance="350" swimtime="00:06:08.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="349" reactiontime="+122" swimtime="00:03:13.25" resultid="3736" heatid="8095" lane="4" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.53" />
                    <SPLIT distance="100" swimtime="00:01:33.77" />
                    <SPLIT distance="150" swimtime="00:02:24.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="300" reactiontime="+132" swimtime="00:08:16.67" resultid="3737" heatid="8166" lane="1" entrytime="00:08:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.79" />
                    <SPLIT distance="100" swimtime="00:02:00.11" />
                    <SPLIT distance="150" swimtime="00:03:13.42" />
                    <SPLIT distance="200" swimtime="00:04:27.74" />
                    <SPLIT distance="250" swimtime="00:05:32.19" />
                    <SPLIT distance="300" swimtime="00:06:36.21" />
                    <SPLIT distance="350" swimtime="00:07:26.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-08-04" firstname="Wojciech" gender="M" lastname="Staruch" nation="POL" athleteid="3750">
              <RESULTS>
                <RESULT eventid="1075" points="443" reactiontime="+93" swimtime="00:03:32.86" resultid="3751" heatid="7947" lane="2" entrytime="00:03:35.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.36" />
                    <SPLIT distance="100" swimtime="00:01:44.94" />
                    <SPLIT distance="150" swimtime="00:02:43.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="438" reactiontime="+70" swimtime="00:00:39.42" resultid="3752" heatid="7964" lane="9" entrytime="00:00:39.12" />
                <RESULT eventid="1228" points="526" reactiontime="+83" swimtime="00:00:42.55" resultid="3753" heatid="8003" lane="1" entrytime="00:00:42.34" />
                <RESULT eventid="1258" points="390" reactiontime="+104" swimtime="00:03:52.22" resultid="3754" heatid="8015" lane="8" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.81" />
                    <SPLIT distance="100" swimtime="00:01:52.51" />
                    <SPLIT distance="150" swimtime="00:02:54.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="487" reactiontime="+80" swimtime="00:03:47.36" resultid="3755" heatid="8073" lane="2" entrytime="00:03:34.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.30" />
                    <SPLIT distance="100" swimtime="00:01:46.96" />
                    <SPLIT distance="150" swimtime="00:02:45.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="412" reactiontime="+77" swimtime="00:01:36.16" resultid="3756" heatid="8083" lane="9" entrytime="00:01:32.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="484" reactiontime="+86" swimtime="00:01:40.99" resultid="3757" heatid="8127" lane="2" entrytime="00:01:35.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="425" reactiontime="+118" swimtime="00:07:49.14" resultid="3758" heatid="8166" lane="8" entrytime="00:08:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.54" />
                    <SPLIT distance="100" swimtime="00:01:50.74" />
                    <SPLIT distance="150" swimtime="00:02:54.51" />
                    <SPLIT distance="200" swimtime="00:03:59.01" />
                    <SPLIT distance="250" swimtime="00:05:01.21" />
                    <SPLIT distance="300" swimtime="00:06:03.07" />
                    <SPLIT distance="350" swimtime="00:06:57.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-27" firstname="Wojciech" gender="M" lastname="Korpetta" nation="POL" athleteid="3726">
              <RESULTS>
                <RESULT eventid="1105" points="264" reactiontime="+133" swimtime="00:00:44.43" resultid="3727" heatid="7961" lane="4" />
                <RESULT eventid="1165" points="492" reactiontime="+127" swimtime="00:24:58.91" resultid="3728" heatid="8145" lane="4" entrytime="00:26:03.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.87" />
                    <SPLIT distance="100" swimtime="00:01:37.59" />
                    <SPLIT distance="150" swimtime="00:02:28.48" />
                    <SPLIT distance="200" swimtime="00:03:19.97" />
                    <SPLIT distance="250" swimtime="00:04:11.09" />
                    <SPLIT distance="300" swimtime="00:05:02.71" />
                    <SPLIT distance="350" swimtime="00:05:53.57" />
                    <SPLIT distance="400" swimtime="00:06:44.89" />
                    <SPLIT distance="450" swimtime="00:07:35.03" />
                    <SPLIT distance="500" swimtime="00:08:25.95" />
                    <SPLIT distance="550" swimtime="00:09:16.35" />
                    <SPLIT distance="600" swimtime="00:10:07.47" />
                    <SPLIT distance="650" swimtime="00:10:57.66" />
                    <SPLIT distance="700" swimtime="00:11:48.06" />
                    <SPLIT distance="750" swimtime="00:12:38.11" />
                    <SPLIT distance="800" swimtime="00:13:28.78" />
                    <SPLIT distance="850" swimtime="00:14:18.80" />
                    <SPLIT distance="900" swimtime="00:15:09.62" />
                    <SPLIT distance="950" swimtime="00:16:00.06" />
                    <SPLIT distance="1000" swimtime="00:16:50.21" />
                    <SPLIT distance="1050" swimtime="00:17:39.25" />
                    <SPLIT distance="1100" swimtime="00:18:29.48" />
                    <SPLIT distance="1150" swimtime="00:19:19.21" />
                    <SPLIT distance="1200" swimtime="00:20:09.31" />
                    <SPLIT distance="1250" swimtime="00:20:58.76" />
                    <SPLIT distance="1300" swimtime="00:21:48.30" />
                    <SPLIT distance="1350" swimtime="00:22:37.71" />
                    <SPLIT distance="1400" swimtime="00:23:26.92" />
                    <SPLIT distance="1450" swimtime="00:24:14.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="545" reactiontime="+72" swimtime="00:03:15.97" resultid="3729" heatid="8024" lane="3" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.50" />
                    <SPLIT distance="100" swimtime="00:01:36.37" />
                    <SPLIT distance="150" swimtime="00:02:26.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="492" reactiontime="+75" swimtime="00:01:31.14" resultid="3730" heatid="8038" lane="3" entrytime="00:01:32.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="432" reactiontime="+118" swimtime="00:03:00.01" resultid="3731" heatid="8093" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.11" />
                    <SPLIT distance="100" swimtime="00:01:26.78" />
                    <SPLIT distance="150" swimtime="00:02:14.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="472" reactiontime="+71" swimtime="00:00:41.71" resultid="3732" heatid="8111" lane="6" entrytime="00:00:41.17" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1614" reactiontime="+60" swimtime="00:02:50.95" resultid="3759" heatid="8133" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.36" />
                    <SPLIT distance="100" swimtime="00:01:33.70" />
                    <SPLIT distance="150" swimtime="00:02:13.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3726" number="1" reactiontime="+60" />
                    <RELAYPOSITION athleteid="3738" number="2" />
                    <RELAYPOSITION athleteid="3750" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="3743" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="LTU" clubid="6409" name="Kaisiadoriu p.k. &quot;PLAUKIAM&quot;">
          <CONTACT city="Vilnius" email="alex@gedwood.eu" name="Aleksandras Zamorskis" phone="+370 65609220" street="Fizikø 14-59" zip="VNO" />
          <ATHLETES>
            <ATHLETE birthdate="1971-04-22" firstname="Aleksandras" gender="M" lastname="Zamorskis" nation="LTU" athleteid="6410">
              <RESULTS>
                <RESULT eventid="1228" points="880" reactiontime="+67" swimtime="00:00:31.83" resultid="6411" heatid="8009" lane="7" entrytime="00:00:33.00" />
                <RESULT eventid="1402" points="882" reactiontime="+75" swimtime="00:02:37.28" resultid="6412" heatid="8077" lane="6" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.78" />
                    <SPLIT distance="100" swimtime="00:01:15.81" />
                    <SPLIT distance="150" swimtime="00:01:56.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="889" reactiontime="+60" swimtime="00:01:11.47" resultid="6413" heatid="8132" lane="8" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-01-14" firstname="Eimantas" gender="M" lastname="Frankonis" nation="LTU" athleteid="6414">
              <RESULTS>
                <RESULT eventid="1198" points="558" reactiontime="+77" swimtime="00:01:07.83" resultid="6415" heatid="7988" lane="8" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="553" reactiontime="+67" swimtime="00:03:07.22" resultid="6416" heatid="8076" lane="9" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.36" />
                    <SPLIT distance="100" swimtime="00:01:30.58" />
                    <SPLIT distance="150" swimtime="00:02:19.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="598" reactiontime="+75" swimtime="00:01:21.79" resultid="6417" heatid="8130" lane="6" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-05-01" firstname="Mindaugas" gender="M" lastname="Sakys" nation="LTU" athleteid="6427">
              <RESULTS>
                <RESULT eventid="1288" points="620" reactiontime="+72" swimtime="00:02:39.06" resultid="6428" heatid="8027" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.90" />
                    <SPLIT distance="100" swimtime="00:01:15.45" />
                    <SPLIT distance="150" swimtime="00:01:57.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="654" reactiontime="+78" swimtime="00:01:12.51" resultid="6429" heatid="8042" lane="9" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="540" reactiontime="+83" swimtime="00:00:34.98" resultid="6430" heatid="8115" lane="9" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-08-22" firstname="Gintas" gender="M" lastname="Kanapickas" nation="LTU" athleteid="6423">
              <RESULTS>
                <RESULT eventid="1198" points="533" reactiontime="+72" swimtime="00:01:11.13" resultid="6424" heatid="7986" lane="6" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="524" reactiontime="+86" swimtime="00:05:37.96" resultid="6425" heatid="8153" lane="2" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                    <SPLIT distance="100" swimtime="00:01:15.36" />
                    <SPLIT distance="150" swimtime="00:01:57.86" />
                    <SPLIT distance="200" swimtime="00:02:41.46" />
                    <SPLIT distance="250" swimtime="00:03:25.63" />
                    <SPLIT distance="300" swimtime="00:04:10.20" />
                    <SPLIT distance="350" swimtime="00:04:55.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="569" reactiontime="+80" swimtime="00:02:35.93" resultid="6426" heatid="8098" lane="4" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                    <SPLIT distance="100" swimtime="00:01:13.70" />
                    <SPLIT distance="150" swimtime="00:01:54.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-07-20" firstname="Raimondas" gender="M" lastname="Gincas" nation="LTU" athleteid="6418">
              <RESULTS>
                <RESULT eventid="1198" points="809" reactiontime="+71" swimtime="00:00:58.29" resultid="6419" heatid="7992" lane="6" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="804" reactiontime="+69" swimtime="00:00:26.43" resultid="6420" heatid="8064" lane="4" entrytime="00:00:26.00" />
                <RESULT eventid="1432" points="604" reactiontime="+69" swimtime="00:05:00.89" resultid="6421" heatid="8151" lane="6" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.08" />
                    <SPLIT distance="100" swimtime="00:01:09.97" />
                    <SPLIT distance="150" swimtime="00:01:47.78" />
                    <SPLIT distance="200" swimtime="00:02:26.41" />
                    <SPLIT distance="250" swimtime="00:03:04.89" />
                    <SPLIT distance="300" swimtime="00:03:43.92" />
                    <SPLIT distance="350" swimtime="00:04:22.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="703" reactiontime="+72" swimtime="00:02:13.24" resultid="6422" heatid="8102" lane="0" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.73" />
                    <SPLIT distance="100" swimtime="00:01:03.29" />
                    <SPLIT distance="150" swimtime="00:01:37.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1318" reactiontime="+70" swimtime="00:04:08.96" resultid="6431" heatid="8031" lane="2" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.81" />
                    <SPLIT distance="100" swimtime="00:00:58.52" />
                    <SPLIT distance="150" swimtime="00:01:29.14" />
                    <SPLIT distance="200" swimtime="00:02:05.34" />
                    <SPLIT distance="250" swimtime="00:02:35.61" />
                    <SPLIT distance="300" swimtime="00:03:08.43" />
                    <SPLIT distance="350" swimtime="00:03:37.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6410" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="6414" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="6427" number="3" reactiontime="+28" />
                    <RELAYPOSITION athleteid="6418" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="LTU" clubid="4703" name="Kauno Takas">
          <CONTACT city="Kaunas" email="abicka@takas.lt" internet="www.klubastakas.lt" name="Linas Kersevicius" phone="+37068780249" street="Lentvario g. 19" zip="44439" />
          <ATHLETES>
            <ATHLETE birthdate="1961-12-26" firstname="Arlandas Antanas" gender="M" lastname="Juodeska" nation="LTU" athleteid="4708">
              <RESULTS>
                <RESULT eventid="1075" points="576" reactiontime="+76" swimtime="00:02:53.26" resultid="4709" heatid="7950" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                    <SPLIT distance="100" swimtime="00:01:20.85" />
                    <SPLIT distance="150" swimtime="00:02:13.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="633" reactiontime="+74" swimtime="00:00:37.46" resultid="4710" heatid="8006" lane="9" entrytime="00:00:38.00" />
                <RESULT eventid="1288" points="643" reactiontime="+70" swimtime="00:02:52.14" resultid="4711" heatid="8026" lane="7" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                    <SPLIT distance="100" swimtime="00:01:23.99" />
                    <SPLIT distance="150" swimtime="00:02:09.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="618" reactiontime="+67" swimtime="00:01:17.29" resultid="4712" heatid="8040" lane="4" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="575" reactiontime="+79" swimtime="00:03:12.45" resultid="4713" heatid="8075" lane="1" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.15" />
                    <SPLIT distance="100" swimtime="00:01:34.59" />
                    <SPLIT distance="150" swimtime="00:02:24.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="765" reactiontime="+67" swimtime="00:00:33.37" resultid="4714" heatid="8114" lane="0" entrytime="00:00:34.00" />
                <RESULT eventid="1569" points="644" reactiontime="+73" swimtime="00:01:23.93" resultid="4715" heatid="8129" lane="6" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-06-18" firstname="Linas" gender="M" lastname="Kersevicius" nation="LTU" athleteid="4716">
              <RESULTS>
                <RESULT eventid="1075" points="576" reactiontime="+89" swimtime="00:02:39.14" resultid="4717" heatid="7952" lane="0" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                    <SPLIT distance="100" swimtime="00:01:13.92" />
                    <SPLIT distance="150" swimtime="00:02:01.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="673" reactiontime="+77" swimtime="00:02:34.75" resultid="4718" heatid="8028" lane="9" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                    <SPLIT distance="100" swimtime="00:01:14.14" />
                    <SPLIT distance="150" swimtime="00:01:54.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="728" reactiontime="+77" swimtime="00:01:09.97" resultid="4719" heatid="8042" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="707" reactiontime="+72" swimtime="00:00:31.98" resultid="4720" heatid="8116" lane="8" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02001" nation="POL" region="DOL" clubid="4268" name="Klub Sportowy REKIN Świebodzice" shortname="Klub Sportowy REKIN Świebodzic">
          <CONTACT city="Świebodzice" email="winiar182@wp.pl" internet="www.klubrekin.pl" name="WINIARCZYK Krzysztof" phone="606626274" state="DOL" street="Mieszka Starego 4" zip="58-160" />
          <ATHLETES>
            <ATHLETE birthdate="1982-11-09" firstname="Karol" gender="M" lastname="Żemier" nation="POL" athleteid="4293">
              <RESULTS>
                <RESULT eventid="1075" points="710" reactiontime="+78" swimtime="00:02:27.48" resultid="4294" heatid="7953" lane="1" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.98" />
                    <SPLIT distance="100" swimtime="00:01:06.39" />
                    <SPLIT distance="150" swimtime="00:01:50.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="732" reactiontime="+74" swimtime="00:00:27.75" resultid="4295" heatid="7971" lane="4" entrytime="00:00:27.90" entrycourse="SCM" />
                <RESULT eventid="1228" points="655" reactiontime="+74" swimtime="00:00:33.60" resultid="4296" heatid="8009" lane="1" entrytime="00:00:33.50" />
                <RESULT eventid="1258" points="621" reactiontime="+79" swimtime="00:02:35.14" resultid="4297" heatid="8017" lane="2" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                    <SPLIT distance="100" swimtime="00:01:06.14" />
                    <SPLIT distance="150" swimtime="00:01:46.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="692" reactiontime="+75" swimtime="00:00:26.28" resultid="4298" heatid="8064" lane="0" entrytime="00:00:26.20" />
                <RESULT eventid="1462" points="733" reactiontime="+79" swimtime="00:01:02.86" resultid="4299" heatid="8086" lane="9" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="683" reactiontime="+64" swimtime="00:00:29.54" resultid="4300" heatid="8117" lane="2" entrytime="00:00:29.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-04-16" firstname="Filip" gender="M" lastname="Żemier" nation="POL" athleteid="4287">
              <RESULTS>
                <RESULT eventid="1105" points="543" reactiontime="+68" swimtime="00:00:30.66" resultid="4288" heatid="7972" lane="9" entrytime="00:00:27.90" entrycourse="SCM" />
                <RESULT eventid="1198" points="534" reactiontime="+68" swimtime="00:01:02.64" resultid="4289" heatid="7992" lane="3" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="388" reactiontime="+67" swimtime="00:00:40.02" resultid="4290" heatid="8009" lane="0" entrytime="00:00:33.60" />
                <RESULT eventid="1372" points="636" reactiontime="+69" swimtime="00:00:27.03" resultid="4291" heatid="8064" lane="7" entrytime="00:00:26.10" />
                <RESULT eventid="1569" points="400" reactiontime="+72" swimtime="00:01:28.39" resultid="4292" heatid="8131" lane="0" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-12-22" firstname="Jacek" gender="M" lastname="Hankus" nation="POL" athleteid="4269">
              <RESULTS>
                <RESULT eventid="1105" points="723" reactiontime="+75" swimtime="00:00:27.93" resultid="4270" heatid="7972" lane="1" entrytime="00:00:27.50" entrycourse="SCM" />
                <RESULT eventid="1198" points="644" reactiontime="+73" swimtime="00:00:59.86" resultid="4271" heatid="7992" lane="8" entrytime="00:00:58.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="547" reactiontime="+74" swimtime="00:00:35.82" resultid="4272" heatid="8008" lane="4" entrytime="00:00:33.80" />
                <RESULT eventid="1342" points="659" reactiontime="+68" swimtime="00:01:08.07" resultid="4273" heatid="8043" lane="7" entrytime="00:01:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="642" reactiontime="+73" swimtime="00:00:26.83" resultid="4274" heatid="8064" lane="9" entrytime="00:00:26.20" />
                <RESULT eventid="1539" points="631" reactiontime="+61" swimtime="00:00:31.22" resultid="4275" heatid="8117" lane="8" entrytime="00:00:29.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-10-23" firstname="Piotr" gender="M" lastname="Tatarynowicz" nation="POL" athleteid="4276">
              <RESULTS>
                <RESULT eventid="1288" points="732" reactiontime="+68" swimtime="00:02:26.32" resultid="4277" heatid="8028" lane="7" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.52" />
                    <SPLIT distance="100" swimtime="00:01:09.64" />
                    <SPLIT distance="150" swimtime="00:01:47.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="633" reactiontime="+69" swimtime="00:01:05.86" resultid="4278" heatid="8043" lane="3" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="660" reactiontime="+69" swimtime="00:00:29.88" resultid="4279" heatid="8117" lane="7" entrytime="00:00:29.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-06-21" firstname="Alfred" gender="M" lastname="Żemier" nation="POL" athleteid="4280">
              <RESULTS>
                <RESULT eventid="1075" points="597" reactiontime="+79" swimtime="00:02:36.27" resultid="4281" heatid="7953" lane="0" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.27" />
                    <SPLIT distance="100" swimtime="00:01:10.72" />
                    <SPLIT distance="150" swimtime="00:01:58.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="642" reactiontime="+78" swimtime="00:00:58.91" resultid="4282" heatid="7993" lane="0" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="499" reactiontime="+63" swimtime="00:00:36.78" resultid="4283" heatid="8009" lane="9" entrytime="00:00:33.70" />
                <RESULT eventid="1342" points="546" reactiontime="+73" swimtime="00:01:09.16" resultid="4284" heatid="8043" lane="1" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="692" reactiontime="+77" swimtime="00:00:26.28" resultid="4285" heatid="8065" lane="0" entrytime="00:00:26.00" />
                <RESULT eventid="1539" points="583" reactiontime="+64" swimtime="00:00:31.14" resultid="4286" heatid="8117" lane="9" entrytime="00:00:29.90" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" name="Rekin Świebodzice" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1318" reactiontime="+75" swimtime="00:03:56.13" resultid="4301" heatid="8031" lane="6" entrytime="00:03:59.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.78" />
                    <SPLIT distance="100" swimtime="00:00:58.70" />
                    <SPLIT distance="150" swimtime="00:01:26.20" />
                    <SPLIT distance="200" swimtime="00:01:57.37" />
                    <SPLIT distance="250" swimtime="00:02:24.16" />
                    <SPLIT distance="300" swimtime="00:02:55.24" />
                    <SPLIT distance="350" swimtime="00:03:22.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4293" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="4287" number="2" reactiontime="+67" />
                    <RELAYPOSITION athleteid="4269" number="3" reactiontime="+25" />
                    <RELAYPOSITION athleteid="4280" number="4" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="501013" nation="POL" region="WAR" clubid="3572" name="KP Victory Masters Elbląg">
          <CONTACT city="Elbląg" email="waldi-m@wp.pl" name="Maciesza Waldemar" phone="608338265" state="WAR-M" street="ul. Bema 42" zip="82-300" />
          <ATHLETES>
            <ATHLETE birthdate="1965-12-25" firstname="Waldemar" gender="M" lastname="Maciesza" nation="POL" athleteid="3573">
              <RESULTS>
                <RESULT eventid="1198" points="390" reactiontime="+104" swimtime="00:01:18.90" resultid="3574" heatid="7983" lane="5" entrytime="00:01:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="384" reactiontime="+90" swimtime="00:00:44.27" resultid="3575" heatid="8002" lane="6" entrytime="00:00:45.00" entrycourse="LCM" />
                <RESULT eventid="1402" points="328" reactiontime="+76" swimtime="00:03:51.93" resultid="3576" heatid="8071" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.67" />
                    <SPLIT distance="100" swimtime="00:01:50.58" />
                    <SPLIT distance="150" swimtime="00:02:51.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="298" reactiontime="+101" swimtime="00:03:13.46" resultid="3577" heatid="8095" lane="1" entrytime="00:03:15.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.66" />
                    <SPLIT distance="100" swimtime="00:01:34.93" />
                    <SPLIT distance="150" swimtime="00:02:25.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="339" reactiontime="+93" swimtime="00:01:43.95" resultid="3578" heatid="8126" lane="6" entrytime="00:01:42.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PŁYWAK" nation="POL" region="WAR" clubid="3579" name="KPiRS &quot;PŁYWAK&quot; Płock">
          <CONTACT city="Płock" email="pawel.powichrowski@wp.pl" name="Powichrowski Paweł" phone="603694397" state="MAZ" street="Wiatraki 11 b" zip="09-402" />
          <ATHLETES>
            <ATHLETE birthdate="1995-04-28" firstname="Karolina" gender="F" lastname="Kowalska" nation="POL" athleteid="3588">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="3589" heatid="7942" lane="4" entrytime="00:03:20.00" />
                <RESULT eventid="1090" status="DNS" swimtime="00:00:00.00" resultid="3590" heatid="7959" lane="0" entrytime="00:00:35.00" />
                <RESULT eventid="1181" status="DNS" swimtime="00:00:00.00" resultid="3591" heatid="7978" lane="0" entrytime="00:01:12.00" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="3592" heatid="8021" lane="3" entrytime="00:02:40.00" />
                <RESULT eventid="1326" status="DNS" swimtime="00:00:00.00" resultid="3593" heatid="8032" lane="7" />
                <RESULT eventid="1357" status="DNS" swimtime="00:00:00.00" resultid="3594" heatid="8048" lane="3" entrytime="00:00:32.00" />
                <RESULT eventid="1554" status="DNS" swimtime="00:00:00.00" resultid="3595" heatid="8121" lane="3" entrytime="00:01:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-09" firstname="Piotr" gender="M" lastname="Mikuła" nation="POL" athleteid="3580">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="3581" heatid="7953" lane="8" entrytime="00:02:25.00" />
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="3582" heatid="7969" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="3583" heatid="7980" lane="5" />
                <RESULT eventid="1228" status="DNS" swimtime="00:00:00.00" resultid="3584" heatid="8010" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="1372" status="DNS" swimtime="00:00:00.00" resultid="3585" heatid="8065" lane="5" entrytime="00:00:24.00" />
                <RESULT eventid="1509" status="DNS" swimtime="00:00:00.00" resultid="3587" heatid="8101" lane="6" entrytime="00:02:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-07-04" firstname="Agata" gender="F" lastname="Olejniczak" nation="POL" athleteid="3596">
              <RESULTS>
                <RESULT eventid="1058" points="552" reactiontime="+90" swimtime="00:02:58.58" resultid="3597" heatid="7943" lane="9" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                    <SPLIT distance="100" swimtime="00:01:27.05" />
                    <SPLIT distance="150" swimtime="00:02:18.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="599" reactiontime="+89" swimtime="00:00:39.84" resultid="3598" heatid="7999" lane="2" entrytime="00:00:39.00" />
                <RESULT eventid="1273" points="424" reactiontime="+89" swimtime="00:03:12.86" resultid="3599" heatid="8021" lane="5" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.27" />
                    <SPLIT distance="100" swimtime="00:01:30.14" />
                    <SPLIT distance="150" swimtime="00:02:20.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="760" reactiontime="+88" swimtime="00:00:29.17" resultid="3600" heatid="8050" lane="0" entrytime="00:00:29.00" />
                <RESULT eventid="1387" points="501" reactiontime="+93" swimtime="00:03:18.84" resultid="3601" heatid="8069" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.60" />
                    <SPLIT distance="100" swimtime="00:01:35.30" />
                    <SPLIT distance="150" swimtime="00:02:27.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="571" reactiontime="+91" swimtime="00:01:29.16" resultid="3602" heatid="8122" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-06-30" firstname="Łukasz" gender="M" lastname="Szypryt" nation="POL" athleteid="3603">
              <RESULTS>
                <RESULT eventid="1075" points="410" reactiontime="+82" swimtime="00:02:49.46" resultid="3604" heatid="7951" lane="7" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.94" />
                    <SPLIT distance="100" swimtime="00:01:15.39" />
                    <SPLIT distance="150" swimtime="00:02:03.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="523" reactiontime="+79" swimtime="00:00:36.35" resultid="3605" heatid="8010" lane="7" entrytime="00:00:32.00" />
                <RESULT eventid="1288" points="365" reactiontime="+83" swimtime="00:02:53.23" resultid="3606" heatid="8028" lane="0" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.41" />
                    <SPLIT distance="100" swimtime="00:01:20.08" />
                    <SPLIT distance="150" swimtime="00:02:04.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="431" reactiontime="+81" swimtime="00:01:18.40" resultid="3607" heatid="8042" lane="3" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="470" reactiontime="+85" swimtime="00:03:08.24" resultid="3608" heatid="8076" lane="4" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.81" />
                    <SPLIT distance="100" swimtime="00:01:31.88" />
                    <SPLIT distance="150" swimtime="00:02:20.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="366" reactiontime="+85" swimtime="00:01:30.40" resultid="3609" heatid="8132" lane="7" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="438" reactiontime="+86" swimtime="00:06:15.63" resultid="3610" heatid="8163" lane="4" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.31" />
                    <SPLIT distance="100" swimtime="00:01:24.42" />
                    <SPLIT distance="150" swimtime="00:02:14.84" />
                    <SPLIT distance="200" swimtime="00:03:05.01" />
                    <SPLIT distance="250" swimtime="00:03:52.97" />
                    <SPLIT distance="300" swimtime="00:04:43.25" />
                    <SPLIT distance="350" swimtime="00:05:29.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01910" nation="POL" region="POM" clubid="3295" name="KS Delfin Gdynia">
          <ATHLETES>
            <ATHLETE birthdate="1971-11-04" firstname="Jakub" gender="M" lastname="Mańczak" nation="POL" license="101910200065" athleteid="3296">
              <RESULTS>
                <RESULT eventid="1105" points="657" reactiontime="+71" swimtime="00:00:29.78" resultid="3297" heatid="7970" lane="8" entrytime="00:00:29.50" />
                <RESULT eventid="1258" points="469" reactiontime="+86" swimtime="00:02:50.29" resultid="3298" heatid="8016" lane="4" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.87" />
                    <SPLIT distance="100" swimtime="00:01:18.22" />
                    <SPLIT distance="150" swimtime="00:02:05.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="699" reactiontime="+70" swimtime="00:00:27.69" resultid="3299" heatid="8062" lane="2" entrytime="00:00:27.60" />
                <RESULT eventid="1462" points="632" reactiontime="+72" swimtime="00:01:08.37" resultid="3300" heatid="8085" lane="8" entrytime="00:01:09.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="EXOBO" nation="POL" region="WIE" clubid="6436" name="Ks Extreme Team Oborniki">
          <CONTACT city="OBORNIKI" email="janwol@poczta.onet.pl" name="WOLNIEWICZ" phone="791064667" state="WIE" street="CZARNKOWSKA 84" zip="64-600" />
          <ATHLETES>
            <ATHLETE birthdate="1948-12-22" firstname="Janusz" gender="M" lastname="Wolniewicz" nation="POL" athleteid="6437">
              <RESULTS>
                <RESULT eventid="1165" points="340" reactiontime="+109" swimtime="00:30:01.29" resultid="6438" heatid="8145" lane="7" entrytime="00:28:22.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.71" />
                    <SPLIT distance="100" swimtime="00:01:43.13" />
                    <SPLIT distance="150" swimtime="00:02:40.28" />
                    <SPLIT distance="200" swimtime="00:03:38.63" />
                    <SPLIT distance="250" swimtime="00:04:38.61" />
                    <SPLIT distance="300" swimtime="00:05:37.93" />
                    <SPLIT distance="350" swimtime="00:06:37.25" />
                    <SPLIT distance="400" swimtime="00:07:37.42" />
                    <SPLIT distance="450" swimtime="00:08:37.84" />
                    <SPLIT distance="500" swimtime="00:09:37.04" />
                    <SPLIT distance="550" swimtime="00:10:36.55" />
                    <SPLIT distance="600" swimtime="00:11:35.83" />
                    <SPLIT distance="650" swimtime="00:12:35.18" />
                    <SPLIT distance="700" swimtime="00:13:35.14" />
                    <SPLIT distance="750" swimtime="00:14:35.35" />
                    <SPLIT distance="800" swimtime="00:15:35.67" />
                    <SPLIT distance="850" swimtime="00:16:36.84" />
                    <SPLIT distance="900" swimtime="00:17:38.30" />
                    <SPLIT distance="950" swimtime="00:18:40.43" />
                    <SPLIT distance="1000" swimtime="00:19:42.78" />
                    <SPLIT distance="1050" swimtime="00:20:45.32" />
                    <SPLIT distance="1100" swimtime="00:21:47.30" />
                    <SPLIT distance="1150" swimtime="00:22:50.66" />
                    <SPLIT distance="1200" swimtime="00:23:52.75" />
                    <SPLIT distance="1250" swimtime="00:24:53.69" />
                    <SPLIT distance="1300" swimtime="00:25:56.89" />
                    <SPLIT distance="1350" swimtime="00:26:59.82" />
                    <SPLIT distance="1400" swimtime="00:28:03.04" />
                    <SPLIT distance="1450" swimtime="00:29:03.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="467" reactiontime="+96" swimtime="00:01:25.05" resultid="6439" heatid="7983" lane="1" entrytime="00:01:23.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="346" reactiontime="+90" swimtime="00:07:37.47" resultid="6440" heatid="8155" lane="7" entrytime="00:06:59.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.87" />
                    <SPLIT distance="100" swimtime="00:01:42.40" />
                    <SPLIT distance="150" swimtime="00:02:41.68" />
                    <SPLIT distance="200" swimtime="00:03:41.61" />
                    <SPLIT distance="250" swimtime="00:04:41.55" />
                    <SPLIT distance="300" swimtime="00:05:42.48" />
                    <SPLIT distance="350" swimtime="00:06:41.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="396" reactiontime="+98" swimtime="00:03:24.92" resultid="6441" heatid="8096" lane="8" entrytime="00:03:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.81" />
                    <SPLIT distance="100" swimtime="00:01:35.58" />
                    <SPLIT distance="150" swimtime="00:02:30.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAPOL" nation="POL" region="DOL" clubid="3616" name="KS Masters Polkowice">
          <CONTACT city="Polkowice" email="bogdan.jawor@gmail.com" name="Jawor Bogdan" phone="519102742" state="DOL" street="ul.Kolejowa 6/5" zip="59-100" />
          <ATHLETES>
            <ATHLETE birthdate="1968-01-02" firstname="Pavlo" gender="M" lastname="Vechirko" nation="POL" athleteid="3629">
              <RESULTS>
                <RESULT eventid="1228" points="469" swimtime="00:00:38.48" resultid="3630" heatid="8007" lane="0" entrytime="00:00:37.00" entrycourse="LCM" />
                <RESULT eventid="1288" points="524" reactiontime="+82" swimtime="00:02:55.65" resultid="3631" heatid="8027" lane="9" entrytime="00:02:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.54" />
                    <SPLIT distance="100" swimtime="00:01:24.03" />
                    <SPLIT distance="150" swimtime="00:02:09.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="495" reactiontime="+79" swimtime="00:01:20.73" resultid="3632" heatid="8041" lane="2" entrytime="00:01:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" status="DNS" swimtime="00:00:00.00" resultid="3633" heatid="8075" lane="4" entrytime="00:03:05.00" entrycourse="LCM" />
                <RESULT eventid="1539" points="507" reactiontime="+82" swimtime="00:00:36.66" resultid="3634" heatid="8113" lane="6" entrytime="00:00:35.00" entrycourse="LCM" />
                <RESULT eventid="1569" points="484" reactiontime="+101" swimtime="00:01:27.73" resultid="3635" heatid="8130" lane="9" entrytime="00:01:24.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-04-23" firstname="Bogdan" gender="M" lastname="Jawor" nation="POL" athleteid="3644">
              <RESULTS>
                <RESULT eventid="1075" points="245" reactiontime="+95" swimtime="00:04:24.65" resultid="3645" heatid="7945" lane="3" entrytime="00:04:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.28" />
                    <SPLIT distance="100" swimtime="00:02:04.67" />
                    <SPLIT distance="150" swimtime="00:03:20.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="133" reactiontime="+95" swimtime="00:00:59.74" resultid="3646" heatid="7962" lane="5" entrytime="00:00:53.00" entrycourse="LCM" />
                <RESULT eventid="1228" points="293" reactiontime="+99" swimtime="00:00:54.57" resultid="3647" heatid="8001" lane="9" entrytime="00:00:54.00" entrycourse="LCM" />
                <RESULT eventid="1288" points="267" reactiontime="+92" swimtime="00:04:09.85" resultid="3648" heatid="8023" lane="7" entrytime="00:04:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.73" />
                    <SPLIT distance="100" swimtime="00:02:00.93" />
                    <SPLIT distance="150" swimtime="00:03:06.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="267" reactiontime="+85" swimtime="00:01:54.54" resultid="3649" heatid="8037" lane="8" entrytime="00:02:07.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="306" reactiontime="+107" swimtime="00:04:41.14" resultid="3650" heatid="8071" lane="5" entrytime="00:04:26.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.14" />
                    <SPLIT distance="100" swimtime="00:02:14.81" />
                    <SPLIT distance="150" swimtime="00:03:29.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="262" reactiontime="+98" swimtime="00:00:52.33" resultid="3651" heatid="8109" lane="8" entrytime="00:01:00.00" entrycourse="LCM" />
                <RESULT eventid="1569" points="277" reactiontime="+100" swimtime="00:02:06.21" resultid="3652" heatid="8125" lane="6" entrytime="00:02:03.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-05-30" firstname="Grażyna" gender="F" lastname="Grzegorzewska" nation="POL" athleteid="3621">
              <RESULTS>
                <RESULT eventid="1090" points="234" reactiontime="+94" swimtime="00:00:56.84" resultid="3622" heatid="7955" lane="7" entrytime="00:00:56.00" entrycourse="LCM" />
                <RESULT eventid="1120" points="430" reactiontime="+106" swimtime="00:15:36.60" resultid="3623" heatid="8137" lane="0" entrytime="00:15:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.05" />
                    <SPLIT distance="100" swimtime="00:01:47.55" />
                    <SPLIT distance="150" swimtime="00:02:47.16" />
                    <SPLIT distance="200" swimtime="00:03:47.54" />
                    <SPLIT distance="250" swimtime="00:04:47.04" />
                    <SPLIT distance="300" swimtime="00:05:46.55" />
                    <SPLIT distance="350" swimtime="00:06:46.04" />
                    <SPLIT distance="400" swimtime="00:07:45.10" />
                    <SPLIT distance="450" swimtime="00:08:44.79" />
                    <SPLIT distance="500" swimtime="00:09:44.23" />
                    <SPLIT distance="550" swimtime="00:10:44.16" />
                    <SPLIT distance="600" swimtime="00:11:43.93" />
                    <SPLIT distance="650" swimtime="00:12:43.52" />
                    <SPLIT distance="700" swimtime="00:13:43.33" />
                    <SPLIT distance="750" swimtime="00:14:42.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="391" reactiontime="+91" swimtime="00:01:36.11" resultid="3624" heatid="7974" lane="6" entrytime="00:01:35.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="459" reactiontime="+83" swimtime="00:00:40.89" resultid="3625" heatid="8045" lane="6" entrytime="00:00:42.00" entrycourse="LCM" />
                <RESULT eventid="1417" points="449" reactiontime="+96" swimtime="00:07:35.45" resultid="3626" heatid="8149" lane="0" entrytime="00:07:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.08" />
                    <SPLIT distance="100" swimtime="00:01:43.97" />
                    <SPLIT distance="150" swimtime="00:02:42.14" />
                    <SPLIT distance="200" swimtime="00:03:41.26" />
                    <SPLIT distance="250" swimtime="00:04:39.87" />
                    <SPLIT distance="300" swimtime="00:05:39.95" />
                    <SPLIT distance="350" swimtime="00:06:39.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="406" reactiontime="+95" swimtime="00:03:34.55" resultid="3627" heatid="8088" lane="0" entrytime="00:03:35.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.00" />
                    <SPLIT distance="100" swimtime="00:01:39.24" />
                    <SPLIT distance="150" swimtime="00:02:37.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="325" reactiontime="+82" swimtime="00:00:58.36" resultid="3628" heatid="8104" lane="8" entrytime="00:00:56.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-05-26" firstname="Zygmunt" gender="M" lastname="Pawlaczek" nation="POL" athleteid="3636">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="3637" heatid="7945" lane="5" entrytime="00:04:12.00" entrycourse="LCM" />
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="3638" heatid="7982" lane="3" entrytime="00:01:28.00" entrycourse="LCM" />
                <RESULT eventid="1228" status="DNS" swimtime="00:00:00.00" resultid="3639" heatid="8001" lane="2" entrytime="00:00:50.00" entrycourse="LCM" />
                <RESULT eventid="1342" status="DNS" swimtime="00:00:00.00" resultid="3640" heatid="8037" lane="5" entrytime="00:01:55.00" entrycourse="LCM" />
                <RESULT eventid="1372" status="DNS" swimtime="00:00:00.00" resultid="3641" heatid="8053" lane="2" entrytime="00:00:38.00" entrycourse="LCM" />
                <RESULT eventid="1509" status="DNS" swimtime="00:00:00.00" resultid="3642" heatid="8094" lane="4" entrytime="00:03:30.00" entrycourse="LCM" />
                <RESULT eventid="1539" status="DNS" swimtime="00:00:00.00" resultid="3643" heatid="8110" lane="6" entrytime="00:00:47.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WIE" nation="POL" region="WIE" clubid="3653" name="KS Warta Poznań">
          <CONTACT city="POZNAŃ" email="jacek.thiem@gmail.com" name="THIEM JACEK" phone="502499565" state="WIE" street="OS. DĘBINA 19 M 34" zip="61-450" />
          <ATHLETES>
            <ATHLETE birthdate="1969-07-07" firstname="Elżbieta" gender="F" lastname="Krakowiak" nation="POL" license="100115600356" athleteid="3663">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1357" points="870" reactiontime="+85" swimtime="00:00:29.69" resultid="3664" heatid="8049" lane="2" entrytime="00:00:31.00" />
                <RESULT eventid="1417" points="779" reactiontime="+90" swimtime="00:05:09.00" resultid="3665" heatid="8147" lane="2" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                    <SPLIT distance="100" swimtime="00:01:12.57" />
                    <SPLIT distance="150" swimtime="00:01:51.00" />
                    <SPLIT distance="200" swimtime="00:02:30.22" />
                    <SPLIT distance="250" swimtime="00:03:09.54" />
                    <SPLIT distance="300" swimtime="00:03:49.71" />
                    <SPLIT distance="350" swimtime="00:04:29.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="832" reactiontime="+89" swimtime="00:02:24.46" resultid="3666" heatid="8091" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                    <SPLIT distance="100" swimtime="00:01:09.58" />
                    <SPLIT distance="150" swimtime="00:01:47.21" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1584" points="826" reactiontime="+91" swimtime="00:05:54.47" resultid="3667" heatid="8159" lane="2" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                    <SPLIT distance="100" swimtime="00:01:19.30" />
                    <SPLIT distance="150" swimtime="00:02:05.77" />
                    <SPLIT distance="200" swimtime="00:02:51.65" />
                    <SPLIT distance="250" swimtime="00:03:43.15" />
                    <SPLIT distance="300" swimtime="00:04:35.17" />
                    <SPLIT distance="350" swimtime="00:05:15.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-22" firstname="Małgorzata" gender="F" lastname="Putowska" nation="POL" athleteid="3668">
              <RESULTS>
                <RESULT eventid="1090" points="274" reactiontime="+79" swimtime="00:00:46.55" resultid="3669" heatid="7955" lane="4" entrytime="00:00:49.53" />
                <RESULT eventid="1213" points="515" reactiontime="+86" swimtime="00:00:47.08" resultid="3670" heatid="7996" lane="6" entrytime="00:00:46.44" />
                <RESULT eventid="1273" points="320" reactiontime="+90" swimtime="00:04:03.92" resultid="3671" heatid="8019" lane="0" entrytime="00:03:58.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.49" />
                    <SPLIT distance="100" swimtime="00:01:58.12" />
                    <SPLIT distance="150" swimtime="00:03:01.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="327" reactiontime="+69" swimtime="00:01:49.42" resultid="3672" heatid="8033" lane="1" entrytime="00:01:47.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1387" points="435" reactiontime="+87" swimtime="00:04:01.66" resultid="3673" heatid="8067" lane="4" entrytime="00:03:53.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.69" />
                    <SPLIT distance="100" swimtime="00:01:54.97" />
                    <SPLIT distance="150" swimtime="00:02:59.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="413" reactiontime="+78" swimtime="00:01:52.08" resultid="3674" heatid="8120" lane="6" entrytime="00:01:44.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-07-23" firstname="Przemysław" gender="M" lastname="Kuca" nation="POL" license="S00115200198" athleteid="3703">
              <RESULTS>
                <RESULT eventid="1075" points="880" reactiontime="+67" swimtime="00:02:15.22" resultid="3704" heatid="7953" lane="4" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.88" />
                    <SPLIT distance="100" swimtime="00:01:04.49" />
                    <SPLIT distance="150" swimtime="00:01:45.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="756" reactiontime="+69" swimtime="00:00:27.71" resultid="3705" heatid="7972" lane="0" entrytime="00:00:27.66" />
                <RESULT eventid="1198" points="822" reactiontime="+72" swimtime="00:00:55.20" resultid="3706" heatid="7993" lane="6" entrytime="00:00:55.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="889" swimtime="00:02:11.06" resultid="3707" heatid="8017" lane="4" entrytime="00:02:10.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.99" />
                    <SPLIT distance="100" swimtime="00:01:02.09" />
                    <SPLIT distance="150" swimtime="00:01:36.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="743" reactiontime="+67" swimtime="00:04:23.76" resultid="3708" heatid="8151" lane="4" entrytime="00:04:23.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.27" />
                    <SPLIT distance="100" swimtime="00:01:01.82" />
                    <SPLIT distance="150" swimtime="00:01:35.01" />
                    <SPLIT distance="200" swimtime="00:02:09.05" />
                    <SPLIT distance="250" swimtime="00:02:42.90" />
                    <SPLIT distance="300" swimtime="00:03:17.53" />
                    <SPLIT distance="350" swimtime="00:03:51.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="866" reactiontime="+70" swimtime="00:00:59.23" resultid="3709" heatid="8086" lane="5" entrytime="00:00:58.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="831" reactiontime="+70" swimtime="00:02:03.01" resultid="3710" heatid="8102" lane="4" entrytime="00:02:04.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.02" />
                    <SPLIT distance="100" swimtime="00:00:59.13" />
                    <SPLIT distance="150" swimtime="00:01:31.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="860" reactiontime="+73" swimtime="00:04:54.13" resultid="3711" heatid="8162" lane="4" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.71" />
                    <SPLIT distance="100" swimtime="00:01:02.30" />
                    <SPLIT distance="150" swimtime="00:01:42.41" />
                    <SPLIT distance="200" swimtime="00:02:21.20" />
                    <SPLIT distance="250" swimtime="00:03:04.14" />
                    <SPLIT distance="300" swimtime="00:03:48.22" />
                    <SPLIT distance="350" swimtime="00:04:21.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-05-01" firstname="Kevin" gender="M" lastname="Mrotek" nation="POL" athleteid="3712">
              <RESULTS>
                <RESULT eventid="1075" points="521" swimtime="00:02:41.02" resultid="3713" heatid="7952" lane="9" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.40" />
                    <SPLIT distance="100" swimtime="00:01:12.50" />
                    <SPLIT distance="150" swimtime="00:02:01.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="562" reactiontime="+60" swimtime="00:00:30.58" resultid="3714" heatid="7970" lane="9" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-02" firstname="Paweł" gender="M" lastname="Olszewski" nation="POL" license="100115700350" athleteid="3697">
              <RESULTS>
                <RESULT eventid="1105" points="763" reactiontime="+76" swimtime="00:00:30.40" resultid="3698" heatid="7967" lane="5" entrytime="00:00:32.50" />
                <RESULT eventid="1198" points="858" reactiontime="+79" swimtime="00:01:00.70" resultid="3699" heatid="7990" lane="6" entrytime="00:01:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="909" reactiontime="+78" swimtime="00:02:13.42" resultid="3701" heatid="8101" lane="2" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.45" />
                    <SPLIT distance="100" swimtime="00:01:04.21" />
                    <SPLIT distance="150" swimtime="00:01:38.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="672" reactiontime="+65" swimtime="00:00:34.83" resultid="3702" heatid="8114" lane="1" entrytime="00:00:34.00" />
                <RESULT eventid="1432" points="794" reactiontime="+84" swimtime="00:04:54.31" resultid="8289" heatid="8156" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                    <SPLIT distance="100" swimtime="00:01:11.29" />
                    <SPLIT distance="150" swimtime="00:01:48.96" />
                    <SPLIT distance="200" swimtime="00:02:26.98" />
                    <SPLIT distance="250" swimtime="00:03:04.31" />
                    <SPLIT distance="300" swimtime="00:03:41.65" />
                    <SPLIT distance="350" swimtime="00:04:18.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-02-17" firstname="Jacek" gender="M" lastname="Thiem" nation="POL" license="100115700345" athleteid="3684">
              <RESULTS>
                <RESULT eventid="1135" points="352" reactiontime="+107" swimtime="00:13:17.81" resultid="3685" heatid="8140" lane="1" entrytime="00:13:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.97" />
                    <SPLIT distance="100" swimtime="00:01:31.70" />
                    <SPLIT distance="150" swimtime="00:02:21.26" />
                    <SPLIT distance="200" swimtime="00:03:11.78" />
                    <SPLIT distance="250" swimtime="00:04:02.95" />
                    <SPLIT distance="300" swimtime="00:04:54.09" />
                    <SPLIT distance="350" swimtime="00:05:45.54" />
                    <SPLIT distance="400" swimtime="00:06:37.52" />
                    <SPLIT distance="450" swimtime="00:07:28.97" />
                    <SPLIT distance="500" swimtime="00:08:20.87" />
                    <SPLIT distance="550" swimtime="00:09:12.61" />
                    <SPLIT distance="600" swimtime="00:10:03.81" />
                    <SPLIT distance="650" swimtime="00:10:54.77" />
                    <SPLIT distance="700" swimtime="00:11:45.39" />
                    <SPLIT distance="750" swimtime="00:12:33.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="423" reactiontime="+108" swimtime="00:03:21.79" resultid="3686" heatid="8016" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.83" />
                    <SPLIT distance="100" swimtime="00:01:31.43" />
                    <SPLIT distance="150" swimtime="00:02:24.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="425" reactiontime="+105" swimtime="00:01:24.68" resultid="3687" heatid="8083" lane="3" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="406" reactiontime="+106" swimtime="00:02:54.49" resultid="3688" heatid="8096" lane="6" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                    <SPLIT distance="100" swimtime="00:01:26.04" />
                    <SPLIT distance="150" swimtime="00:02:11.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="359" reactiontime="+111" swimtime="00:07:28.18" resultid="3689" heatid="8166" lane="3" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.06" />
                    <SPLIT distance="100" swimtime="00:01:40.92" />
                    <SPLIT distance="150" swimtime="00:02:44.45" />
                    <SPLIT distance="200" swimtime="00:03:47.18" />
                    <SPLIT distance="250" swimtime="00:04:50.05" />
                    <SPLIT distance="300" swimtime="00:05:52.54" />
                    <SPLIT distance="350" swimtime="00:06:41.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-05-08" firstname="Anna" gender="F" lastname="Kotecka" nation="POL" license="100115600357" athleteid="3690">
              <RESULTS>
                <RESULT eventid="1150" points="683" swimtime="00:24:57.73" resultid="3691" heatid="8142" lane="2" entrytime="00:30:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.27" />
                    <SPLIT distance="100" swimtime="00:01:32.20" />
                    <SPLIT distance="150" swimtime="00:02:21.31" />
                    <SPLIT distance="200" swimtime="00:03:10.63" />
                    <SPLIT distance="250" swimtime="00:04:00.36" />
                    <SPLIT distance="300" swimtime="00:04:49.87" />
                    <SPLIT distance="350" swimtime="00:05:39.79" />
                    <SPLIT distance="400" swimtime="00:06:30.56" />
                    <SPLIT distance="450" swimtime="00:07:20.34" />
                    <SPLIT distance="500" swimtime="00:08:10.37" />
                    <SPLIT distance="550" swimtime="00:09:00.58" />
                    <SPLIT distance="600" swimtime="00:09:51.40" />
                    <SPLIT distance="650" swimtime="00:10:42.16" />
                    <SPLIT distance="700" swimtime="00:11:32.89" />
                    <SPLIT distance="750" swimtime="00:12:22.65" />
                    <SPLIT distance="800" swimtime="00:13:13.19" />
                    <SPLIT distance="850" swimtime="00:14:03.33" />
                    <SPLIT distance="900" swimtime="00:14:53.77" />
                    <SPLIT distance="950" swimtime="00:15:44.38" />
                    <SPLIT distance="1000" swimtime="00:16:34.67" />
                    <SPLIT distance="1050" swimtime="00:17:24.23" />
                    <SPLIT distance="1100" swimtime="00:18:14.37" />
                    <SPLIT distance="1150" swimtime="00:19:05.20" />
                    <SPLIT distance="1200" swimtime="00:19:55.97" />
                    <SPLIT distance="1250" swimtime="00:20:46.78" />
                    <SPLIT distance="1300" swimtime="00:21:37.88" />
                    <SPLIT distance="1350" swimtime="00:22:28.17" />
                    <SPLIT distance="1400" swimtime="00:23:19.20" />
                    <SPLIT distance="1450" swimtime="00:24:09.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="392" swimtime="00:01:27.71" resultid="3692" heatid="7975" lane="9" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="391" reactiontime="+87" swimtime="00:01:43.07" resultid="3693" heatid="8033" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="406" swimtime="00:06:32.92" resultid="3694" heatid="8148" lane="2" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.27" />
                    <SPLIT distance="100" swimtime="00:01:31.66" />
                    <SPLIT distance="150" swimtime="00:02:20.86" />
                    <SPLIT distance="200" swimtime="00:03:12.19" />
                    <SPLIT distance="250" swimtime="00:04:02.99" />
                    <SPLIT distance="300" swimtime="00:04:54.16" />
                    <SPLIT distance="350" swimtime="00:05:44.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="394" swimtime="00:03:08.32" resultid="3695" heatid="8089" lane="6" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.51" />
                    <SPLIT distance="100" swimtime="00:01:28.75" />
                    <SPLIT distance="150" swimtime="00:02:18.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="354" reactiontime="+104" swimtime="00:00:48.56" resultid="3696" heatid="8105" lane="9" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-07-02" firstname="Tomasz" gender="M" lastname="Tomaszewski" nation="POL" athleteid="3675">
              <RESULTS>
                <RESULT eventid="1288" points="564" reactiontime="+80" swimtime="00:02:39.65" resultid="3676" heatid="8027" lane="2" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                    <SPLIT distance="100" swimtime="00:01:13.46" />
                    <SPLIT distance="150" swimtime="00:01:55.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="547" reactiontime="+71" swimtime="00:01:09.11" resultid="3677" heatid="8042" lane="8" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="579" reactiontime="+65" swimtime="00:00:31.21" resultid="3678" heatid="8116" lane="2" entrytime="00:00:30.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-26" firstname="Stanisław" gender="M" lastname="Kaczmarek" nation="POL" license="100115700354" athleteid="3654">
              <RESULTS>
                <RESULT eventid="1075" points="821" reactiontime="+76" swimtime="00:02:24.29" resultid="3655" heatid="7953" lane="7" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.05" />
                    <SPLIT distance="100" swimtime="00:01:09.66" />
                    <SPLIT distance="150" swimtime="00:01:51.20" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1165" points="795" reactiontime="+85" swimtime="00:18:29.55" resultid="3656" heatid="8143" lane="4" entrytime="00:17:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.73" />
                    <SPLIT distance="100" swimtime="00:01:07.50" />
                    <SPLIT distance="150" swimtime="00:01:44.33" />
                    <SPLIT distance="200" swimtime="00:02:20.82" />
                    <SPLIT distance="250" swimtime="00:02:57.36" />
                    <SPLIT distance="300" swimtime="00:03:34.16" />
                    <SPLIT distance="350" swimtime="00:04:10.99" />
                    <SPLIT distance="400" swimtime="00:04:48.08" />
                    <SPLIT distance="450" swimtime="00:05:24.96" />
                    <SPLIT distance="500" swimtime="00:06:02.11" />
                    <SPLIT distance="550" swimtime="00:06:39.41" />
                    <SPLIT distance="600" swimtime="00:07:16.37" />
                    <SPLIT distance="650" swimtime="00:07:53.39" />
                    <SPLIT distance="700" swimtime="00:08:30.52" />
                    <SPLIT distance="750" swimtime="00:09:07.93" />
                    <SPLIT distance="800" swimtime="00:09:45.38" />
                    <SPLIT distance="850" swimtime="00:10:22.85" />
                    <SPLIT distance="900" swimtime="00:11:00.20" />
                    <SPLIT distance="950" swimtime="00:11:37.82" />
                    <SPLIT distance="1000" swimtime="00:12:15.81" />
                    <SPLIT distance="1050" swimtime="00:12:53.22" />
                    <SPLIT distance="1100" swimtime="00:13:30.93" />
                    <SPLIT distance="1150" swimtime="00:14:08.52" />
                    <SPLIT distance="1200" swimtime="00:14:46.26" />
                    <SPLIT distance="1250" swimtime="00:15:24.02" />
                    <SPLIT distance="1300" swimtime="00:16:01.77" />
                    <SPLIT distance="1350" swimtime="00:16:39.48" />
                    <SPLIT distance="1400" swimtime="00:17:16.97" />
                    <SPLIT distance="1450" swimtime="00:17:54.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="736" reactiontime="+81" swimtime="00:02:29.05" resultid="3657" heatid="8017" lane="6" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                    <SPLIT distance="100" swimtime="00:01:08.80" />
                    <SPLIT distance="150" swimtime="00:01:48.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="652" reactiontime="+81" swimtime="00:02:33.96" resultid="3658" heatid="8027" lane="4" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                    <SPLIT distance="100" swimtime="00:01:16.87" />
                    <SPLIT distance="150" swimtime="00:01:56.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="798" reactiontime="+78" swimtime="00:04:36.53" resultid="3659" heatid="8151" lane="5" entrytime="00:04:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.80" />
                    <SPLIT distance="100" swimtime="00:01:05.44" />
                    <SPLIT distance="150" swimtime="00:01:40.66" />
                    <SPLIT distance="200" swimtime="00:02:16.56" />
                    <SPLIT distance="250" swimtime="00:02:52.28" />
                    <SPLIT distance="300" swimtime="00:03:27.73" />
                    <SPLIT distance="350" swimtime="00:04:02.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="745" reactiontime="+77" swimtime="00:01:04.21" resultid="3660" heatid="8086" lane="8" entrytime="00:01:04.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="711" reactiontime="+79" swimtime="00:02:09.60" resultid="3661" heatid="8102" lane="3" entrytime="00:02:08.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.57" />
                    <SPLIT distance="100" swimtime="00:01:02.77" />
                    <SPLIT distance="150" swimtime="00:01:36.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="766" reactiontime="+81" swimtime="00:05:19.01" resultid="3662" heatid="8162" lane="3" entrytime="00:05:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                    <SPLIT distance="100" swimtime="00:01:08.35" />
                    <SPLIT distance="150" swimtime="00:01:54.14" />
                    <SPLIT distance="200" swimtime="00:02:38.00" />
                    <SPLIT distance="250" swimtime="00:03:23.19" />
                    <SPLIT distance="300" swimtime="00:04:09.30" />
                    <SPLIT distance="350" swimtime="00:04:46.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-19" firstname="Przemysław" gender="M" lastname="Waraczewski" nation="POL" license="1001155700344" athleteid="3679">
              <RESULTS>
                <RESULT eventid="1075" points="500" reactiontime="+80" swimtime="00:03:01.66" resultid="3680" heatid="7950" lane="0" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.06" />
                    <SPLIT distance="100" swimtime="00:01:29.91" />
                    <SPLIT distance="150" swimtime="00:02:20.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="586" reactiontime="+79" swimtime="00:00:38.45" resultid="3681" heatid="8004" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="1402" points="582" reactiontime="+81" swimtime="00:03:11.68" resultid="3682" heatid="8075" lane="0" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.91" />
                    <SPLIT distance="100" swimtime="00:01:32.43" />
                    <SPLIT distance="150" swimtime="00:02:21.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="579" reactiontime="+80" swimtime="00:01:26.94" resultid="3683" heatid="8129" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-27" firstname="Dariusz" gender="M" lastname="Janyga" nation="POL" license="100115700346" athleteid="3715">
              <RESULTS>
                <RESULT eventid="1165" points="537" reactiontime="+88" swimtime="00:21:08.55" resultid="3716" heatid="8143" lane="9" entrytime="00:21:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                    <SPLIT distance="100" swimtime="00:01:19.65" />
                    <SPLIT distance="150" swimtime="00:02:01.56" />
                    <SPLIT distance="200" swimtime="00:02:44.87" />
                    <SPLIT distance="250" swimtime="00:03:27.36" />
                    <SPLIT distance="300" swimtime="00:04:10.79" />
                    <SPLIT distance="350" swimtime="00:04:53.34" />
                    <SPLIT distance="400" swimtime="00:05:36.19" />
                    <SPLIT distance="450" swimtime="00:06:18.91" />
                    <SPLIT distance="500" swimtime="00:07:02.21" />
                    <SPLIT distance="550" swimtime="00:07:44.79" />
                    <SPLIT distance="600" swimtime="00:08:27.51" />
                    <SPLIT distance="650" swimtime="00:09:09.43" />
                    <SPLIT distance="700" swimtime="00:09:51.97" />
                    <SPLIT distance="750" swimtime="00:10:34.73" />
                    <SPLIT distance="800" swimtime="00:11:17.41" />
                    <SPLIT distance="850" swimtime="00:12:00.24" />
                    <SPLIT distance="900" swimtime="00:12:42.99" />
                    <SPLIT distance="950" swimtime="00:13:25.74" />
                    <SPLIT distance="1000" swimtime="00:14:08.75" />
                    <SPLIT distance="1050" swimtime="00:14:51.74" />
                    <SPLIT distance="1100" swimtime="00:15:34.65" />
                    <SPLIT distance="1150" swimtime="00:16:17.74" />
                    <SPLIT distance="1200" swimtime="00:17:01.03" />
                    <SPLIT distance="1250" swimtime="00:17:44.00" />
                    <SPLIT distance="1300" swimtime="00:18:26.13" />
                    <SPLIT distance="1350" swimtime="00:19:08.36" />
                    <SPLIT distance="1400" swimtime="00:19:50.63" />
                    <SPLIT distance="1450" swimtime="00:20:31.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="652" reactiontime="+79" swimtime="00:02:43.26" resultid="3717" heatid="8026" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.96" />
                    <SPLIT distance="100" swimtime="00:01:20.83" />
                    <SPLIT distance="150" swimtime="00:02:03.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="637" reactiontime="+81" swimtime="00:01:14.24" resultid="3718" heatid="8041" lane="0" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="532" reactiontime="+94" swimtime="00:05:16.05" resultid="3719" heatid="8152" lane="2" entrytime="00:05:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                    <SPLIT distance="100" swimtime="00:01:15.07" />
                    <SPLIT distance="150" swimtime="00:01:55.35" />
                    <SPLIT distance="200" swimtime="00:02:36.08" />
                    <SPLIT distance="250" swimtime="00:03:16.39" />
                    <SPLIT distance="300" swimtime="00:03:57.23" />
                    <SPLIT distance="350" swimtime="00:04:37.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="656" reactiontime="+80" swimtime="00:00:33.64" resultid="3720" heatid="8114" lane="9" entrytime="00:00:34.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="3722" heatid="8030" lane="7" entrytime="00:04:50.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3679" number="1" />
                    <RELAYPOSITION athleteid="3684" number="2" />
                    <RELAYPOSITION athleteid="3715" number="3" />
                    <RELAYPOSITION athleteid="3697" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1614" reactiontime="+105" swimtime="00:02:19.87" resultid="3721" heatid="8134" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.64" />
                    <SPLIT distance="100" swimtime="00:01:21.73" />
                    <SPLIT distance="150" swimtime="00:01:51.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3690" number="1" reactiontime="+105" />
                    <RELAYPOSITION athleteid="3654" number="2" />
                    <RELAYPOSITION athleteid="3675" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="3663" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="03315" nation="POL" region="PO" clubid="3760" name="KU AZS UAM Poznań">
          <CONTACT city="Poznań" email="kukowalazs@gmail.com" name="Kowalik" phone="603965223" state="WLKP" street="Zagajnikowa 9" zip="61-602" />
          <ATHLETES>
            <ATHLETE birthdate="1991-01-05" firstname="Piotr" gender="M" lastname="Kowalik" nation="POL" license="103315700017" athleteid="3769">
              <RESULTS>
                <RESULT eventid="1105" points="1032" reactiontime="+62" swimtime="00:00:24.98" resultid="3770" heatid="7972" lane="4" entrytime="00:00:24.72" />
                <RESULT eventid="1228" points="682" reactiontime="+66" swimtime="00:00:33.16" resultid="3771" heatid="8006" lane="7" entrytime="00:00:37.50" />
                <RESULT eventid="1372" points="814" reactiontime="+69" swimtime="00:00:24.66" resultid="3772" heatid="8065" lane="6" entrytime="00:00:24.44" />
                <RESULT eventid="1539" points="848" reactiontime="+50" swimtime="00:00:28.78" resultid="3773" heatid="8117" lane="5" entrytime="00:00:28.57" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-04-18" firstname="Karolina" gender="F" lastname="Stadnik" nation="POL" license="103315100003" athleteid="3761">
              <RESULTS>
                <RESULT eventid="1090" points="811" reactiontime="+76" swimtime="00:00:30.34" resultid="3762" heatid="7958" lane="4" entrytime="00:00:36.00" />
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1181" points="924" reactiontime="+77" swimtime="00:01:00.31" resultid="3763" heatid="7979" lane="6" entrytime="00:01:01.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="668" reactiontime="+73" swimtime="00:00:37.34" resultid="3764" heatid="7999" lane="5" entrytime="00:00:37.00" />
                <RESULT comment="Rekord Polski Masters" eventid="1326" points="821" reactiontime="+73" swimtime="00:01:12.39" resultid="3765" heatid="8035" lane="6" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1357" points="941" reactiontime="+74" swimtime="00:00:27.60" resultid="3766" heatid="8050" lane="4" entrytime="00:00:27.43" />
                <RESULT comment="Rekord Polski Masters" eventid="1493" points="845" reactiontime="+82" swimtime="00:02:16.36" resultid="3767" heatid="8092" lane="3" entrytime="00:02:19.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.83" />
                    <SPLIT distance="100" swimtime="00:01:05.54" />
                    <SPLIT distance="150" swimtime="00:01:41.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="898" reactiontime="+70" swimtime="00:00:32.23" resultid="3768" heatid="8107" lane="2" entrytime="00:00:33.07" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="CYP" clubid="3778" name="Limassol Nautical Club">
          <CONTACT name="Larrys Fylactou" />
          <ATHLETES>
            <ATHLETE birthdate="1964-01-29" firstname="Larrys" gender="M" lastname="Fylactou" nation="CYP" athleteid="3779">
              <RESULTS>
                <RESULT eventid="1075" points="700" reactiontime="+76" swimtime="00:02:42.41" resultid="3780" heatid="7952" lane="8" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                    <SPLIT distance="100" swimtime="00:01:17.23" />
                    <SPLIT distance="150" swimtime="00:02:06.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="689" reactiontime="+79" swimtime="00:00:31.45" resultid="3781" heatid="7968" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="1198" points="853" reactiontime="+71" swimtime="00:01:00.81" resultid="3782" heatid="7989" lane="5" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="608" swimtime="00:00:37.98" resultid="3783" heatid="8007" lane="9" entrytime="00:00:37.00" />
                <RESULT eventid="1342" points="593" reactiontime="+81" swimtime="00:01:18.35" resultid="3784" heatid="8040" lane="8" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="794" reactiontime="+75" swimtime="00:00:27.43" resultid="3785" heatid="8063" lane="9" entrytime="00:00:27.00" />
                <RESULT eventid="1539" points="710" reactiontime="+70" swimtime="00:00:34.20" resultid="3786" heatid="8114" lane="8" entrytime="00:00:34.00" />
                <RESULT eventid="1569" points="597" reactiontime="+80" swimtime="00:01:26.05" resultid="3787" heatid="8128" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="ZAC" clubid="3799" name="Marlin Gryfino">
          <CONTACT city="Gryfino" email="u210@wp.pl" name="Rosiak  Paweł" phone="512129733" state="ZACH" street="Iwaszkiewicza" zip="74-101" />
          <ATHLETES>
            <ATHLETE birthdate="1963-04-08" firstname="Dariusz" gender="M" lastname="Bauer" nation="POL" athleteid="3808">
              <RESULTS>
                <RESULT eventid="1165" points="230" reactiontime="+121" swimtime="00:29:35.26" resultid="3809" heatid="8145" lane="2" entrytime="00:28:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.20" />
                    <SPLIT distance="100" swimtime="00:01:43.52" />
                    <SPLIT distance="200" swimtime="00:03:38.74" />
                    <SPLIT distance="300" swimtime="00:05:38.14" />
                    <SPLIT distance="350" swimtime="00:06:37.40" />
                    <SPLIT distance="400" swimtime="00:07:37.35" />
                    <SPLIT distance="450" swimtime="00:08:36.37" />
                    <SPLIT distance="500" swimtime="00:09:36.36" />
                    <SPLIT distance="550" swimtime="00:12:34.52" />
                    <SPLIT distance="600" swimtime="00:11:34.14" />
                    <SPLIT distance="700" swimtime="00:15:33.15" />
                    <SPLIT distance="800" swimtime="00:17:32.11" />
                    <SPLIT distance="850" swimtime="00:18:32.37" />
                    <SPLIT distance="900" swimtime="00:19:32.50" />
                    <SPLIT distance="950" swimtime="00:20:32.91" />
                    <SPLIT distance="1000" swimtime="00:21:33.05" />
                    <SPLIT distance="1100" swimtime="00:23:33.67" />
                    <SPLIT distance="1200" swimtime="00:25:34.52" />
                    <SPLIT distance="1300" swimtime="00:27:35.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="244" reactiontime="+109" swimtime="00:01:32.30" resultid="3810" heatid="7983" lane="7" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="305" swimtime="00:00:47.77" resultid="3811" heatid="8002" lane="9" entrytime="00:00:48.00" />
                <RESULT eventid="1372" points="273" reactiontime="+102" swimtime="00:00:39.14" resultid="3812" heatid="8054" lane="3" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-16" firstname="Paweł" gender="M" lastname="Rosiak" nation="POL" athleteid="3800">
              <RESULTS>
                <RESULT comment="O4 - Start wykonany przed sygnałem (przedwczesny start)" eventid="1105" reactiontime="+71" status="DSQ" swimtime="00:00:41.80" resultid="3801" heatid="7963" lane="4" entrytime="00:00:41.00" />
                <RESULT eventid="1198" points="307" reactiontime="+87" swimtime="00:01:20.46" resultid="3802" heatid="7984" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="346" reactiontime="+83" swimtime="00:00:43.42" resultid="3803" heatid="8003" lane="4" entrytime="00:00:42.00" />
                <RESULT eventid="1372" points="412" reactiontime="+79" swimtime="00:00:33.02" resultid="3804" heatid="8056" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="1402" points="319" reactiontime="+99" swimtime="00:03:40.69" resultid="3805" heatid="8073" lane="7" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.36" />
                    <SPLIT distance="100" swimtime="00:01:47.53" />
                    <SPLIT distance="150" swimtime="00:02:46.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" status="DNS" swimtime="00:00:00.00" resultid="3806" heatid="8111" lane="7" entrytime="00:00:42.00" />
                <RESULT eventid="1569" status="DNS" swimtime="00:00:00.00" resultid="3807" heatid="8127" lane="5" entrytime="00:01:34.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5744" name="Masters Białystok">
          <CONTACT email="mbzgloszenia@gmail.pl" name="DOMINIKA MICHALIK" />
          <ATHLETES>
            <ATHLETE birthdate="1959-01-01" firstname="Joanna" gender="F" lastname="Wasilewicz" nation="POL" athleteid="5752">
              <RESULTS>
                <RESULT eventid="1090" points="416" reactiontime="+75" swimtime="00:00:46.39" resultid="5753" heatid="7956" lane="8" entrytime="00:00:47.00" />
                <RESULT eventid="1181" points="458" reactiontime="+93" swimtime="00:01:29.65" resultid="5754" heatid="7975" lane="1" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="526" reactiontime="+92" swimtime="00:00:38.25" resultid="5755" heatid="8046" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="1493" points="470" reactiontime="+81" swimtime="00:03:21.60" resultid="5756" heatid="8089" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.83" />
                    <SPLIT distance="100" swimtime="00:01:32.66" />
                    <SPLIT distance="150" swimtime="00:02:26.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-01-01" firstname="Andrzej" gender="M" lastname="Twarowski" nation="POL" athleteid="5745">
              <RESULTS>
                <RESULT eventid="1228" points="360" reactiontime="+86" swimtime="00:00:45.23" resultid="5746" heatid="8004" lane="8" entrytime="00:00:41.00" />
                <RESULT eventid="1288" points="465" reactiontime="+72" swimtime="00:03:11.75" resultid="5747" heatid="8024" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.23" />
                    <SPLIT distance="100" swimtime="00:01:33.20" />
                    <SPLIT distance="150" swimtime="00:02:23.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="427" reactiontime="+78" swimtime="00:01:27.45" resultid="5748" heatid="8039" lane="3" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="254" reactiontime="+99" swimtime="00:01:40.52" resultid="5749" heatid="8082" lane="4" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="487" reactiontime="+77" swimtime="00:00:38.79" resultid="5750" heatid="8112" lane="4" entrytime="00:00:37.00" />
                <RESULT eventid="1599" points="390" reactiontime="+95" swimtime="00:07:16.10" resultid="5751" heatid="8165" lane="2" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.42" />
                    <SPLIT distance="100" swimtime="00:01:44.97" />
                    <SPLIT distance="150" swimtime="00:02:41.23" />
                    <SPLIT distance="200" swimtime="00:03:36.06" />
                    <SPLIT distance="250" swimtime="00:04:34.45" />
                    <SPLIT distance="300" swimtime="00:05:33.69" />
                    <SPLIT distance="350" swimtime="00:06:26.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Mirosław" gender="M" lastname="Matusik" nation="POL" athleteid="5763">
              <RESULTS>
                <RESULT eventid="1105" points="502" reactiontime="+97" swimtime="00:00:35.89" resultid="5764" heatid="7965" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1198" points="507" reactiontime="+93" swimtime="00:01:16.19" resultid="5765" heatid="7985" lane="8" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="494" reactiontime="+91" swimtime="00:00:33.64" resultid="5766" heatid="8055" lane="7" entrytime="00:00:33.00" />
                <RESULT eventid="1462" status="DNS" swimtime="00:00:00.00" resultid="5767" heatid="8083" lane="1" entrytime="00:01:30.00" />
                <RESULT eventid="1509" points="495" reactiontime="+99" swimtime="00:02:52.02" resultid="5768" heatid="8097" lane="0" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                    <SPLIT distance="100" swimtime="00:01:24.39" />
                    <SPLIT distance="150" swimtime="00:02:10.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-01" firstname="Dominika" gender="F" lastname="Michalik" nation="POL" athleteid="5757">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1150" points="786" reactiontime="+82" swimtime="00:20:26.29" resultid="5758" heatid="8142" lane="4" entrytime="00:20:29.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                    <SPLIT distance="100" swimtime="00:01:13.05" />
                    <SPLIT distance="150" swimtime="00:01:52.72" />
                    <SPLIT distance="200" swimtime="00:02:33.03" />
                    <SPLIT distance="250" swimtime="00:03:13.97" />
                    <SPLIT distance="300" swimtime="00:03:54.91" />
                    <SPLIT distance="350" swimtime="00:04:36.00" />
                    <SPLIT distance="400" swimtime="00:05:17.19" />
                    <SPLIT distance="450" swimtime="00:05:58.59" />
                    <SPLIT distance="500" swimtime="00:06:39.73" />
                    <SPLIT distance="550" swimtime="00:07:20.25" />
                    <SPLIT distance="600" swimtime="00:08:01.93" />
                    <SPLIT distance="650" swimtime="00:08:43.19" />
                    <SPLIT distance="700" swimtime="00:09:24.69" />
                    <SPLIT distance="750" swimtime="00:10:04.69" />
                    <SPLIT distance="800" swimtime="00:10:44.56" />
                    <SPLIT distance="850" swimtime="00:11:26.35" />
                    <SPLIT distance="900" swimtime="00:12:07.88" />
                    <SPLIT distance="950" swimtime="00:12:50.31" />
                    <SPLIT distance="1000" swimtime="00:13:32.72" />
                    <SPLIT distance="1050" swimtime="00:14:14.32" />
                    <SPLIT distance="1100" swimtime="00:14:56.97" />
                    <SPLIT distance="1150" swimtime="00:15:39.05" />
                    <SPLIT distance="1200" swimtime="00:16:20.88" />
                    <SPLIT distance="1250" swimtime="00:17:03.22" />
                    <SPLIT distance="1300" swimtime="00:17:45.46" />
                    <SPLIT distance="1350" swimtime="00:18:26.74" />
                    <SPLIT distance="1400" swimtime="00:19:08.23" />
                    <SPLIT distance="1450" swimtime="00:19:49.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="741" swimtime="00:01:05.97" resultid="5759" heatid="7979" lane="9" entrytime="00:01:06.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="814" reactiontime="+78" swimtime="00:05:04.54" resultid="5760" heatid="8147" lane="5" entrytime="00:05:01.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.12" />
                    <SPLIT distance="100" swimtime="00:01:11.50" />
                    <SPLIT distance="150" swimtime="00:01:50.09" />
                    <SPLIT distance="200" swimtime="00:02:29.12" />
                    <SPLIT distance="250" swimtime="00:03:08.29" />
                    <SPLIT distance="300" swimtime="00:03:47.54" />
                    <SPLIT distance="350" swimtime="00:04:26.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="744" reactiontime="+80" swimtime="00:02:26.15" resultid="5761" heatid="8092" lane="7" entrytime="00:02:22.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                    <SPLIT distance="100" swimtime="00:01:09.07" />
                    <SPLIT distance="150" swimtime="00:01:47.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1584" points="706" reactiontime="+86" swimtime="00:06:01.75" resultid="5762" heatid="8159" lane="3" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.11" />
                    <SPLIT distance="100" swimtime="00:01:19.19" />
                    <SPLIT distance="150" swimtime="00:02:07.05" />
                    <SPLIT distance="200" swimtime="00:02:53.82" />
                    <SPLIT distance="250" swimtime="00:03:48.42" />
                    <SPLIT distance="300" swimtime="00:04:42.92" />
                    <SPLIT distance="350" swimtime="00:05:24.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2176" name="Masters Chełm">
          <CONTACT name="Golik Janusz" />
          <ATHLETES>
            <ATHLETE birthdate="1941-10-11" firstname="Janusz" gender="M" lastname="Golik" nation="POL" athleteid="2182">
              <RESULTS>
                <RESULT eventid="1105" points="341" reactiontime="+125" swimtime="00:00:47.89" resultid="2183" heatid="7963" lane="0" entrytime="00:00:48.00" />
                <RESULT eventid="1228" points="604" reactiontime="+103" swimtime="00:00:45.09" resultid="2184" heatid="8003" lane="9" entrytime="00:00:43.50" />
                <RESULT eventid="1258" points="186" reactiontime="+107" swimtime="00:05:22.53" resultid="2185" heatid="8014" lane="6" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.65" />
                    <SPLIT distance="100" swimtime="00:02:31.65" />
                    <SPLIT distance="150" swimtime="00:03:58.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="418" reactiontime="+111" swimtime="00:04:17.52" resultid="2186" heatid="8072" lane="1" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.46" />
                    <SPLIT distance="100" swimtime="00:02:06.62" />
                    <SPLIT distance="150" swimtime="00:03:13.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="329" reactiontime="+96" swimtime="00:01:54.97" resultid="2187" heatid="8082" lane="7" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="207" reactiontime="+110" swimtime="00:04:18.13" resultid="2188" heatid="8094" lane="0" entrytime="00:04:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.55" />
                    <SPLIT distance="100" swimtime="00:02:03.27" />
                    <SPLIT distance="150" swimtime="00:03:11.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="552" reactiontime="+98" swimtime="00:01:45.88" resultid="2189" heatid="8126" lane="2" entrytime="00:01:44.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAGOR" nation="POL" region="LBS" clubid="3839" name="Masters Gorzów">
          <CONTACT city="Klodawa Gorzowska" email="mastersgorzow@onet.eu" name="Wojciechowicz Marek" phone="602891603" state="LBS" street="Skalna 2" zip="66-415" />
          <ATHLETES>
            <ATHLETE birthdate="1974-02-20" firstname="Artur" gender="M" lastname="Rutkowski" nation="POL" license="ARUT" athleteid="3862">
              <RESULTS>
                <RESULT eventid="1075" points="484" reactiontime="+84" swimtime="00:02:48.55" resultid="3863" heatid="7951" lane="8" entrytime="00:02:48.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                    <SPLIT distance="100" swimtime="00:01:19.06" />
                    <SPLIT distance="150" swimtime="00:02:09.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="421" reactiontime="+82" swimtime="00:02:56.57" resultid="3865" heatid="8016" lane="6" entrytime="00:02:52.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                    <SPLIT distance="100" swimtime="00:01:20.40" />
                    <SPLIT distance="150" swimtime="00:02:07.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="445" reactiontime="+83" swimtime="00:06:10.66" resultid="3866" heatid="8163" lane="0" entrytime="00:06:04.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                    <SPLIT distance="100" swimtime="00:01:24.14" />
                    <SPLIT distance="150" swimtime="00:02:11.10" />
                    <SPLIT distance="200" swimtime="00:02:59.66" />
                    <SPLIT distance="250" swimtime="00:03:52.72" />
                    <SPLIT distance="300" swimtime="00:04:48.31" />
                    <SPLIT distance="350" swimtime="00:05:30.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-02-25" firstname="Tomasz" gender="M" lastname="Szymanowski" nation="POL" license="TSZYM" athleteid="3856">
              <RESULTS>
                <RESULT comment="O4 - Start wykonany przed sygnałem (przedwczesny start)" eventid="1198" status="DSQ" swimtime="00:01:03.63" resultid="3857" heatid="7989" lane="9" entrytime="00:01:04.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="533" reactiontime="+96" swimtime="00:02:44.66" resultid="3858" heatid="8026" lane="4" entrytime="00:02:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.48" />
                    <SPLIT distance="100" swimtime="00:01:18.40" />
                    <SPLIT distance="150" swimtime="00:02:01.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="580" reactiontime="+85" swimtime="00:01:14.36" resultid="3859" heatid="8041" lane="8" entrytime="00:01:16.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="513" reactiontime="+89" swimtime="00:00:29.39" resultid="3860" heatid="8060" lane="4" entrytime="00:00:28.30" entrycourse="LCM" />
                <RESULT eventid="1539" points="653" reactiontime="+76" swimtime="00:00:32.50" resultid="3861" heatid="8115" lane="6" entrytime="00:00:33.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-07-15" firstname="Marian" gender="M" lastname="Lasowy" nation="POL" license="MLAS" athleteid="3852">
              <RESULTS>
                <RESULT eventid="1165" points="372" reactiontime="+123" swimtime="00:28:28.49" resultid="3853" heatid="8145" lane="1" entrytime="00:29:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.43" />
                    <SPLIT distance="100" swimtime="00:01:41.25" />
                    <SPLIT distance="150" swimtime="00:02:36.61" />
                    <SPLIT distance="200" swimtime="00:03:32.42" />
                    <SPLIT distance="250" swimtime="00:04:29.16" />
                    <SPLIT distance="300" swimtime="00:05:25.97" />
                    <SPLIT distance="350" swimtime="00:06:22.85" />
                    <SPLIT distance="400" swimtime="00:07:20.64" />
                    <SPLIT distance="450" swimtime="00:08:17.42" />
                    <SPLIT distance="500" swimtime="00:09:14.61" />
                    <SPLIT distance="550" swimtime="00:10:12.62" />
                    <SPLIT distance="600" swimtime="00:11:09.50" />
                    <SPLIT distance="650" swimtime="00:12:07.26" />
                    <SPLIT distance="700" swimtime="00:13:05.30" />
                    <SPLIT distance="750" swimtime="00:14:03.86" />
                    <SPLIT distance="800" swimtime="00:15:02.07" />
                    <SPLIT distance="850" swimtime="00:15:59.40" />
                    <SPLIT distance="900" swimtime="00:16:57.82" />
                    <SPLIT distance="950" swimtime="00:17:55.16" />
                    <SPLIT distance="1000" swimtime="00:18:53.61" />
                    <SPLIT distance="1050" swimtime="00:19:50.85" />
                    <SPLIT distance="1100" swimtime="00:20:47.91" />
                    <SPLIT distance="1150" swimtime="00:21:46.22" />
                    <SPLIT distance="1200" swimtime="00:22:44.57" />
                    <SPLIT distance="1250" swimtime="00:23:44.56" />
                    <SPLIT distance="1300" swimtime="00:24:42.80" />
                    <SPLIT distance="1350" swimtime="00:25:40.19" />
                    <SPLIT distance="1400" swimtime="00:26:38.16" />
                    <SPLIT distance="1450" swimtime="00:27:35.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="349" reactiontime="+121" swimtime="00:03:21.16" resultid="3854" heatid="8095" lane="0" entrytime="00:03:22.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.48" />
                    <SPLIT distance="100" swimtime="00:01:36.46" />
                    <SPLIT distance="150" swimtime="00:02:29.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="343" reactiontime="+122" swimtime="00:01:53.21" resultid="3855" heatid="8126" lane="0" entrytime="00:01:52.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-05-08" firstname="Dawid" gender="M" lastname="Borus" nation="POL" license="DABOR" athleteid="3847">
              <RESULTS>
                <RESULT eventid="1288" points="647" reactiontime="+69" swimtime="00:02:43.70" resultid="3848" heatid="8028" lane="8" entrytime="00:02:28.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.46" />
                    <SPLIT distance="100" swimtime="00:01:17.59" />
                    <SPLIT distance="150" swimtime="00:02:00.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="666" reactiontime="+69" swimtime="00:01:13.16" resultid="3849" heatid="8041" lane="4" entrytime="00:01:12.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" status="DNS" swimtime="00:00:00.00" resultid="3850" heatid="8060" lane="2" entrytime="00:00:28.50" entrycourse="LCM" />
                <RESULT eventid="1539" status="DNS" swimtime="00:00:00.00" resultid="3851" heatid="8115" lane="8" entrytime="00:00:33.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-12-12" firstname="Marek" gender="M" lastname="Wojciechowicz" nation="POL" license="MWOJ" athleteid="3840">
              <RESULTS>
                <RESULT eventid="1075" points="630" reactiontime="+90" swimtime="00:02:50.08" resultid="3841" heatid="7951" lane="0" entrytime="00:02:48.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                    <SPLIT distance="100" swimtime="00:01:18.45" />
                    <SPLIT distance="150" swimtime="00:02:09.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="492" reactiontime="+106" swimtime="00:21:46.20" resultid="3842" heatid="8144" lane="7" entrytime="00:23:03.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                    <SPLIT distance="100" swimtime="00:01:19.47" />
                    <SPLIT distance="150" swimtime="00:02:03.77" />
                    <SPLIT distance="200" swimtime="00:02:48.26" />
                    <SPLIT distance="250" swimtime="00:03:32.62" />
                    <SPLIT distance="300" swimtime="00:04:17.30" />
                    <SPLIT distance="350" swimtime="00:05:01.12" />
                    <SPLIT distance="400" swimtime="00:05:45.19" />
                    <SPLIT distance="450" swimtime="00:06:28.90" />
                    <SPLIT distance="500" swimtime="00:07:13.19" />
                    <SPLIT distance="550" swimtime="00:07:57.09" />
                    <SPLIT distance="600" swimtime="00:08:41.49" />
                    <SPLIT distance="650" swimtime="00:09:25.53" />
                    <SPLIT distance="700" swimtime="00:10:09.96" />
                    <SPLIT distance="750" swimtime="00:10:54.01" />
                    <SPLIT distance="800" swimtime="00:11:38.51" />
                    <SPLIT distance="850" swimtime="00:12:21.65" />
                    <SPLIT distance="900" swimtime="00:13:05.58" />
                    <SPLIT distance="950" swimtime="00:13:49.01" />
                    <SPLIT distance="1000" swimtime="00:14:32.73" />
                    <SPLIT distance="1050" swimtime="00:15:15.94" />
                    <SPLIT distance="1100" swimtime="00:15:59.93" />
                    <SPLIT distance="1150" swimtime="00:16:43.33" />
                    <SPLIT distance="1200" swimtime="00:17:27.39" />
                    <SPLIT distance="1250" swimtime="00:18:11.18" />
                    <SPLIT distance="1300" swimtime="00:18:55.70" />
                    <SPLIT distance="1350" swimtime="00:19:39.28" />
                    <SPLIT distance="1400" swimtime="00:20:23.54" />
                    <SPLIT distance="1450" swimtime="00:21:06.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="649" reactiontime="+85" swimtime="00:01:04.49" resultid="3843" heatid="7989" lane="1" entrytime="00:01:04.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="655" reactiontime="+81" swimtime="00:00:28.97" resultid="3844" heatid="8060" lane="3" entrytime="00:00:28.50" entrycourse="LCM" />
                <RESULT eventid="1432" points="482" reactiontime="+83" swimtime="00:05:26.64" resultid="3845" heatid="8152" lane="8" entrytime="00:05:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                    <SPLIT distance="100" swimtime="00:01:12.53" />
                    <SPLIT distance="150" swimtime="00:01:54.08" />
                    <SPLIT distance="200" swimtime="00:02:36.59" />
                    <SPLIT distance="250" swimtime="00:03:19.35" />
                    <SPLIT distance="300" swimtime="00:04:02.49" />
                    <SPLIT distance="350" swimtime="00:04:44.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="520" reactiontime="+97" swimtime="00:02:28.37" resultid="3846" heatid="8100" lane="7" entrytime="00:02:23.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.99" />
                    <SPLIT distance="100" swimtime="00:01:10.30" />
                    <SPLIT distance="150" swimtime="00:01:49.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1318" reactiontime="+95" swimtime="00:04:30.46" resultid="3867" heatid="8030" lane="3" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                    <SPLIT distance="100" swimtime="00:01:04.82" />
                    <SPLIT distance="150" swimtime="00:01:35.82" />
                    <SPLIT distance="200" swimtime="00:02:11.56" />
                    <SPLIT distance="250" swimtime="00:02:42.61" />
                    <SPLIT distance="300" swimtime="00:03:16.79" />
                    <SPLIT distance="350" swimtime="00:03:51.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3847" number="1" reactiontime="+95" />
                    <RELAYPOSITION athleteid="3862" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="3856" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="3840" number="4" reactiontime="+66" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="KORONA KRA" nation="POL" region="MAL" clubid="3868" name="Masters Korona Kraków">
          <CONTACT city="Kraków" email="masterskorona@wp.pl" name="Mariola Kuliś" phone="500677133" state="MAŁ" />
          <ATHLETES>
            <ATHLETE birthdate="1981-02-26" firstname="Anna" gender="F" lastname="Kasprzykowska" nation="POL" athleteid="3885">
              <RESULTS>
                <RESULT eventid="1090" points="148" reactiontime="+94" swimtime="00:00:55.32" resultid="3886" heatid="7955" lane="5" entrytime="00:00:51.00" />
                <RESULT eventid="1243" points="129" reactiontime="+90" swimtime="00:04:50.14" resultid="3887" heatid="8011" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.33" />
                    <SPLIT distance="100" swimtime="00:02:23.09" />
                    <SPLIT distance="150" swimtime="00:03:42.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="196" reactiontime="+91" swimtime="00:00:46.70" resultid="3888" heatid="8045" lane="8" entrytime="00:00:45.00" />
                <RESULT eventid="1493" points="156" reactiontime="+85" swimtime="00:03:57.04" resultid="3889" heatid="8087" lane="4" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.68" />
                    <SPLIT distance="100" swimtime="00:01:54.89" />
                    <SPLIT distance="150" swimtime="00:02:56.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-26" firstname="Marta" gender="F" lastname="Wysocka" nation="POL" athleteid="3934">
              <RESULTS>
                <RESULT eventid="1213" points="734" swimtime="00:00:42.50" resultid="3935" heatid="7998" lane="6" entrytime="00:00:41.00" />
                <RESULT eventid="1387" points="905" reactiontime="+93" swimtime="00:03:18.49" resultid="3936" heatid="8070" lane="8" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.64" />
                    <SPLIT distance="100" swimtime="00:01:35.71" />
                    <SPLIT distance="150" swimtime="00:02:26.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="782" reactiontime="+87" swimtime="00:01:32.69" resultid="3937" heatid="8122" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-05-06" firstname="Matteo" gender="M" lastname="Morlupi" nation="POL" athleteid="3916">
              <RESULTS>
                <RESULT eventid="1198" points="312" reactiontime="+83" swimtime="00:01:16.63" resultid="3917" heatid="7985" lane="9" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="396" reactiontime="+98" swimtime="00:00:39.75" resultid="3918" heatid="8006" lane="8" entrytime="00:00:38.00" />
                <RESULT eventid="1372" points="394" reactiontime="+92" swimtime="00:00:32.09" resultid="3919" heatid="8056" lane="1" entrytime="00:00:32.00" />
                <RESULT eventid="1402" points="353" reactiontime="+96" swimtime="00:03:34.11" resultid="3920" heatid="8074" lane="5" entrytime="00:03:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.14" />
                    <SPLIT distance="100" swimtime="00:01:40.01" />
                    <SPLIT distance="150" swimtime="00:02:38.32" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K15 - Brak dotknięcia ściany obydwoma rozłączonymi dłońmi przy nawrocie lub na zakończenie wyścigu" eventid="1569" reactiontime="+87" status="DSQ" swimtime="00:01:31.88" resultid="3921" heatid="8129" lane="0" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-10-22" firstname="Maria" gender="F" lastname="Mleczko" nation="POL" athleteid="3907">
              <RESULTS>
                <RESULT eventid="1058" points="157" reactiontime="+125" swimtime="00:05:43.13" resultid="3908" heatid="7941" lane="3" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.37" />
                    <SPLIT distance="100" swimtime="00:02:58.80" />
                    <SPLIT distance="150" swimtime="00:04:29.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="100" reactiontime="+110" swimtime="00:01:17.01" resultid="3909" heatid="7955" lane="0" entrytime="00:01:16.00" />
                <RESULT eventid="1181" points="148" reactiontime="+102" swimtime="00:02:15.84" resultid="3910" heatid="7973" lane="5" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="266" reactiontime="+112" swimtime="00:01:04.56" resultid="3911" heatid="7995" lane="0" entrytime="00:01:05.00" />
                <RESULT eventid="1387" points="229" reactiontime="+107" swimtime="00:05:37.93" resultid="3912" heatid="8067" lane="9" entrytime="00:05:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.41" />
                    <SPLIT distance="100" swimtime="00:02:44.55" />
                    <SPLIT distance="150" swimtime="00:04:16.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="91" reactiontime="+103" swimtime="00:03:12.00" resultid="3913" heatid="8078" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:25.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="171" reactiontime="+108" swimtime="00:04:51.89" resultid="3914" heatid="8087" lane="6" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.98" />
                    <SPLIT distance="100" swimtime="00:02:21.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="270" reactiontime="+106" swimtime="00:02:27.51" resultid="3915" heatid="8119" lane="1" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-08-26" firstname="Andrzej" gender="M" lastname="Mleczko" nation="POL" athleteid="3898">
              <RESULTS>
                <RESULT eventid="1075" points="400" reactiontime="+138" swimtime="00:03:44.76" resultid="3899" heatid="7947" lane="0" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.51" />
                    <SPLIT distance="100" swimtime="00:01:49.96" />
                    <SPLIT distance="150" swimtime="00:02:57.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="430" reactiontime="+122" swimtime="00:14:28.84" resultid="3900" heatid="8140" lane="8" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.08" />
                    <SPLIT distance="100" swimtime="00:01:40.86" />
                    <SPLIT distance="150" swimtime="00:02:36.57" />
                    <SPLIT distance="200" swimtime="00:03:32.90" />
                    <SPLIT distance="250" swimtime="00:04:28.86" />
                    <SPLIT distance="300" swimtime="00:05:24.96" />
                    <SPLIT distance="350" swimtime="00:06:20.41" />
                    <SPLIT distance="400" swimtime="00:07:15.50" />
                    <SPLIT distance="450" swimtime="00:08:10.46" />
                    <SPLIT distance="500" swimtime="00:09:05.23" />
                    <SPLIT distance="550" swimtime="00:10:00.06" />
                    <SPLIT distance="600" swimtime="00:10:55.25" />
                    <SPLIT distance="650" swimtime="00:11:50.37" />
                    <SPLIT distance="700" swimtime="00:12:45.80" />
                    <SPLIT distance="750" swimtime="00:13:40.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="678" reactiontime="+113" swimtime="00:01:15.11" resultid="3901" heatid="7984" lane="3" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="245" reactiontime="+128" swimtime="00:04:41.11" resultid="3902" heatid="8014" lane="5" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.32" />
                    <SPLIT distance="100" swimtime="00:02:08.34" />
                    <SPLIT distance="150" swimtime="00:03:20.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="616" reactiontime="+129" swimtime="00:00:33.83" resultid="3903" heatid="8055" lane="0" entrytime="00:00:34.00" />
                <RESULT eventid="1432" points="451" reactiontime="+123" swimtime="00:06:58.96" resultid="3904" heatid="8155" lane="6" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.40" />
                    <SPLIT distance="100" swimtime="00:01:43.21" />
                    <SPLIT distance="150" swimtime="00:02:39.23" />
                    <SPLIT distance="200" swimtime="00:03:32.99" />
                    <SPLIT distance="250" swimtime="00:04:26.73" />
                    <SPLIT distance="300" swimtime="00:05:19.92" />
                    <SPLIT distance="350" swimtime="00:06:11.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="538" reactiontime="+129" swimtime="00:03:04.96" resultid="3905" heatid="8096" lane="2" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.27" />
                    <SPLIT distance="100" swimtime="00:01:26.48" />
                    <SPLIT distance="150" swimtime="00:02:15.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="337" reactiontime="+124" swimtime="00:09:01.86" resultid="3906" heatid="8167" lane="3" entrytime="00:08:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.17" />
                    <SPLIT distance="100" swimtime="00:02:08.25" />
                    <SPLIT distance="150" swimtime="00:03:19.82" />
                    <SPLIT distance="200" swimtime="00:04:32.40" />
                    <SPLIT distance="250" swimtime="00:05:47.23" />
                    <SPLIT distance="300" swimtime="00:07:02.11" />
                    <SPLIT distance="350" swimtime="00:08:04.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-12-07" firstname="Robert" gender="M" lastname="Kominiak" nation="POL" athleteid="3938">
              <RESULTS>
                <RESULT eventid="1075" points="570" reactiontime="+85" swimtime="00:02:53.91" resultid="3939" heatid="7951" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.89" />
                    <SPLIT distance="100" swimtime="00:01:21.09" />
                    <SPLIT distance="150" swimtime="00:02:09.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="635" reactiontime="+70" swimtime="00:00:32.32" resultid="3940" heatid="7969" lane="9" entrytime="00:00:31.00" />
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1228" points="823" reactiontime="+77" swimtime="00:00:34.33" resultid="3941" heatid="8009" lane="4" entrytime="00:00:33.00" />
                <RESULT comment="K16 - Niejednoczesne dotknięcie ściany dłońmi przy nawrocie lub na zakończenie wyścigu" eventid="1402" reactiontime="+77" status="DSQ" swimtime="00:03:09.19" resultid="3942" heatid="8076" lane="3" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.31" />
                    <SPLIT distance="100" swimtime="00:01:28.82" />
                    <SPLIT distance="150" swimtime="00:02:18.48" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1569" points="778" reactiontime="+74" swimtime="00:01:18.80" resultid="3943" heatid="8131" lane="1" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-05-16" firstname="Tadeusz" gender="M" lastname="Krawczyk" nation="POL" athleteid="3890">
              <RESULTS>
                <RESULT eventid="1075" points="140" reactiontime="+121" swimtime="00:05:48.70" resultid="3891" heatid="7945" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.45" />
                    <SPLIT distance="100" swimtime="00:02:51.46" />
                    <SPLIT distance="150" swimtime="00:04:49.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="60" reactiontime="+118" swimtime="00:01:25.45" resultid="3892" heatid="7961" lane="5" />
                <RESULT eventid="1198" points="234" reactiontime="+119" swimtime="00:01:46.72" resultid="3893" heatid="7981" lane="6" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="117" reactiontime="+97" swimtime="00:02:37.92" resultid="3894" heatid="8036" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="233" reactiontime="+115" swimtime="00:00:46.22" resultid="3895" heatid="8052" lane="6" entrytime="00:00:47.00" />
                <RESULT eventid="1509" points="205" reactiontime="+117" swimtime="00:04:19.24" resultid="3896" heatid="8093" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.50" />
                    <SPLIT distance="100" swimtime="00:01:59.95" />
                    <SPLIT distance="150" swimtime="00:03:13.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="143" reactiontime="+99" swimtime="00:01:06.64" resultid="3897" heatid="8109" lane="9" entrytime="00:01:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-04-22" firstname="Alicja" gender="F" lastname="Romańska" nation="POL" athleteid="3944">
              <RESULTS>
                <RESULT eventid="1090" points="142" reactiontime="+102" swimtime="00:00:56.98" resultid="3945" heatid="7954" lane="3" />
                <RESULT eventid="1120" points="295" reactiontime="+99" swimtime="00:14:42.92" resultid="3946" heatid="8137" lane="7" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.86" />
                    <SPLIT distance="100" swimtime="00:01:45.90" />
                    <SPLIT distance="150" swimtime="00:02:42.32" />
                    <SPLIT distance="200" swimtime="00:03:39.70" />
                    <SPLIT distance="250" swimtime="00:04:35.67" />
                    <SPLIT distance="300" swimtime="00:05:31.44" />
                    <SPLIT distance="350" swimtime="00:06:27.58" />
                    <SPLIT distance="400" swimtime="00:07:23.46" />
                    <SPLIT distance="450" swimtime="00:08:18.24" />
                    <SPLIT distance="500" swimtime="00:09:13.76" />
                    <SPLIT distance="550" swimtime="00:10:09.12" />
                    <SPLIT distance="600" swimtime="00:11:04.76" />
                    <SPLIT distance="650" swimtime="00:12:00.38" />
                    <SPLIT distance="700" swimtime="00:12:55.44" />
                    <SPLIT distance="750" swimtime="00:13:49.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="203" reactiontime="+98" swimtime="00:01:43.48" resultid="3947" heatid="7974" lane="1" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="249" reactiontime="+89" swimtime="00:00:43.74" resultid="3948" heatid="8045" lane="0" entrytime="00:00:47.00" />
                <RESULT eventid="1417" points="258" reactiontime="+86" swimtime="00:07:24.16" resultid="3949" heatid="8149" lane="6" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.82" />
                    <SPLIT distance="100" swimtime="00:01:46.34" />
                    <SPLIT distance="150" swimtime="00:02:44.15" />
                    <SPLIT distance="200" swimtime="00:03:41.46" />
                    <SPLIT distance="250" swimtime="00:04:38.32" />
                    <SPLIT distance="300" swimtime="00:05:35.34" />
                    <SPLIT distance="350" swimtime="00:06:30.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-08-18" firstname="Jadwiga" gender="F" lastname="Górecka - Burkot" nation="POL" athleteid="3880">
              <RESULTS>
                <RESULT eventid="1090" points="603" reactiontime="+84" swimtime="00:00:40.99" resultid="3881" heatid="7956" lane="4" entrytime="00:00:41.00" />
                <RESULT eventid="1181" points="606" reactiontime="+82" swimtime="00:01:21.70" resultid="3882" heatid="7975" lane="5" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="686" reactiontime="+78" swimtime="00:00:35.01" resultid="3883" heatid="8046" lane="3" entrytime="00:00:36.00" />
                <RESULT eventid="1493" points="573" reactiontime="+69" swimtime="00:03:08.78" resultid="3884" heatid="8088" lane="8" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.33" />
                    <SPLIT distance="100" swimtime="00:01:31.71" />
                    <SPLIT distance="150" swimtime="00:02:21.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-07-04" firstname="Stanisław" gender="M" lastname="Waga" nation="POL" athleteid="3926">
              <RESULTS>
                <RESULT eventid="1165" points="397" reactiontime="+106" swimtime="00:32:00.62" resultid="3927" heatid="8146" lane="5" entrytime="00:43:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.10" />
                    <SPLIT distance="100" swimtime="00:01:56.28" />
                    <SPLIT distance="150" swimtime="00:03:02.00" />
                    <SPLIT distance="200" swimtime="00:04:09.26" />
                    <SPLIT distance="250" swimtime="00:05:16.85" />
                    <SPLIT distance="300" swimtime="00:06:23.03" />
                    <SPLIT distance="350" swimtime="00:07:28.53" />
                    <SPLIT distance="400" swimtime="00:08:33.64" />
                    <SPLIT distance="450" swimtime="00:09:40.12" />
                    <SPLIT distance="500" swimtime="00:10:45.18" />
                    <SPLIT distance="550" swimtime="00:11:50.68" />
                    <SPLIT distance="600" swimtime="00:12:55.29" />
                    <SPLIT distance="650" swimtime="00:14:00.32" />
                    <SPLIT distance="700" swimtime="00:15:05.09" />
                    <SPLIT distance="750" swimtime="00:16:09.38" />
                    <SPLIT distance="800" swimtime="00:17:13.26" />
                    <SPLIT distance="850" swimtime="00:18:17.63" />
                    <SPLIT distance="900" swimtime="00:19:21.70" />
                    <SPLIT distance="950" swimtime="00:20:25.98" />
                    <SPLIT distance="1000" swimtime="00:21:30.16" />
                    <SPLIT distance="1050" swimtime="00:22:32.77" />
                    <SPLIT distance="1100" swimtime="00:23:37.23" />
                    <SPLIT distance="1150" swimtime="00:24:40.86" />
                    <SPLIT distance="1200" swimtime="00:25:44.15" />
                    <SPLIT distance="1250" swimtime="00:26:46.94" />
                    <SPLIT distance="1300" swimtime="00:27:50.47" />
                    <SPLIT distance="1350" swimtime="00:28:55.40" />
                    <SPLIT distance="1400" swimtime="00:29:58.89" />
                    <SPLIT distance="1450" swimtime="00:30:59.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="349" reactiontime="+89" swimtime="00:01:43.29" resultid="3928" heatid="7981" lane="3" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="211" reactiontime="+99" swimtime="00:01:06.37" resultid="3929" heatid="8000" lane="7" entrytime="00:01:15.00" />
                <RESULT eventid="1372" points="344" reactiontime="+105" swimtime="00:00:44.87" resultid="3930" heatid="8052" lane="5" entrytime="00:00:45.00" />
                <RESULT eventid="1432" points="326" reactiontime="+97" swimtime="00:08:19.44" resultid="3931" heatid="8156" lane="2" entrytime="00:11:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.17" />
                    <SPLIT distance="100" swimtime="00:01:50.37" />
                    <SPLIT distance="150" swimtime="00:02:54.63" />
                    <SPLIT distance="200" swimtime="00:04:01.00" />
                    <SPLIT distance="250" swimtime="00:05:06.48" />
                    <SPLIT distance="300" swimtime="00:06:12.70" />
                    <SPLIT distance="350" swimtime="00:07:17.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="336" reactiontime="+105" swimtime="00:03:49.74" resultid="3932" heatid="8094" lane="3" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.34" />
                    <SPLIT distance="100" swimtime="00:01:47.76" />
                    <SPLIT distance="150" swimtime="00:02:48.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="227" reactiontime="+103" swimtime="00:02:27.38" resultid="3933" heatid="8124" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-03-26" firstname="Józef" gender="M" lastname="Śmigielski" nation="POL" athleteid="3922">
              <RESULTS>
                <RESULT eventid="1288" points="232" reactiontime="+104" swimtime="00:04:21.82" resultid="3923" heatid="8023" lane="2" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.34" />
                    <SPLIT distance="100" swimtime="00:02:05.34" />
                    <SPLIT distance="150" swimtime="00:03:13.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="168" reactiontime="+120" swimtime="00:02:13.77" resultid="3924" heatid="8037" lane="0" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="175" reactiontime="+101" swimtime="00:00:59.83" resultid="3925" heatid="8109" lane="1" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-07-27" firstname="Mariola" gender="F" lastname="Kuliś" nation="POL" athleteid="3872">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1090" points="778" reactiontime="+70" swimtime="00:00:32.94" resultid="3873" heatid="7960" lane="9" entrytime="00:00:34.00" />
                <RESULT eventid="1181" points="741" reactiontime="+78" swimtime="00:01:09.31" resultid="3874" heatid="7978" lane="8" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1213" points="971" reactiontime="+66" swimtime="00:00:36.95" resultid="3875" heatid="7999" lane="6" entrytime="00:00:38.50" />
                <RESULT eventid="1326" points="762" reactiontime="+66" swimtime="00:01:20.00" resultid="3876" heatid="8033" lane="7" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.98" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1357" points="854" reactiontime="+75" swimtime="00:00:29.88" resultid="3877" heatid="8048" lane="2" entrytime="00:00:32.00" />
                <RESULT eventid="1524" points="777" reactiontime="+62" swimtime="00:00:36.09" resultid="3878" heatid="8104" lane="2" entrytime="00:00:55.00" />
                <RESULT comment="Rekord Polski Masters" eventid="1554" points="789" reactiontime="+77" swimtime="00:01:26.70" resultid="3879" heatid="8123" lane="1" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="280" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1318" swimtime="00:07:01.39" resultid="3950" heatid="8030" lane="8" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.29" />
                    <SPLIT distance="100" swimtime="00:02:06.09" />
                    <SPLIT distance="150" swimtime="00:02:44.19" />
                    <SPLIT distance="200" swimtime="00:03:24.65" />
                    <SPLIT distance="250" swimtime="00:04:11.98" />
                    <SPLIT distance="300" swimtime="00:05:13.10" />
                    <SPLIT distance="350" swimtime="00:06:03.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3922" number="1" />
                    <RELAYPOSITION athleteid="3898" number="2" reactiontime="+73" />
                    <RELAYPOSITION athleteid="3890" number="3" reactiontime="+76" />
                    <RELAYPOSITION athleteid="3926" number="4" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1614" reactiontime="+65" swimtime="00:02:23.73" resultid="3951" heatid="8134" lane="7" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                    <SPLIT distance="100" swimtime="00:01:18.70" />
                    <SPLIT distance="150" swimtime="00:01:49.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3872" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="3934" number="2" />
                    <RELAYPOSITION athleteid="3938" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="3898" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1614" reactiontime="+89" swimtime="00:03:36.23" resultid="3952" heatid="8133" lane="7" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.01" />
                    <SPLIT distance="100" swimtime="00:02:07.58" />
                    <SPLIT distance="150" swimtime="00:02:52.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3922" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="3907" number="2" />
                    <RELAYPOSITION athleteid="3880" number="3" reactiontime="+67" />
                    <RELAYPOSITION athleteid="3926" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MASKRAS" nation="POL" region="LU" clubid="2144" name="Masters Krasnik">
          <CONTACT city="Kraśnik" email="jurek@krasnik.info" internet="www.masterskrasnik.za.pl" name="Michalczyk Jerzy" phone="601 69 89 77" state="LUB." street="Żwirki i Wigury 2" zip="23-204" />
          <ATHLETES>
            <ATHLETE birthdate="1971-03-04" firstname="Mirosław" gender="M" lastname="Leszczyński" nation="POL" athleteid="2150">
              <RESULTS>
                <RESULT eventid="1228" points="493" reactiontime="+91" swimtime="00:00:38.60" resultid="2151" heatid="8005" lane="9" entrytime="00:00:40.00" />
                <RESULT eventid="1402" points="559" reactiontime="+86" swimtime="00:03:03.06" resultid="2152" heatid="8075" lane="7" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.07" />
                    <SPLIT distance="100" swimtime="00:01:28.68" />
                    <SPLIT distance="150" swimtime="00:02:16.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="499" reactiontime="+90" swimtime="00:01:26.63" resultid="2153" heatid="8125" lane="8" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-09" firstname="Jerzy" gender="M" lastname="Michalczyk" nation="POL" athleteid="2170">
              <RESULTS>
                <RESULT eventid="1075" points="262" reactiontime="+93" swimtime="00:04:02.29" resultid="2171" heatid="7945" lane="4" entrytime="00:04:05.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.73" />
                    <SPLIT distance="100" swimtime="00:01:56.21" />
                    <SPLIT distance="150" swimtime="00:03:06.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="211" reactiontime="+96" swimtime="00:00:52.10" resultid="2172" heatid="8001" lane="1" entrytime="00:00:50.00" />
                <RESULT eventid="1258" points="150" reactiontime="+98" swimtime="00:04:51.90" resultid="2173" heatid="8014" lane="0" entrytime="00:04:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.77" />
                    <SPLIT distance="100" swimtime="00:02:12.01" />
                    <SPLIT distance="150" swimtime="00:03:32.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="268" swimtime="00:04:16.64" resultid="2174" heatid="8071" lane="6" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.57" />
                    <SPLIT distance="100" swimtime="00:02:05.42" />
                    <SPLIT distance="150" swimtime="00:03:13.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="227" reactiontime="+88" swimtime="00:01:59.25" resultid="2175" heatid="8126" lane="9" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-09-07" firstname="Andrzej" gender="M" lastname="Cis" nation="POL" athleteid="2154">
              <RESULTS>
                <RESULT eventid="1075" points="405" reactiontime="+69" swimtime="00:03:29.40" resultid="2155" heatid="7948" lane="5" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.07" />
                    <SPLIT distance="100" swimtime="00:01:40.95" />
                    <SPLIT distance="150" swimtime="00:02:44.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="402" reactiontime="+75" swimtime="00:13:49.99" resultid="2156" heatid="8140" lane="6" entrytime="00:13:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.38" />
                    <SPLIT distance="100" swimtime="00:01:33.84" />
                    <SPLIT distance="150" swimtime="00:02:25.28" />
                    <SPLIT distance="200" swimtime="00:03:18.80" />
                    <SPLIT distance="250" swimtime="00:04:11.92" />
                    <SPLIT distance="300" swimtime="00:05:06.03" />
                    <SPLIT distance="350" swimtime="00:06:00.72" />
                    <SPLIT distance="400" swimtime="00:06:55.21" />
                    <SPLIT distance="450" swimtime="00:07:49.36" />
                    <SPLIT distance="500" swimtime="00:08:42.17" />
                    <SPLIT distance="550" swimtime="00:09:35.90" />
                    <SPLIT distance="600" swimtime="00:10:28.79" />
                    <SPLIT distance="650" swimtime="00:11:22.31" />
                    <SPLIT distance="700" swimtime="00:12:13.94" />
                    <SPLIT distance="750" swimtime="00:13:05.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="565" reactiontime="+82" swimtime="00:01:13.49" resultid="2157" heatid="7986" lane="0" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="522" reactiontime="+69" swimtime="00:03:18.86" resultid="2158" heatid="8025" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.25" />
                    <SPLIT distance="100" swimtime="00:01:38.25" />
                    <SPLIT distance="150" swimtime="00:02:32.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="223" reactiontime="+90" swimtime="00:01:58.54" resultid="2159" heatid="8039" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="569" reactiontime="+66" swimtime="00:00:32.11" resultid="2160" heatid="8057" lane="0" entrytime="00:00:30.00" />
                <RESULT eventid="1539" points="547" reactiontime="+60" swimtime="00:00:39.71" resultid="2161" heatid="8112" lane="7" entrytime="00:00:38.00" />
                <RESULT eventid="1599" status="DNS" swimtime="00:00:00.00" resultid="2162" heatid="8165" lane="0" entrytime="00:07:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-11-05" firstname="Krzysztof" gender="M" lastname="Samonek" nation="POL" athleteid="2163">
              <RESULTS>
                <RESULT eventid="1075" points="296" reactiontime="+97" swimtime="00:03:52.56" resultid="2164" heatid="7946" lane="9" entrytime="00:04:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.01" />
                    <SPLIT distance="100" swimtime="00:01:51.23" />
                    <SPLIT distance="150" swimtime="00:03:00.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="176" reactiontime="+106" swimtime="00:04:36.46" resultid="2165" heatid="8014" lane="8" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.57" />
                    <SPLIT distance="100" swimtime="00:02:14.27" />
                    <SPLIT distance="150" swimtime="00:03:30.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="347" reactiontime="+86" swimtime="00:03:47.90" resultid="2166" heatid="8023" lane="5" entrytime="00:04:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.91" />
                    <SPLIT distance="100" swimtime="00:01:53.79" />
                    <SPLIT distance="150" swimtime="00:02:53.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" status="DNS" swimtime="00:00:00.00" resultid="2167" heatid="8037" lane="6" entrytime="00:01:57.00" />
                <RESULT eventid="1462" points="165" reactiontime="+93" swimtime="00:01:57.67" resultid="2168" heatid="8082" lane="1" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="281" reactiontime="+96" swimtime="00:08:27.90" resultid="2169" heatid="8166" lane="9" entrytime="00:08:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.55" />
                    <SPLIT distance="100" swimtime="00:02:04.28" />
                    <SPLIT distance="150" swimtime="00:03:09.73" />
                    <SPLIT distance="200" swimtime="00:04:10.24" />
                    <SPLIT distance="250" swimtime="00:05:23.54" />
                    <SPLIT distance="300" swimtime="00:06:35.87" />
                    <SPLIT distance="350" swimtime="00:07:33.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-02-09" firstname="Marcin" gender="M" lastname="Mazurek" nation="POL" athleteid="2145">
              <RESULTS>
                <RESULT eventid="1198" points="374" reactiontime="+85" swimtime="00:01:15.39" resultid="2146" heatid="7985" lane="0" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="429" reactiontime="+83" swimtime="00:00:32.59" resultid="2147" heatid="8059" lane="7" entrytime="00:00:29.00" />
                <RESULT eventid="1432" points="281" reactiontime="+91" swimtime="00:06:28.02" resultid="2148" heatid="8153" lane="9" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                    <SPLIT distance="100" swimtime="00:01:23.94" />
                    <SPLIT distance="150" swimtime="00:02:11.41" />
                    <SPLIT distance="200" swimtime="00:03:00.82" />
                    <SPLIT distance="250" swimtime="00:03:51.84" />
                    <SPLIT distance="300" swimtime="00:04:44.05" />
                    <SPLIT distance="350" swimtime="00:05:37.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="309" reactiontime="+86" swimtime="00:02:55.12" resultid="2149" heatid="8097" lane="6" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.92" />
                    <SPLIT distance="100" swimtime="00:01:22.37" />
                    <SPLIT distance="150" swimtime="00:02:09.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3990" name="Masters Szczecinek">
          <CONTACT name="Andrzej Wojnicz" />
          <ATHLETES>
            <ATHLETE birthdate="1933-02-19" firstname="Zbigniew" gender="M" lastname="Ludwiczak" nation="POL" athleteid="4014">
              <RESULTS>
                <RESULT eventid="1135" points="404" swimtime="00:19:04.24" resultid="4015" heatid="8141" lane="3" entrytime="00:18:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.14" />
                    <SPLIT distance="100" swimtime="00:02:10.40" />
                    <SPLIT distance="150" swimtime="00:03:20.95" />
                    <SPLIT distance="200" swimtime="00:04:32.57" />
                    <SPLIT distance="250" swimtime="00:05:43.10" />
                    <SPLIT distance="300" swimtime="00:06:54.52" />
                    <SPLIT distance="350" swimtime="00:08:06.78" />
                    <SPLIT distance="400" swimtime="00:09:18.74" />
                    <SPLIT distance="450" swimtime="00:10:31.00" />
                    <SPLIT distance="500" swimtime="00:11:44.04" />
                    <SPLIT distance="550" swimtime="00:12:57.40" />
                    <SPLIT distance="600" swimtime="00:14:12.34" />
                    <SPLIT distance="650" swimtime="00:15:26.25" />
                    <SPLIT distance="700" swimtime="00:16:41.89" />
                    <SPLIT distance="750" swimtime="00:17:55.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="374" swimtime="00:01:57.78" resultid="4016" heatid="7981" lane="7" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="362" reactiontime="+113" swimtime="00:05:13.67" resultid="4017" heatid="8023" lane="1" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.36" />
                    <SPLIT distance="100" swimtime="00:02:36.23" />
                    <SPLIT distance="150" swimtime="00:03:58.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="406" reactiontime="+122" swimtime="00:02:16.57" resultid="4018" heatid="8036" lane="5" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="422" swimtime="00:09:03.04" resultid="4019" heatid="8156" lane="6" entrytime="00:08:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.38" />
                    <SPLIT distance="100" swimtime="00:02:07.58" />
                    <SPLIT distance="150" swimtime="00:03:16.56" />
                    <SPLIT distance="200" swimtime="00:04:27.38" />
                    <SPLIT distance="250" swimtime="00:05:37.11" />
                    <SPLIT distance="300" swimtime="00:06:48.03" />
                    <SPLIT distance="350" swimtime="00:07:57.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="420" swimtime="00:04:10.40" resultid="4020" heatid="8094" lane="9" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.49" />
                    <SPLIT distance="100" swimtime="00:02:02.31" />
                    <SPLIT distance="150" swimtime="00:03:06.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="415" reactiontime="+126" swimtime="00:01:00.02" resultid="4021" heatid="8109" lane="7" entrytime="00:00:59.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-11-23" firstname="Krystyna" gender="F" lastname="Witkowska" nation="POL" athleteid="4000">
              <RESULTS>
                <RESULT eventid="1181" points="146" reactiontime="+145" swimtime="00:02:54.04" resultid="4001" heatid="7973" lane="7" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="80" reactiontime="+122" swimtime="00:01:50.40" resultid="4002" heatid="7994" lane="2" entrytime="00:01:44.00" />
                <RESULT eventid="1326" points="131" reactiontime="+111" swimtime="00:03:33.58" resultid="4003" heatid="8032" lane="2" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:40.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="127" reactiontime="+136" swimtime="00:01:19.13" resultid="4004" heatid="8044" lane="6" entrytime="00:01:20.00" />
                <RESULT eventid="1493" points="163" reactiontime="+139" swimtime="00:06:03.68" resultid="4005" heatid="8087" lane="2" entrytime="00:06:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.95" />
                    <SPLIT distance="100" swimtime="00:02:57.62" />
                    <SPLIT distance="150" swimtime="00:04:32.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="103" reactiontime="+69" swimtime="00:01:38.10" resultid="4006" heatid="8103" lane="3" entrytime="00:01:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-03-27" firstname="Ryszard" gender="M" lastname="Przelicki" nation="POL" athleteid="4022">
              <RESULTS>
                <RESULT eventid="1105" points="66" reactiontime="+121" swimtime="00:01:30.48" resultid="4023" heatid="7962" lane="1" entrytime="00:01:23.00" />
                <RESULT eventid="1228" points="150" reactiontime="+110" swimtime="00:01:14.47" resultid="4024" heatid="8000" lane="2" entrytime="00:01:12.00" />
                <RESULT eventid="1372" points="215" reactiontime="+101" swimtime="00:00:52.43" resultid="4025" heatid="8052" lane="7" entrytime="00:00:52.00" />
                <RESULT eventid="1569" points="139" reactiontime="+142" swimtime="00:02:53.55" resultid="4026" heatid="8124" lane="4" entrytime="00:02:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-08-19" firstname="Zofia" gender="F" lastname="Wełk" nation="POL" athleteid="4007">
              <RESULTS>
                <RESULT eventid="1090" points="107" swimtime="00:01:42.99" resultid="4008" heatid="7954" lane="5" entrytime="00:02:40.00" />
                <RESULT eventid="1181" points="66" swimtime="00:03:46.61" resultid="4009" heatid="7973" lane="1" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:45.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="137" swimtime="00:01:32.14" resultid="4010" heatid="7994" lane="6" entrytime="00:01:25.00" />
                <RESULT eventid="1357" points="72" swimtime="00:01:35.38" resultid="4011" heatid="8044" lane="7" entrytime="00:01:29.00" />
                <RESULT eventid="1387" points="248" swimtime="00:06:47.05" resultid="4012" heatid="8066" lane="4" entrytime="00:06:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:33.74" />
                    <SPLIT distance="100" swimtime="00:03:18.63" />
                    <SPLIT distance="150" swimtime="00:05:02.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="231" swimtime="00:03:06.19" resultid="4013" heatid="8118" lane="5" entrytime="00:03:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:30.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-11-25" firstname="Piotr" gender="M" lastname="Wujtiuk" nation="POL" athleteid="4027">
              <RESULTS>
                <RESULT eventid="1198" points="323" reactiontime="+78" swimtime="00:01:19.12" resultid="4028" heatid="7984" lane="9" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="209" reactiontime="+93" swimtime="00:00:51.36" resultid="4029" heatid="8001" lane="7" entrytime="00:00:50.00" />
                <RESULT eventid="1372" points="331" reactiontime="+92" swimtime="00:00:35.51" resultid="4030" heatid="8054" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="1509" points="263" reactiontime="+93" swimtime="00:03:04.80" resultid="4032" heatid="8096" lane="5" entrytime="00:02:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.88" />
                    <SPLIT distance="100" swimtime="00:01:25.96" />
                    <SPLIT distance="150" swimtime="00:02:16.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="169" reactiontime="+89" swimtime="00:00:51.45" resultid="4033" heatid="8110" lane="9" entrytime="00:00:49.00" />
                <RESULT eventid="1432" points="248" reactiontime="+93" swimtime="00:06:44.53" resultid="8290" heatid="8156" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.49" />
                    <SPLIT distance="100" swimtime="00:01:29.29" />
                    <SPLIT distance="150" swimtime="00:02:20.82" />
                    <SPLIT distance="200" swimtime="00:03:13.03" />
                    <SPLIT distance="250" swimtime="00:04:06.84" />
                    <SPLIT distance="300" swimtime="00:05:01.77" />
                    <SPLIT distance="350" swimtime="00:05:54.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" clubid="6037" name="Masters Unia Oświęcim">
          <ATHLETES>
            <ATHLETE birthdate="1966-05-03" firstname="Ilona" gender="F" lastname="Szkudlarz" athleteid="4677">
              <RESULTS>
                <RESULT eventid="1181" points="481" reactiontime="+89" swimtime="00:01:20.06" resultid="4678" heatid="7976" lane="8" entrytime="00:01:20.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="492" reactiontime="+88" swimtime="00:00:46.33" resultid="4679" heatid="7997" lane="5" entrytime="00:00:42.12" />
                <RESULT eventid="1326" points="468" reactiontime="+41" swimtime="00:01:34.05" resultid="4680" heatid="8033" lane="5" entrytime="00:01:36.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="554" reactiontime="+88" swimtime="00:00:34.51" resultid="4681" heatid="8046" lane="7" entrytime="00:00:36.40" />
                <RESULT eventid="1493" points="491" reactiontime="+89" swimtime="00:02:52.19" resultid="4682" heatid="8090" lane="8" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.40" />
                    <SPLIT distance="100" swimtime="00:01:25.93" />
                    <SPLIT distance="150" swimtime="00:02:11.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="521" reactiontime="+91" swimtime="00:01:39.53" resultid="4683" heatid="8121" lane="0" entrytime="00:01:42.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-10" firstname="Jolanta" gender="F" lastname="Płatek" athleteid="4684">
              <RESULTS>
                <RESULT eventid="1273" points="569" reactiontime="+78" swimtime="00:03:05.80" resultid="4685" heatid="8019" lane="4" entrytime="00:03:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.80" />
                    <SPLIT distance="100" swimtime="00:01:31.53" />
                    <SPLIT distance="150" swimtime="00:02:19.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="573" reactiontime="+82" swimtime="00:01:24.34" resultid="4686" heatid="8034" lane="9" entrytime="00:01:30.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="509" reactiontime="+97" swimtime="00:05:53.95" resultid="4687" heatid="8148" lane="1" entrytime="00:06:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.42" />
                    <SPLIT distance="100" swimtime="00:01:24.37" />
                    <SPLIT distance="150" swimtime="00:02:08.90" />
                    <SPLIT distance="200" swimtime="00:02:54.20" />
                    <SPLIT distance="250" swimtime="00:03:39.22" />
                    <SPLIT distance="300" swimtime="00:04:25.06" />
                    <SPLIT distance="350" swimtime="00:05:10.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="668" reactiontime="+80" swimtime="00:00:37.38" resultid="4688" heatid="8105" lane="4" entrytime="00:00:39.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="4034" name="Masters Wisła Kraków">
          <CONTACT email="wislaplywanie@gmail.com" internet="http://www.wislaplywanie.pl/sekcja-masters/" name="Wojciech Wolski" phone="791126323" />
          <ATHLETES>
            <ATHLETE birthdate="1969-01-25" firstname="Jerzy" gender="M" lastname="Korba" nation="POL" athleteid="4059">
              <RESULTS>
                <RESULT eventid="1135" points="544" reactiontime="+94" swimtime="00:10:49.32" resultid="4061" heatid="8139" lane="0" entrytime="00:11:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                    <SPLIT distance="100" swimtime="00:01:12.51" />
                    <SPLIT distance="150" swimtime="00:01:52.17" />
                    <SPLIT distance="200" swimtime="00:02:32.47" />
                    <SPLIT distance="250" swimtime="00:03:13.71" />
                    <SPLIT distance="300" swimtime="00:03:54.68" />
                    <SPLIT distance="350" swimtime="00:04:36.21" />
                    <SPLIT distance="400" swimtime="00:05:18.23" />
                    <SPLIT distance="450" swimtime="00:06:00.13" />
                    <SPLIT distance="500" swimtime="00:06:42.46" />
                    <SPLIT distance="550" swimtime="00:07:24.06" />
                    <SPLIT distance="600" swimtime="00:08:05.51" />
                    <SPLIT distance="650" swimtime="00:08:47.20" />
                    <SPLIT distance="700" swimtime="00:09:28.91" />
                    <SPLIT distance="750" swimtime="00:10:10.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="724" reactiontime="+78" swimtime="00:01:02.18" resultid="4062" heatid="7990" lane="1" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="513" reactiontime="+88" swimtime="00:00:37.35" resultid="4063" heatid="8005" lane="5" entrytime="00:00:38.00" />
                <RESULT eventid="1372" points="733" reactiontime="+78" swimtime="00:00:27.90" resultid="4064" heatid="8061" lane="2" entrytime="00:00:28.00" />
                <RESULT eventid="1599" points="607" reactiontime="+98" swimtime="00:06:08.79" resultid="4066" heatid="8164" lane="6" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.31" />
                    <SPLIT distance="100" swimtime="00:01:29.80" />
                    <SPLIT distance="150" swimtime="00:02:20.16" />
                    <SPLIT distance="200" swimtime="00:03:08.45" />
                    <SPLIT distance="250" swimtime="00:04:02.03" />
                    <SPLIT distance="300" swimtime="00:04:54.35" />
                    <SPLIT distance="350" swimtime="00:05:34.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-08-25" firstname="Tomasz" gender="M" lastname="doniec" nation="POL" athleteid="4049">
              <RESULTS>
                <RESULT eventid="1075" points="218" reactiontime="+103" swimtime="00:03:39.87" resultid="4050" heatid="7945" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.55" />
                    <SPLIT distance="100" swimtime="00:01:58.75" />
                    <SPLIT distance="150" swimtime="00:02:53.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="478" reactiontime="+95" swimtime="00:00:39.00" resultid="4051" heatid="8005" lane="3" entrytime="00:00:38.25" />
                <RESULT eventid="1402" points="352" reactiontime="+111" swimtime="00:03:33.61" resultid="4052" heatid="8074" lane="9" entrytime="00:03:25.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.45" />
                    <SPLIT distance="100" swimtime="00:01:44.07" />
                    <SPLIT distance="150" swimtime="00:02:42.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="423" reactiontime="+99" swimtime="00:01:31.53" resultid="4053" heatid="8129" lane="9" entrytime="00:01:29.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1930-05-04" firstname="Stanisław" gender="M" lastname="Krokoszyński" nation="POL" athleteid="4083">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1075" points="818" reactiontime="+118" swimtime="00:04:14.16" resultid="4084" heatid="7946" lane="0" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.38" />
                    <SPLIT distance="100" swimtime="00:02:07.03" />
                    <SPLIT distance="150" swimtime="00:03:18.71" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski, Rekord Polski" eventid="1105" points="624" reactiontime="+111" swimtime="00:01:03.73" resultid="4085" heatid="7962" lane="2" entrytime="00:01:02.00" />
                <RESULT comment="Rekord Polski" eventid="1198" points="1003" reactiontime="+121" swimtime="00:01:35.99" resultid="4086" heatid="7982" lane="8" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.33" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1228" points="758" reactiontime="+115" swimtime="00:00:56.39" resultid="4087" heatid="8000" lane="4" entrytime="00:01:00.00" />
                <RESULT comment="Rekord Polski Masters" eventid="1372" points="887" reactiontime="+111" swimtime="00:00:41.91" resultid="4088" heatid="8053" lane="0" entrytime="00:00:40.00" />
                <RESULT comment="Rekord Polski Masters" eventid="1432" points="825" reactiontime="+119" swimtime="00:08:01.90" resultid="4089" heatid="8155" lane="9" entrytime="00:07:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.02" />
                    <SPLIT distance="100" swimtime="00:01:47.49" />
                    <SPLIT distance="150" swimtime="00:02:47.74" />
                    <SPLIT distance="200" swimtime="00:03:48.83" />
                    <SPLIT distance="250" swimtime="00:04:50.83" />
                    <SPLIT distance="300" swimtime="00:05:55.70" />
                    <SPLIT distance="350" swimtime="00:06:58.86" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1509" points="987" reactiontime="+113" swimtime="00:03:36.93" resultid="4090" heatid="8096" lane="0" entrytime="00:03:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.72" />
                    <SPLIT distance="100" swimtime="00:01:38.76" />
                    <SPLIT distance="150" swimtime="00:02:37.08" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1569" points="799" reactiontime="+119" swimtime="00:02:05.66" resultid="4091" heatid="8125" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-05-16" firstname="Kamil" gender="M" lastname="Latuszek" nation="POL" athleteid="4078">
              <RESULTS>
                <RESULT eventid="1105" points="644" reactiontime="+76" swimtime="00:00:29.03" resultid="4079" heatid="7969" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1198" points="656" reactiontime="+75" swimtime="00:00:59.51" resultid="4080" heatid="7991" lane="1" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="651" reactiontime="+74" swimtime="00:00:26.71" resultid="4081" heatid="8063" lane="0" entrytime="00:00:27.00" />
                <RESULT eventid="1509" points="541" reactiontime="+70" swimtime="00:02:21.27" resultid="4082" heatid="8101" lane="9" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                    <SPLIT distance="100" swimtime="00:01:08.03" />
                    <SPLIT distance="150" swimtime="00:01:44.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-08-01" firstname="Paulina" gender="F" lastname="Palmowska" nation="POL" athleteid="4072">
              <RESULTS>
                <RESULT eventid="1058" points="647" reactiontime="+67" swimtime="00:02:49.45" resultid="4073" heatid="7944" lane="6" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.60" />
                    <SPLIT distance="100" swimtime="00:01:18.28" />
                    <SPLIT distance="150" swimtime="00:02:08.86" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1273" points="674" reactiontime="+71" swimtime="00:02:43.57" resultid="4074" heatid="8021" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                    <SPLIT distance="100" swimtime="00:01:18.04" />
                    <SPLIT distance="150" swimtime="00:02:01.43" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1326" points="793" reactiontime="+69" swimtime="00:01:14.73" resultid="4075" heatid="8035" lane="3" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1524" points="759" reactiontime="+72" swimtime="00:00:34.97" resultid="4076" heatid="8107" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1584" points="608" reactiontime="+66" swimtime="00:06:05.86" resultid="4077" heatid="8160" lane="3" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                    <SPLIT distance="100" swimtime="00:01:24.80" />
                    <SPLIT distance="150" swimtime="00:02:13.11" />
                    <SPLIT distance="200" swimtime="00:03:00.53" />
                    <SPLIT distance="250" swimtime="00:03:51.38" />
                    <SPLIT distance="300" swimtime="00:04:42.78" />
                    <SPLIT distance="350" swimtime="00:05:25.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-02-07" firstname="Bogdan" gender="M" lastname="Szczurek" nation="POL" athleteid="4118">
              <RESULTS>
                <RESULT eventid="1198" points="126" reactiontime="+154" swimtime="00:02:01.65" resultid="4119" heatid="7980" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="169" reactiontime="+139" swimtime="00:00:49.37" resultid="4120" heatid="8051" lane="5" />
                <RESULT eventid="1509" points="132" swimtime="00:04:37.77" resultid="4121" heatid="8093" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.71" />
                    <SPLIT distance="100" swimtime="00:02:03.51" />
                    <SPLIT distance="150" swimtime="00:03:16.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-11-06" firstname="Malgorzata" gender="F" lastname="Wach" nation="POL" athleteid="4114">
              <RESULTS>
                <RESULT eventid="1273" points="434" reactiontime="+69" swimtime="00:03:23.23" resultid="4115" heatid="8019" lane="1" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.48" />
                    <SPLIT distance="100" swimtime="00:01:37.02" />
                    <SPLIT distance="150" swimtime="00:02:31.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="397" reactiontime="+89" swimtime="00:06:24.47" resultid="4116" heatid="8149" lane="7" entrytime="00:07:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.72" />
                    <SPLIT distance="100" swimtime="00:01:31.45" />
                    <SPLIT distance="150" swimtime="00:02:20.91" />
                    <SPLIT distance="200" swimtime="00:03:10.33" />
                    <SPLIT distance="250" swimtime="00:03:59.96" />
                    <SPLIT distance="300" swimtime="00:04:49.56" />
                    <SPLIT distance="350" swimtime="00:05:38.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="396" reactiontime="+76" swimtime="00:03:01.50" resultid="4117" heatid="8089" lane="7" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.75" />
                    <SPLIT distance="100" swimtime="00:01:27.59" />
                    <SPLIT distance="150" swimtime="00:02:16.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-09-10" firstname="Janusz" gender="M" lastname="Mrozik" nation="POL" athleteid="4067">
              <RESULTS>
                <RESULT eventid="1288" points="172" reactiontime="+113" swimtime="00:05:04.24" resultid="4068" heatid="8022" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.43" />
                    <SPLIT distance="100" swimtime="00:02:29.17" />
                    <SPLIT distance="150" swimtime="00:03:49.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="140" reactiontime="+97" swimtime="00:02:23.66" resultid="4069" heatid="8036" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="174" reactiontime="+115" swimtime="00:05:19.96" resultid="4070" heatid="8071" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.18" />
                    <SPLIT distance="100" swimtime="00:02:33.23" />
                    <SPLIT distance="150" swimtime="00:03:59.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="133" reactiontime="+140" swimtime="00:02:35.08" resultid="4071" heatid="8124" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-08-01" firstname="Grzegorz" gender="M" lastname="Grzybczyk" nation="POL" athleteid="4099">
              <RESULTS>
                <RESULT eventid="1105" points="105" reactiontime="+113" swimtime="00:00:53.98" resultid="4100" heatid="7962" lane="0" />
                <RESULT eventid="1198" points="176" reactiontime="+92" swimtime="00:01:32.62" resultid="4101" heatid="7982" lane="0" entrytime="00:01:35.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="162" reactiontime="+99" swimtime="00:00:53.55" resultid="4102" heatid="8001" lane="0" entrytime="00:00:52.48" />
                <RESULT eventid="1342" points="100" reactiontime="+95" swimtime="00:02:13.26" resultid="4103" heatid="8037" lane="1" entrytime="00:02:03.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="197" reactiontime="+91" swimtime="00:04:19.84" resultid="4104" heatid="8071" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.69" />
                    <SPLIT distance="100" swimtime="00:02:04.26" />
                    <SPLIT distance="150" swimtime="00:03:13.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="124" reactiontime="+89" swimtime="00:00:56.49" resultid="4105" heatid="8109" lane="6" entrytime="00:00:54.59" />
                <RESULT eventid="1569" points="150" reactiontime="+101" swimtime="00:02:05.07" resultid="4106" heatid="8125" lane="3" entrytime="00:01:57.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-04" firstname="Małgorzata" gender="F" lastname="Skalska" nation="POL" athleteid="4092">
              <RESULTS>
                <RESULT eventid="1181" points="293" reactiontime="+93" swimtime="00:01:29.87" resultid="4093" heatid="7973" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="345" reactiontime="+66" swimtime="00:00:47.93" resultid="4094" heatid="7996" lane="4" entrytime="00:00:46.24" />
                <RESULT eventid="1357" points="335" reactiontime="+75" swimtime="00:00:39.49" resultid="4095" heatid="8044" lane="1" />
                <RESULT eventid="1387" points="402" reactiontime="+74" swimtime="00:03:46.52" resultid="4096" heatid="8068" lane="1" entrytime="00:03:46.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.69" />
                    <SPLIT distance="100" swimtime="00:01:50.78" />
                    <SPLIT distance="150" swimtime="00:02:49.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="257" reactiontime="+76" swimtime="00:03:28.06" resultid="4097" heatid="8089" lane="0" entrytime="00:03:18.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.89" />
                    <SPLIT distance="100" swimtime="00:01:41.58" />
                    <SPLIT distance="150" swimtime="00:02:36.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="371" reactiontime="+77" swimtime="00:01:44.86" resultid="4098" heatid="8120" lane="4" entrytime="00:01:43.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-11-11" firstname="Paulina" gender="F" lastname="Palka" nation="POL" athleteid="4054">
              <RESULTS>
                <RESULT eventid="1090" points="481" reactiontime="+72" swimtime="00:00:35.56" resultid="4055" heatid="7958" lane="6" entrytime="00:00:36.50" />
                <RESULT eventid="1273" points="595" reactiontime="+55" swimtime="00:02:52.20" resultid="4056" heatid="8021" lane="9" entrytime="00:02:52.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.08" />
                    <SPLIT distance="100" swimtime="00:01:23.37" />
                    <SPLIT distance="150" swimtime="00:02:08.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="663" reactiontime="+61" swimtime="00:01:17.45" resultid="4057" heatid="8035" lane="0" entrytime="00:01:18.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="664" reactiontime="+57" swimtime="00:00:35.75" resultid="4058" heatid="8106" lane="5" entrytime="00:00:36.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-05-28" firstname="Marta" gender="F" lastname="Wolska" nation="POL" athleteid="4042">
              <RESULTS>
                <RESULT eventid="1213" points="200" reactiontime="+132" swimtime="00:01:02.52" resultid="4043" heatid="7995" lane="7" entrytime="00:00:58.69" />
                <RESULT eventid="1273" points="212" reactiontime="+93" swimtime="00:04:26.58" resultid="4044" heatid="8018" lane="3" entrytime="00:04:18.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.05" />
                    <SPLIT distance="100" swimtime="00:02:06.43" />
                    <SPLIT distance="150" swimtime="00:03:18.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="170" reactiontime="+79" swimtime="00:02:11.73" resultid="4045" heatid="8033" lane="9" entrytime="00:01:58.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1387" points="205" reactiontime="+119" swimtime="00:04:49.67" resultid="4046" heatid="8067" lane="8" entrytime="00:04:37.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.07" />
                    <SPLIT distance="100" swimtime="00:02:19.68" />
                    <SPLIT distance="150" swimtime="00:03:34.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="192" reactiontime="+98" swimtime="00:00:57.44" resultid="4047" heatid="8104" lane="1" entrytime="00:00:56.09" />
                <RESULT eventid="1554" points="208" reactiontime="+125" swimtime="00:02:15.07" resultid="4048" heatid="8119" lane="2" entrytime="00:02:13.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-28" firstname="Wojciech" gender="M" lastname="Wolski" nation="POL" athleteid="4035">
              <RESULTS>
                <RESULT eventid="1075" points="468" reactiontime="+92" swimtime="00:03:07.81" resultid="4036" heatid="7949" lane="4" entrytime="00:02:59.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.95" />
                    <SPLIT distance="100" swimtime="00:01:30.76" />
                    <SPLIT distance="150" swimtime="00:02:23.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="306" reactiontime="+94" swimtime="00:03:26.56" resultid="4037" heatid="8013" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.16" />
                    <SPLIT distance="100" swimtime="00:01:31.20" />
                    <SPLIT distance="150" swimtime="00:02:29.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="439" reactiontime="+86" swimtime="00:03:22.15" resultid="4038" heatid="8075" lane="8" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.38" />
                    <SPLIT distance="100" swimtime="00:01:36.14" />
                    <SPLIT distance="150" swimtime="00:02:30.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="348" reactiontime="+87" swimtime="00:01:26.45" resultid="4039" heatid="8084" lane="0" entrytime="00:01:24.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="428" reactiontime="+82" swimtime="00:01:31.42" resultid="4040" heatid="8129" lane="1" entrytime="00:01:25.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="440" reactiontime="+86" swimtime="00:06:50.54" resultid="4041" heatid="8165" lane="3" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.55" />
                    <SPLIT distance="100" swimtime="00:01:31.47" />
                    <SPLIT distance="150" swimtime="00:02:29.02" />
                    <SPLIT distance="200" swimtime="00:03:26.05" />
                    <SPLIT distance="250" swimtime="00:04:20.75" />
                    <SPLIT distance="300" swimtime="00:05:15.26" />
                    <SPLIT distance="350" swimtime="00:06:01.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-08-23" firstname="Magdalena" gender="F" lastname="Drab" nation="POL" athleteid="4107">
              <RESULTS>
                <RESULT eventid="1181" points="873" reactiontime="+82" swimtime="00:01:01.38" resultid="4108" heatid="7979" lane="4" entrytime="00:01:00.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="827" reactiontime="+82" swimtime="00:00:35.79" resultid="4109" heatid="7999" lane="4" entrytime="00:00:35.64" />
                <RESULT eventid="1357" points="810" reactiontime="+78" swimtime="00:00:28.55" resultid="4110" heatid="8050" lane="6" entrytime="00:00:28.76" />
                <RESULT eventid="1387" points="816" reactiontime="+85" swimtime="00:02:48.98" resultid="4111" heatid="8070" lane="4" entrytime="00:02:48.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="100" swimtime="00:01:20.33" />
                    <SPLIT distance="150" swimtime="00:02:04.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="893" reactiontime="+81" swimtime="00:02:13.03" resultid="4112" heatid="8092" lane="5" entrytime="00:02:13.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.53" />
                    <SPLIT distance="100" swimtime="00:01:04.62" />
                    <SPLIT distance="150" swimtime="00:01:39.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="834" reactiontime="+82" swimtime="00:01:18.59" resultid="4113" heatid="8123" lane="4" entrytime="00:01:16.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="4172" name="MASTERS Zdzieszowice">
          <CONTACT name="Jajuga" />
          <ATHLETES>
            <ATHLETE birthdate="1979-02-08" firstname="Przemysław" gender="M" lastname="Osiwała" nation="POL" athleteid="4176">
              <RESULTS>
                <RESULT eventid="1105" points="478" reactiontime="+93" swimtime="00:00:32.63" resultid="4177" heatid="7970" lane="0" entrytime="00:00:29.86" />
                <RESULT eventid="1198" points="524" reactiontime="+82" swimtime="00:01:04.45" resultid="4178" heatid="7991" lane="6" entrytime="00:00:59.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="535" reactiontime="+89" swimtime="00:00:28.98" resultid="4179" heatid="8062" lane="1" entrytime="00:00:27.78" />
                <RESULT eventid="1462" status="DNS" swimtime="00:00:00.00" resultid="4180" heatid="8085" lane="1" entrytime="00:01:09.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-15" firstname="Dawid" gender="M" lastname="Jajuga" nation="POL" athleteid="4181">
              <RESULTS>
                <RESULT eventid="1165" points="487" reactiontime="+89" swimtime="00:20:56.25" resultid="4182" heatid="8143" lane="6" entrytime="00:20:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                    <SPLIT distance="100" swimtime="00:01:13.67" />
                    <SPLIT distance="150" swimtime="00:01:53.69" />
                    <SPLIT distance="200" swimtime="00:02:34.30" />
                    <SPLIT distance="250" swimtime="00:03:15.35" />
                    <SPLIT distance="300" swimtime="00:03:56.32" />
                    <SPLIT distance="350" swimtime="00:04:37.33" />
                    <SPLIT distance="400" swimtime="00:05:18.81" />
                    <SPLIT distance="450" swimtime="00:06:00.59" />
                    <SPLIT distance="500" swimtime="00:06:42.80" />
                    <SPLIT distance="550" swimtime="00:07:24.78" />
                    <SPLIT distance="600" swimtime="00:08:07.15" />
                    <SPLIT distance="650" swimtime="00:08:49.41" />
                    <SPLIT distance="700" swimtime="00:09:31.71" />
                    <SPLIT distance="750" swimtime="00:10:13.75" />
                    <SPLIT distance="800" swimtime="00:10:56.15" />
                    <SPLIT distance="850" swimtime="00:11:38.87" />
                    <SPLIT distance="900" swimtime="00:12:21.27" />
                    <SPLIT distance="950" swimtime="00:13:03.88" />
                    <SPLIT distance="1000" swimtime="00:13:45.46" />
                    <SPLIT distance="1050" swimtime="00:14:28.35" />
                    <SPLIT distance="1100" swimtime="00:15:10.82" />
                    <SPLIT distance="1150" swimtime="00:15:54.42" />
                    <SPLIT distance="1200" swimtime="00:16:37.78" />
                    <SPLIT distance="1250" swimtime="00:17:20.96" />
                    <SPLIT distance="1300" swimtime="00:18:04.31" />
                    <SPLIT distance="1350" swimtime="00:18:47.62" />
                    <SPLIT distance="1400" swimtime="00:19:30.80" />
                    <SPLIT distance="1450" swimtime="00:20:14.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="522" reactiontime="+83" swimtime="00:02:39.13" resultid="4183" heatid="8016" lane="3" entrytime="00:02:50.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                    <SPLIT distance="100" swimtime="00:01:11.90" />
                    <SPLIT distance="150" swimtime="00:01:53.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="566" reactiontime="+82" swimtime="00:05:03.22" resultid="4184" heatid="8151" lane="7" entrytime="00:04:45.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                    <SPLIT distance="100" swimtime="00:01:10.57" />
                    <SPLIT distance="150" swimtime="00:01:48.44" />
                    <SPLIT distance="200" swimtime="00:02:27.41" />
                    <SPLIT distance="250" swimtime="00:03:05.61" />
                    <SPLIT distance="300" swimtime="00:03:44.08" />
                    <SPLIT distance="350" swimtime="00:04:23.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="601" reactiontime="+76" swimtime="00:05:38.01" resultid="4185" heatid="8163" lane="6" entrytime="00:05:55.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                    <SPLIT distance="100" swimtime="00:01:09.55" />
                    <SPLIT distance="150" swimtime="00:01:54.42" />
                    <SPLIT distance="200" swimtime="00:02:37.76" />
                    <SPLIT distance="250" swimtime="00:03:26.78" />
                    <SPLIT distance="300" swimtime="00:04:16.79" />
                    <SPLIT distance="350" swimtime="00:04:57.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="4122" name="Masters Łódź">
          <CONTACT email="sport@masterslodz.pl" internet="http://masterslodz.pl" name="Trudnos Rafał" />
          <ATHLETES>
            <ATHLETE birthdate="1983-01-01" firstname="Jakub" gender="M" lastname="Sidorowicz" nation="POL" athleteid="4141">
              <RESULTS>
                <RESULT eventid="1075" points="228" reactiontime="+84" swimtime="00:03:35.27" resultid="4142" heatid="7950" lane="9" entrytime="00:02:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.20" />
                    <SPLIT distance="100" swimtime="00:01:40.02" />
                    <SPLIT distance="150" swimtime="00:02:42.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" status="DNS" swimtime="00:00:00.00" resultid="4143" heatid="8004" lane="9" entrytime="00:00:42.00" />
                <RESULT eventid="1342" status="DNS" swimtime="00:00:00.00" resultid="4144" heatid="8038" lane="1" entrytime="00:01:40.00" />
                <RESULT eventid="1402" status="DNS" swimtime="00:00:00.00" resultid="4145" heatid="8074" lane="4" entrytime="00:03:10.15" />
                <RESULT eventid="1539" points="222" reactiontime="+72" swimtime="00:00:42.93" resultid="4146" heatid="8112" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1569" points="258" reactiontime="+106" swimtime="00:01:42.31" resultid="4147" heatid="8127" lane="0" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-01" firstname="Artur" gender="M" lastname="Frąckowiak" nation="POL" athleteid="4163">
              <RESULTS>
                <RESULT eventid="1075" points="617" reactiontime="+85" swimtime="00:02:38.64" resultid="4164" heatid="7950" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                    <SPLIT distance="100" swimtime="00:01:14.68" />
                    <SPLIT distance="150" swimtime="00:02:01.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="596" reactiontime="+81" swimtime="00:00:30.32" resultid="4165" heatid="7968" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="1198" points="586" reactiontime="+81" swimtime="00:01:02.10" resultid="4166" heatid="7989" lane="6" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="465" reactiontime="+79" swimtime="00:00:37.69" resultid="4167" heatid="8006" lane="4" entrytime="00:00:37.00" />
                <RESULT eventid="1372" points="590" reactiontime="+73" swimtime="00:00:28.04" resultid="4168" heatid="8061" lane="3" entrytime="00:00:28.00" />
                <RESULT eventid="1432" points="522" reactiontime="+92" swimtime="00:05:18.56" resultid="4169" heatid="8153" lane="6" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                    <SPLIT distance="100" swimtime="00:01:09.23" />
                    <SPLIT distance="150" swimtime="00:01:48.89" />
                    <SPLIT distance="200" swimtime="00:02:29.94" />
                    <SPLIT distance="250" swimtime="00:03:11.87" />
                    <SPLIT distance="300" swimtime="00:03:54.87" />
                    <SPLIT distance="350" swimtime="00:04:37.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="532" reactiontime="+80" swimtime="00:02:22.75" resultid="4170" heatid="8099" lane="7" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                    <SPLIT distance="100" swimtime="00:01:07.85" />
                    <SPLIT distance="150" swimtime="00:01:46.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-01" firstname="Jakub" gender="M" lastname="Karczmarczyk" nation="POL" athleteid="4157">
              <RESULTS>
                <RESULT eventid="1075" points="414" reactiontime="+103" swimtime="00:03:01.26" resultid="4158" heatid="7949" lane="1" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.81" />
                    <SPLIT distance="100" swimtime="00:01:24.45" />
                    <SPLIT distance="150" swimtime="00:02:18.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="423" reactiontime="+92" swimtime="00:00:38.90" resultid="4159" heatid="8004" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="1372" points="483" reactiontime="+90" swimtime="00:00:29.99" resultid="4160" heatid="8055" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="1402" points="468" reactiontime="+91" swimtime="00:03:14.95" resultid="4161" heatid="8074" lane="3" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.78" />
                    <SPLIT distance="100" swimtime="00:01:33.17" />
                    <SPLIT distance="150" swimtime="00:02:25.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="447" reactiontime="+87" swimtime="00:01:26.87" resultid="4162" heatid="8128" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-01" firstname="Jakub" gender="M" lastname="Gryczyński" nation="POL" athleteid="4148">
              <RESULTS>
                <RESULT eventid="1228" status="DNS" swimtime="00:00:00.00" resultid="4149" heatid="8004" lane="7" entrytime="00:00:41.00" />
                <RESULT eventid="1372" points="424" reactiontime="+85" swimtime="00:00:31.32" resultid="4150" heatid="8056" lane="5" entrytime="00:00:31.00" />
                <RESULT eventid="1569" points="347" reactiontime="+84" swimtime="00:01:34.52" resultid="4151" heatid="8127" lane="4" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-01" firstname="Arkadiusz" gender="M" lastname="Olkowicz" nation="POL" athleteid="4130">
              <RESULTS>
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="4131" heatid="7969" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1135" points="431" reactiontime="+79" swimtime="00:11:48.72" resultid="4132" heatid="8140" lane="5" entrytime="00:11:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                    <SPLIT distance="100" swimtime="00:01:17.12" />
                    <SPLIT distance="150" swimtime="00:01:58.59" />
                    <SPLIT distance="200" swimtime="00:02:41.70" />
                    <SPLIT distance="250" swimtime="00:03:26.02" />
                    <SPLIT distance="300" swimtime="00:04:11.66" />
                    <SPLIT distance="350" swimtime="00:04:57.82" />
                    <SPLIT distance="400" swimtime="00:05:43.67" />
                    <SPLIT distance="450" swimtime="00:06:29.66" />
                    <SPLIT distance="500" swimtime="00:07:15.78" />
                    <SPLIT distance="550" swimtime="00:08:01.39" />
                    <SPLIT distance="600" swimtime="00:08:48.56" />
                    <SPLIT distance="650" swimtime="00:09:34.81" />
                    <SPLIT distance="700" swimtime="00:10:21.37" />
                    <SPLIT distance="750" swimtime="00:11:05.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="344" reactiontime="+78" swimtime="00:00:33.56" resultid="4133" heatid="8060" lane="6" entrytime="00:00:28.50" />
                <RESULT eventid="1432" status="DNS" swimtime="00:00:00.00" resultid="4134" heatid="8153" lane="3" entrytime="00:05:30.00" />
                <RESULT eventid="1539" points="473" reactiontime="+82" swimtime="00:00:36.19" resultid="4135" heatid="8113" lane="5" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-01" firstname="Wojciech" gender="M" lastname="Zdzieszyński" nation="POL" athleteid="4136">
              <RESULTS>
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="4137" heatid="7969" lane="8" entrytime="00:00:31.00" />
                <RESULT eventid="1198" points="540" reactiontime="+96" swimtime="00:01:03.81" resultid="4138" heatid="7990" lane="4" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="653" reactiontime="+90" swimtime="00:00:27.11" resultid="4139" heatid="8064" lane="3" entrytime="00:00:26.00" />
                <RESULT eventid="1509" points="342" reactiontime="+98" swimtime="00:02:45.33" resultid="4140" heatid="8101" lane="7" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                    <SPLIT distance="100" swimtime="00:01:11.26" />
                    <SPLIT distance="150" swimtime="00:01:57.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-01" firstname="Łukasz" gender="M" lastname="Raj" nation="POL" athleteid="4152">
              <RESULTS>
                <RESULT eventid="1198" points="323" reactiontime="+85" swimtime="00:01:15.75" resultid="4153" heatid="7988" lane="2" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" status="DNS" swimtime="00:00:00.00" resultid="4154" heatid="8006" lane="3" entrytime="00:00:37.00" />
                <RESULT comment="O4 - Start wykonany przed sygnałem (przedwczesny start)" eventid="1372" reactiontime="+48" status="DSQ" swimtime="00:00:31.57" resultid="4155" heatid="8061" lane="5" entrytime="00:00:28.00" />
                <RESULT eventid="1539" points="335" reactiontime="+94" swimtime="00:00:40.60" resultid="4156" heatid="8113" lane="3" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1318" reactiontime="+81" swimtime="00:04:23.72" resultid="4171" heatid="8030" lane="6" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.68" />
                    <SPLIT distance="100" swimtime="00:01:02.48" />
                    <SPLIT distance="150" swimtime="00:01:35.06" />
                    <SPLIT distance="200" swimtime="00:02:12.19" />
                    <SPLIT distance="250" swimtime="00:02:44.31" />
                    <SPLIT distance="300" swimtime="00:03:00.11" />
                    <SPLIT distance="350" swimtime="00:03:49.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4163" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="4157" number="2" reactiontime="+79" />
                    <RELAYPOSITION athleteid="4130" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="4136" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2190" name="MKP Szczecin">
          <CONTACT email="windmuhle@wp.pl" name="Kowalczyk Piotr" />
          <ATHLETES>
            <ATHLETE birthdate="1966-08-10" firstname="Małgorzata" gender="F" lastname="Serbin" nation="POL" athleteid="3020">
              <RESULTS>
                <RESULT eventid="1120" points="683" reactiontime="+76" swimtime="00:10:59.21" resultid="3021" heatid="8136" lane="6" entrytime="00:10:41.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                    <SPLIT distance="100" swimtime="00:01:16.21" />
                    <SPLIT distance="150" swimtime="00:01:56.95" />
                    <SPLIT distance="200" swimtime="00:02:38.70" />
                    <SPLIT distance="250" swimtime="00:03:20.37" />
                    <SPLIT distance="300" swimtime="00:04:02.26" />
                    <SPLIT distance="350" swimtime="00:04:44.06" />
                    <SPLIT distance="400" swimtime="00:05:26.12" />
                    <SPLIT distance="450" swimtime="00:06:08.05" />
                    <SPLIT distance="500" swimtime="00:06:50.36" />
                    <SPLIT distance="550" swimtime="00:07:32.38" />
                    <SPLIT distance="600" swimtime="00:08:14.53" />
                    <SPLIT distance="650" swimtime="00:08:56.76" />
                    <SPLIT distance="700" swimtime="00:09:38.81" />
                    <SPLIT distance="750" swimtime="00:10:20.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="704" reactiontime="+77" swimtime="00:02:58.91" resultid="3022" heatid="8020" lane="5" entrytime="00:02:54.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.47" />
                    <SPLIT distance="100" swimtime="00:01:27.89" />
                    <SPLIT distance="150" swimtime="00:02:14.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="647" reactiontime="+78" swimtime="00:05:28.70" resultid="3023" heatid="8147" lane="6" entrytime="00:05:09.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.60" />
                    <SPLIT distance="100" swimtime="00:01:17.48" />
                    <SPLIT distance="150" swimtime="00:01:59.46" />
                    <SPLIT distance="200" swimtime="00:02:42.16" />
                    <SPLIT distance="250" swimtime="00:03:24.83" />
                    <SPLIT distance="300" swimtime="00:04:07.71" />
                    <SPLIT distance="350" swimtime="00:04:49.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-10-31" firstname="Konrad" gender="M" lastname="Tekiel" nation="POL" athleteid="3025">
              <RESULTS>
                <RESULT eventid="1372" status="DNS" swimtime="00:00:00.00" resultid="3026" heatid="8052" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-05-23" firstname="Paweł" gender="M" lastname="Radziński" nation="POL" athleteid="2198">
              <RESULTS>
                <RESULT eventid="1432" points="639" reactiontime="+79" swimtime="00:04:51.25" resultid="2201" heatid="8151" lane="3" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                    <SPLIT distance="100" swimtime="00:01:07.13" />
                    <SPLIT distance="150" swimtime="00:01:45.00" />
                    <SPLIT distance="200" swimtime="00:02:22.82" />
                    <SPLIT distance="250" swimtime="00:03:00.44" />
                    <SPLIT distance="300" swimtime="00:03:38.40" />
                    <SPLIT distance="350" swimtime="00:04:15.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="674" reactiontime="+80" swimtime="00:02:11.28" resultid="2202" heatid="8102" lane="2" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.39" />
                    <SPLIT distance="100" swimtime="00:01:02.01" />
                    <SPLIT distance="150" swimtime="00:01:36.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="642" reactiontime="+89" swimtime="00:10:04.10" resultid="3001" heatid="8139" lane="4" entrytime="00:09:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.67" />
                    <SPLIT distance="100" swimtime="00:01:14.16" />
                    <SPLIT distance="150" swimtime="00:01:51.95" />
                    <SPLIT distance="200" swimtime="00:02:30.26" />
                    <SPLIT distance="250" swimtime="00:03:08.47" />
                    <SPLIT distance="300" swimtime="00:03:46.40" />
                    <SPLIT distance="350" swimtime="00:04:24.36" />
                    <SPLIT distance="400" swimtime="00:05:02.49" />
                    <SPLIT distance="450" swimtime="00:05:42.43" />
                    <SPLIT distance="500" swimtime="00:06:20.50" />
                    <SPLIT distance="550" swimtime="00:06:58.32" />
                    <SPLIT distance="600" swimtime="00:07:36.37" />
                    <SPLIT distance="650" swimtime="00:08:14.33" />
                    <SPLIT distance="700" swimtime="00:08:52.23" />
                    <SPLIT distance="750" swimtime="00:09:28.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-02" firstname="Piotr" gender="M" lastname="Kowalczyk" nation="POL" athleteid="3012">
              <RESULTS>
                <RESULT eventid="1135" points="566" reactiontime="+83" swimtime="00:10:36.28" resultid="3013" heatid="8139" lane="6" entrytime="00:10:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                    <SPLIT distance="100" swimtime="00:01:12.65" />
                    <SPLIT distance="150" swimtime="00:01:51.97" />
                    <SPLIT distance="200" swimtime="00:02:32.34" />
                    <SPLIT distance="250" swimtime="00:03:12.33" />
                    <SPLIT distance="300" swimtime="00:03:52.55" />
                    <SPLIT distance="350" swimtime="00:04:32.87" />
                    <SPLIT distance="400" swimtime="00:05:13.08" />
                    <SPLIT distance="450" swimtime="00:05:53.58" />
                    <SPLIT distance="500" swimtime="00:06:34.60" />
                    <SPLIT distance="550" swimtime="00:07:15.61" />
                    <SPLIT distance="600" swimtime="00:07:56.44" />
                    <SPLIT distance="650" swimtime="00:08:37.88" />
                    <SPLIT distance="700" swimtime="00:09:19.05" />
                    <SPLIT distance="750" swimtime="00:09:58.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="3014" heatid="8026" lane="9" entrytime="00:02:54.00" />
                <RESULT eventid="1432" points="609" reactiontime="+81" swimtime="00:05:00.00" resultid="3015" heatid="8152" lane="5" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                    <SPLIT distance="100" swimtime="00:01:09.65" />
                    <SPLIT distance="150" swimtime="00:01:48.05" />
                    <SPLIT distance="200" swimtime="00:02:27.08" />
                    <SPLIT distance="250" swimtime="00:03:06.16" />
                    <SPLIT distance="300" swimtime="00:03:45.32" />
                    <SPLIT distance="350" swimtime="00:04:24.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-07-26" firstname="Marcin" gender="M" lastname="Gargas" nation="POL" athleteid="3028">
              <RESULTS>
                <RESULT eventid="1372" status="DNS" swimtime="00:00:00.00" resultid="6000" heatid="8054" lane="8" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1935-01-01" firstname="Stefania" gender="F" lastname="Noetzel" nation="POL" athleteid="3016">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1213" points="448" swimtime="00:01:09.73" resultid="3017" heatid="7994" lane="3" entrytime="00:01:10.07" />
                <RESULT comment="Rekord Polski Masters" eventid="1387" points="836" swimtime="00:04:57.21" resultid="3018" heatid="8067" lane="0" entrytime="00:04:58.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.51" />
                    <SPLIT distance="100" swimtime="00:02:23.17" />
                    <SPLIT distance="150" swimtime="00:03:42.37" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1554" points="780" swimtime="00:02:20.32" resultid="3019" heatid="8119" lane="8" entrytime="00:02:21.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-02-09" firstname="Piotr" gender="M" lastname="Nowicki" nation="POL" athleteid="3029">
              <RESULTS>
                <RESULT eventid="1372" status="DNS" swimtime="00:00:00.00" resultid="3030" heatid="8053" lane="5" entrytime="00:00:38.00" />
                <RESULT eventid="1509" status="DNS" swimtime="00:00:00.00" resultid="3032" heatid="8096" lane="9" entrytime="00:03:07.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-09-25" firstname="Sławomir" gender="M" lastname="Grzeszewski" nation="POL" athleteid="3002">
              <RESULTS>
                <RESULT eventid="1075" points="550" reactiontime="+86" swimtime="00:03:18.16" resultid="3003" heatid="7947" lane="3" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                    <SPLIT distance="100" swimtime="00:01:34.84" />
                    <SPLIT distance="150" swimtime="00:02:31.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="578" reactiontime="+67" swimtime="00:00:41.23" resultid="3004" heatid="8002" lane="7" entrytime="00:00:45.00" />
                <RESULT eventid="1402" points="552" reactiontime="+68" swimtime="00:03:38.06" resultid="3005" heatid="8073" lane="9" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.80" />
                    <SPLIT distance="100" swimtime="00:01:43.26" />
                    <SPLIT distance="150" swimtime="00:02:40.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="522" reactiontime="+56" swimtime="00:01:38.46" resultid="3006" heatid="8127" lane="9" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-02-27" firstname="Szymon" gender="M" lastname="Kluczyk" nation="POL" athleteid="3007">
              <RESULTS>
                <RESULT eventid="1165" points="528" reactiontime="+95" swimtime="00:20:22.64" resultid="3008" heatid="8143" lane="5" entrytime="00:19:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.38" />
                    <SPLIT distance="100" swimtime="00:01:12.35" />
                    <SPLIT distance="150" swimtime="00:01:51.15" />
                    <SPLIT distance="200" swimtime="00:02:30.56" />
                    <SPLIT distance="250" swimtime="00:03:10.66" />
                    <SPLIT distance="300" swimtime="00:03:51.04" />
                    <SPLIT distance="350" swimtime="00:04:31.47" />
                    <SPLIT distance="400" swimtime="00:05:12.48" />
                    <SPLIT distance="450" swimtime="00:05:53.24" />
                    <SPLIT distance="500" swimtime="00:06:34.43" />
                    <SPLIT distance="550" swimtime="00:07:15.26" />
                    <SPLIT distance="600" swimtime="00:07:56.69" />
                    <SPLIT distance="650" swimtime="00:08:37.96" />
                    <SPLIT distance="700" swimtime="00:09:19.60" />
                    <SPLIT distance="750" swimtime="00:10:01.21" />
                    <SPLIT distance="800" swimtime="00:10:42.72" />
                    <SPLIT distance="850" swimtime="00:11:23.85" />
                    <SPLIT distance="900" swimtime="00:12:05.41" />
                    <SPLIT distance="950" swimtime="00:12:46.67" />
                    <SPLIT distance="1000" swimtime="00:13:28.44" />
                    <SPLIT distance="1050" swimtime="00:14:10.30" />
                    <SPLIT distance="1100" swimtime="00:14:51.61" />
                    <SPLIT distance="1150" swimtime="00:15:32.79" />
                    <SPLIT distance="1200" swimtime="00:16:14.55" />
                    <SPLIT distance="1250" swimtime="00:16:56.08" />
                    <SPLIT distance="1300" swimtime="00:17:37.57" />
                    <SPLIT distance="1350" swimtime="00:18:19.14" />
                    <SPLIT distance="1400" swimtime="00:19:00.58" />
                    <SPLIT distance="1450" swimtime="00:19:43.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="464" reactiontime="+97" swimtime="00:02:45.52" resultid="3009" heatid="8017" lane="0" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                    <SPLIT distance="100" swimtime="00:01:15.18" />
                    <SPLIT distance="150" swimtime="00:02:04.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="710" reactiontime="+90" swimtime="00:04:41.23" resultid="3010" heatid="8151" lane="1" entrytime="00:04:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                    <SPLIT distance="100" swimtime="00:01:05.40" />
                    <SPLIT distance="150" swimtime="00:01:40.06" />
                    <SPLIT distance="200" swimtime="00:02:15.72" />
                    <SPLIT distance="250" swimtime="00:02:51.71" />
                    <SPLIT distance="300" swimtime="00:03:28.76" />
                    <SPLIT distance="350" swimtime="00:04:05.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="679" reactiontime="+89" swimtime="00:05:24.61" resultid="3011" heatid="8162" lane="6" entrytime="00:05:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                    <SPLIT distance="100" swimtime="00:01:10.92" />
                    <SPLIT distance="150" swimtime="00:01:54.04" />
                    <SPLIT distance="200" swimtime="00:02:35.99" />
                    <SPLIT distance="250" swimtime="00:03:25.10" />
                    <SPLIT distance="300" swimtime="00:04:14.16" />
                    <SPLIT distance="350" swimtime="00:04:49.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="4194" name="MKS Aquatic Gubin">
          <CONTACT name="Ziemowit Patek" />
          <ATHLETES>
            <ATHLETE birthdate="1975-03-29" firstname="Sylwia" gender="F" lastname="Gorockiewicz" nation="POL" athleteid="4199">
              <RESULTS>
                <RESULT eventid="1213" points="234" reactiontime="+99" swimtime="00:00:56.68" resultid="4200" heatid="7995" lane="8" entrytime="00:01:03.69" />
                <RESULT eventid="1387" points="246" reactiontime="+119" swimtime="00:04:31.11" resultid="4201" heatid="8066" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.84" />
                    <SPLIT distance="100" swimtime="00:02:09.49" />
                    <SPLIT distance="150" swimtime="00:03:21.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="222" reactiontime="+114" swimtime="00:02:06.74" resultid="4202" heatid="8119" lane="7" entrytime="00:02:18.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Anna" gender="F" lastname="Krupińska" nation="POL" athleteid="4195">
              <RESULTS>
                <RESULT eventid="1213" points="449" reactiontime="+96" swimtime="00:00:50.22" resultid="4196" heatid="7996" lane="8" entrytime="00:00:49.00" />
                <RESULT eventid="1387" points="539" reactiontime="+104" swimtime="00:04:00.93" resultid="4197" heatid="8067" lane="5" entrytime="00:03:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.04" />
                    <SPLIT distance="100" swimtime="00:01:57.89" />
                    <SPLIT distance="150" swimtime="00:03:00.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="521" reactiontime="+115" swimtime="00:01:51.64" resultid="4198" heatid="8120" lane="1" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00816" nation="POL" region="SZ" clubid="4203" name="MKS Neptun Stargard">
          <CONTACT city="Stargard Szcz." email="prezes@mksneptun.pl" internet="www.mksneptun.pl" name="Miedzyszkolny Klub Sportowy &quot;Neptun&quot;" phone="602731410" state="ZACHO" street="Os. Zachód B 15" zip="73-110" />
          <ATHLETES>
            <ATHLETE birthdate="1972-08-18" firstname="Ireneusz" gender="M" lastname="Drozd" nation="POL" athleteid="4211">
              <RESULTS>
                <RESULT eventid="1105" points="592" reactiontime="+97" swimtime="00:00:30.83" resultid="4212" heatid="7969" lane="2" entrytime="00:00:30.04" />
                <RESULT eventid="1342" status="DNS" swimtime="00:00:00.00" resultid="4213" heatid="8041" lane="6" entrytime="00:01:14.04" />
                <RESULT eventid="1372" status="DNS" swimtime="00:00:00.00" resultid="4214" heatid="8060" lane="0" entrytime="00:00:28.74" />
                <RESULT eventid="1539" status="DNS" swimtime="00:00:00.00" resultid="4215" heatid="8114" lane="4" entrytime="00:00:33.44" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-09-30" firstname="Mateusz" gender="M" lastname="Drozd" nation="POL" athleteid="4204">
              <RESULTS>
                <RESULT eventid="1075" points="788" reactiontime="+74" swimtime="00:02:20.29" resultid="4205" heatid="7953" lane="5" entrytime="00:02:15.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.33" />
                    <SPLIT distance="100" swimtime="00:01:05.25" />
                    <SPLIT distance="150" swimtime="00:01:47.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="814" reactiontime="+70" swimtime="00:00:27.04" resultid="4206" heatid="7972" lane="6" entrytime="00:00:26.20" />
                <RESULT eventid="1198" points="831" reactiontime="+71" swimtime="00:00:55.01" resultid="4207" heatid="7993" lane="5" entrytime="00:00:54.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="647" reactiontime="+82" swimtime="00:01:07.47" resultid="4208" heatid="8043" lane="4" entrytime="00:01:01.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="793" reactiontime="+69" swimtime="00:00:24.88" resultid="4209" heatid="8065" lane="2" entrytime="00:00:24.73" />
                <RESULT eventid="1539" points="739" reactiontime="+75" swimtime="00:00:30.14" resultid="4210" heatid="8117" lane="3" entrytime="00:00:28.62" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="01011" nation="POL" region="SLA" clubid="4216" name="MKS Park Wodny Tarnowskie Góry">
          <CONTACT city="Tarnowskie Góry" email="klubplywacki@gmail.com" name="Macner Dagmara" phone="509 691 784" state="SLA" street="ul. Obwodnica 8" zip="42-600" />
          <ATHLETES>
            <ATHLETE birthdate="1989-07-15" firstname="Mateusz" gender="M" lastname="Kotkowski" nation="POL" athleteid="4217">
              <RESULTS>
                <RESULT eventid="1105" points="697" reactiontime="+75" swimtime="00:00:28.27" resultid="4218" heatid="7971" lane="5" entrytime="00:00:28.00" />
                <RESULT eventid="1198" points="704" reactiontime="+79" swimtime="00:00:58.12" resultid="4219" heatid="7993" lane="9" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="703" reactiontime="+74" swimtime="00:00:26.03" resultid="4220" heatid="8064" lane="5" entrytime="00:00:26.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-12-31" firstname="Kajetan" gender="M" lastname="Smoliński" nation="POL" athleteid="4221">
              <RESULTS>
                <RESULT eventid="1105" points="693" reactiontime="+76" swimtime="00:00:28.33" resultid="4222" heatid="7970" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="1372" points="708" reactiontime="+72" swimtime="00:00:25.97" resultid="4223" heatid="8065" lane="1" entrytime="00:00:25.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2104" name="MOSiR KSZO Ostrowiec Św.">
          <CONTACT name="Różalski Zbigniew" />
          <ATHLETES>
            <ATHLETE birthdate="1945-03-28" firstname="Józef" gender="M" lastname="Różalski" nation="POL" athleteid="2105">
              <RESULTS>
                <RESULT eventid="1075" points="716" reactiontime="+94" swimtime="00:03:22.84" resultid="2106" heatid="7946" lane="4" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.25" />
                    <SPLIT distance="100" swimtime="00:01:36.79" />
                    <SPLIT distance="150" swimtime="00:02:38.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="783" reactiontime="+93" swimtime="00:00:36.33" resultid="2107" heatid="7964" lane="1" entrytime="00:00:38.00" />
                <RESULT eventid="1198" points="594" reactiontime="+91" swimtime="00:01:18.28" resultid="2108" heatid="7983" lane="8" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="659" reactiontime="+91" swimtime="00:00:43.80" resultid="2109" heatid="8002" lane="4" entrytime="00:00:44.00" />
                <RESULT eventid="1372" points="624" reactiontime="+90" swimtime="00:00:33.30" resultid="2110" heatid="8055" lane="8" entrytime="00:00:34.00" />
                <RESULT eventid="1462" points="460" reactiontime="+96" swimtime="00:01:42.89" resultid="2111" heatid="8082" lane="6" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="515" reactiontime="+108" swimtime="00:03:10.71" resultid="2112" heatid="8095" lane="5" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                    <SPLIT distance="100" swimtime="00:01:30.89" />
                    <SPLIT distance="150" swimtime="00:02:21.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="617" reactiontime="+94" swimtime="00:01:42.05" resultid="2113" heatid="8127" lane="8" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOTYL" nation="POL" region="PDK" clubid="4228" name="MOTYL-SENIOR MOSiR Stalowa Wola" shortname="MOTYL -SENIOR MOSiR Stalowa Wo">
          <CONTACT city="Stalowa Wola" email="lorkowska@wp.pl" name="Chmielewski Andrzej" state="PODK" street="Hutnicza 15" zip="37-450" />
          <ATHLETES>
            <ATHLETE birthdate="1967-04-17" firstname="Maria" gender="F" lastname="Petecka" nation="POL" athleteid="4260">
              <RESULTS>
                <RESULT eventid="1058" points="536" reactiontime="+91" swimtime="00:03:12.94" resultid="4261" heatid="7943" lane="0" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.39" />
                    <SPLIT distance="100" swimtime="00:01:35.45" />
                    <SPLIT distance="150" swimtime="00:02:29.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="511" reactiontime="+90" swimtime="00:00:37.90" resultid="4262" heatid="7957" lane="1" entrytime="00:00:39.00" />
                <RESULT eventid="1243" points="363" reactiontime="+95" swimtime="00:03:40.60" resultid="4263" heatid="8012" lane="0" entrytime="00:03:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.95" />
                    <SPLIT distance="100" swimtime="00:01:40.60" />
                    <SPLIT distance="150" swimtime="00:02:38.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1387" points="494" reactiontime="+86" swimtime="00:03:36.14" resultid="4264" heatid="8068" lane="5" entrytime="00:03:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.61" />
                    <SPLIT distance="100" swimtime="00:01:45.34" />
                    <SPLIT distance="150" swimtime="00:02:41.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="359" reactiontime="+89" swimtime="00:01:37.90" resultid="4265" heatid="8078" lane="4" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="443" reactiontime="+91" swimtime="00:02:58.15" resultid="4266" heatid="8089" lane="3" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.45" />
                    <SPLIT distance="100" swimtime="00:01:22.82" />
                    <SPLIT distance="150" swimtime="00:02:10.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="528" reactiontime="+90" swimtime="00:01:39.07" resultid="4267" heatid="8120" lane="3" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-14" firstname="Arkadiusz" gender="M" lastname="Berwecki" nation="POL" athleteid="4229">
              <RESULTS>
                <RESULT eventid="1075" points="821" reactiontime="+73" swimtime="00:02:21.39" resultid="4230" heatid="7953" lane="2" entrytime="00:02:20.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.03" />
                    <SPLIT distance="100" swimtime="00:01:06.17" />
                    <SPLIT distance="150" swimtime="00:01:47.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="820" reactiontime="+71" swimtime="00:00:27.67" resultid="4231" heatid="7972" lane="8" entrytime="00:00:27.59" />
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1198" points="876" reactiontime="+73" swimtime="00:00:56.75" resultid="4232" heatid="7993" lane="7" entrytime="00:00:57.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="702" reactiontime="+80" swimtime="00:02:28.87" resultid="4233" heatid="8017" lane="3" entrytime="00:02:23.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                    <SPLIT distance="100" swimtime="00:01:08.36" />
                    <SPLIT distance="150" swimtime="00:01:46.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="807" reactiontime="+72" swimtime="00:00:26.40" resultid="4234" heatid="8063" lane="4" entrytime="00:00:26.29" />
                <RESULT eventid="1462" points="902" reactiontime="+68" swimtime="00:01:00.73" resultid="4235" heatid="8086" lane="6" entrytime="00:01:00.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="826" reactiontime="+73" swimtime="00:02:06.25" resultid="4236" heatid="8102" lane="5" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.15" />
                    <SPLIT distance="100" swimtime="00:01:01.37" />
                    <SPLIT distance="150" swimtime="00:01:34.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="699" reactiontime="+79" swimtime="00:05:18.88" resultid="4237" heatid="8162" lane="5" entrytime="00:05:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                    <SPLIT distance="100" swimtime="00:01:10.98" />
                    <SPLIT distance="150" swimtime="00:01:51.73" />
                    <SPLIT distance="200" swimtime="00:02:31.79" />
                    <SPLIT distance="250" swimtime="00:03:18.07" />
                    <SPLIT distance="300" swimtime="00:04:04.31" />
                    <SPLIT distance="350" swimtime="00:04:42.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-02-27" firstname="Robert" gender="M" lastname="Lorkowski" nation="POL" athleteid="4254">
              <RESULTS>
                <RESULT eventid="1075" points="749" reactiontime="+92" swimtime="00:02:50.68" resultid="4255" heatid="7950" lane="6" entrytime="00:02:53.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.92" />
                    <SPLIT distance="100" swimtime="00:01:20.49" />
                    <SPLIT distance="150" swimtime="00:02:11.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="701" reactiontime="+93" swimtime="00:01:08.37" resultid="4256" heatid="7986" lane="2" entrytime="00:01:08.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="748" reactiontime="+77" swimtime="00:02:56.39" resultid="4257" heatid="8025" lane="1" entrytime="00:03:02.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                    <SPLIT distance="100" swimtime="00:01:23.31" />
                    <SPLIT distance="150" swimtime="00:02:09.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="742" reactiontime="+76" swimtime="00:01:19.49" resultid="4258" heatid="8040" lane="9" entrytime="00:01:20.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="710" reactiontime="+89" swimtime="00:06:12.81" resultid="4259" heatid="8164" lane="3" entrytime="00:06:18.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.57" />
                    <SPLIT distance="100" swimtime="00:01:28.02" />
                    <SPLIT distance="150" swimtime="00:02:15.46" />
                    <SPLIT distance="200" swimtime="00:03:02.08" />
                    <SPLIT distance="250" swimtime="00:03:56.27" />
                    <SPLIT distance="300" swimtime="00:04:50.52" />
                    <SPLIT distance="350" swimtime="00:05:32.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-08-09" firstname="Włodzimierz" gender="M" lastname="Jarzyna" nation="POL" athleteid="4238">
              <RESULTS>
                <RESULT eventid="1075" points="569" reactiontime="+87" swimtime="00:03:19.85" resultid="4239" heatid="7947" lane="6" entrytime="00:03:31.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.85" />
                    <SPLIT distance="100" swimtime="00:01:38.73" />
                    <SPLIT distance="150" swimtime="00:02:37.68" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1288" points="520" reactiontime="+72" swimtime="00:03:20.15" resultid="4240" heatid="8024" lane="7" entrytime="00:03:33.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.87" />
                    <SPLIT distance="100" swimtime="00:01:36.32" />
                    <SPLIT distance="150" swimtime="00:02:30.96" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1342" points="556" reactiontime="+73" swimtime="00:01:29.74" resultid="4241" heatid="8038" lane="2" entrytime="00:01:35.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="637" reactiontime="+107" swimtime="00:06:13.31" resultid="4242" heatid="8155" lane="4" entrytime="00:06:31.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.92" />
                    <SPLIT distance="100" swimtime="00:01:27.76" />
                    <SPLIT distance="150" swimtime="00:02:16.81" />
                    <SPLIT distance="200" swimtime="00:03:05.76" />
                    <SPLIT distance="250" swimtime="00:03:55.70" />
                    <SPLIT distance="300" swimtime="00:04:44.10" />
                    <SPLIT distance="350" swimtime="00:05:31.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="529" reactiontime="+76" swimtime="00:00:41.42" resultid="4243" heatid="8111" lane="9" entrytime="00:00:44.09" />
                <RESULT eventid="1599" points="704" reactiontime="+100" swimtime="00:07:04.06" resultid="4244" heatid="8166" lane="4" entrytime="00:07:20.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.85" />
                    <SPLIT distance="100" swimtime="00:01:48.50" />
                    <SPLIT distance="150" swimtime="00:02:43.92" />
                    <SPLIT distance="200" swimtime="00:03:34.35" />
                    <SPLIT distance="250" swimtime="00:04:33.72" />
                    <SPLIT distance="300" swimtime="00:05:33.61" />
                    <SPLIT distance="350" swimtime="00:06:20.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-18" firstname="Waldemar" gender="M" lastname="Kalbarczyk" nation="POL" athleteid="4245">
              <RESULTS>
                <RESULT eventid="1075" points="458" reactiontime="+74" swimtime="00:02:51.68" resultid="4246" heatid="7950" lane="8" entrytime="00:02:57.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                    <SPLIT distance="100" swimtime="00:01:21.03" />
                    <SPLIT distance="150" swimtime="00:02:13.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="465" reactiontime="+68" swimtime="00:00:33.43" resultid="4247" heatid="7967" lane="8" entrytime="00:00:32.82" />
                <RESULT eventid="1198" points="510" reactiontime="+81" swimtime="00:01:07.96" resultid="4248" heatid="7986" lane="5" entrytime="00:01:07.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="447" reactiontime="+76" swimtime="00:02:57.40" resultid="4249" heatid="8025" lane="6" entrytime="00:02:59.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.55" />
                    <SPLIT distance="100" swimtime="00:01:25.83" />
                    <SPLIT distance="150" swimtime="00:02:12.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="447" reactiontime="+72" swimtime="00:01:22.29" resultid="4250" heatid="8039" lane="4" entrytime="00:01:20.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="425" reactiontime="+89" swimtime="00:05:38.14" resultid="4251" heatid="8154" lane="4" entrytime="00:05:45.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                    <SPLIT distance="100" swimtime="00:01:15.57" />
                    <SPLIT distance="150" swimtime="00:01:57.87" />
                    <SPLIT distance="200" swimtime="00:02:41.40" />
                    <SPLIT distance="250" swimtime="00:03:25.11" />
                    <SPLIT distance="300" swimtime="00:04:10.20" />
                    <SPLIT distance="350" swimtime="00:04:55.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="429" reactiontime="+86" swimtime="00:02:37.00" resultid="4252" heatid="8098" lane="7" entrytime="00:02:38.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                    <SPLIT distance="100" swimtime="00:01:14.22" />
                    <SPLIT distance="150" swimtime="00:01:55.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="378" reactiontime="+88" swimtime="00:06:31.10" resultid="4253" heatid="8164" lane="2" entrytime="00:06:29.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                    <SPLIT distance="100" swimtime="00:01:32.75" />
                    <SPLIT distance="150" swimtime="00:02:22.21" />
                    <SPLIT distance="200" swimtime="00:03:09.65" />
                    <SPLIT distance="250" swimtime="00:04:05.66" />
                    <SPLIT distance="300" swimtime="00:05:02.10" />
                    <SPLIT distance="350" swimtime="00:05:46.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2739" name="MSwim Szczecin">
          <CONTACT city="WOŁCZKOWO" email="m@mswim.pl" name="KACZANOWSKI MIŁOSZ" phone="888 18 1234" street="SŁONECZNA 5" zip="72-003" />
          <ATHLETES>
            <ATHLETE birthdate="1968-05-22" firstname="Miłosz" gender="M" lastname="Kaczanowski" nation="POL" athleteid="2740">
              <RESULTS>
                <RESULT eventid="1105" points="869" reactiontime="+69" swimtime="00:00:28.53" resultid="2741" heatid="7970" lane="6" entrytime="00:00:29.00" />
                <RESULT eventid="1228" points="588" swimtime="00:00:35.68" resultid="2742" heatid="8007" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="1372" points="759" reactiontime="+65" swimtime="00:00:27.58" resultid="2743" heatid="8062" lane="9" entrytime="00:00:28.00" />
                <RESULT eventid="1539" points="711" reactiontime="+72" swimtime="00:00:32.76" resultid="2744" heatid="8116" lane="0" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-11-14" firstname="Anna" gender="F" lastname="Frankowska" nation="POL" athleteid="2749">
              <RESULTS>
                <RESULT eventid="1213" points="483" reactiontime="+102" swimtime="00:00:46.62" resultid="2750" heatid="7996" lane="2" entrytime="00:00:48.00" />
                <RESULT eventid="1387" points="500" reactiontime="+97" swimtime="00:03:35.32" resultid="2751" heatid="8068" lane="8" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.24" />
                    <SPLIT distance="100" swimtime="00:01:43.60" />
                    <SPLIT distance="150" swimtime="00:02:40.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="534" reactiontime="+97" swimtime="00:01:38.74" resultid="2752" heatid="8120" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-10-02" firstname="Jadwiga" gender="F" lastname="Weber" nation="POL" athleteid="2745">
              <RESULTS>
                <RESULT eventid="1273" points="691" reactiontime="+79" swimtime="00:03:17.44" resultid="2746" heatid="8020" lane="9" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.42" />
                    <SPLIT distance="100" swimtime="00:01:34.42" />
                    <SPLIT distance="150" swimtime="00:02:25.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="719" reactiontime="+80" swimtime="00:01:30.23" resultid="2747" heatid="8034" lane="8" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="665" reactiontime="+79" swimtime="00:00:41.72" resultid="2748" heatid="8105" lane="2" entrytime="00:00:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-12" firstname="Zbigniew" gender="M" lastname="Szozda" nation="POL" athleteid="2753">
              <RESULTS>
                <RESULT eventid="1105" points="544" reactiontime="+87" swimtime="00:00:34.93" resultid="2754" heatid="7964" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="1228" points="402" reactiontime="+94" swimtime="00:00:42.05" resultid="2755" heatid="8004" lane="1" entrytime="00:00:41.00" />
                <RESULT eventid="1288" points="606" reactiontime="+78" swimtime="00:03:09.26" resultid="2756" heatid="8025" lane="9" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.38" />
                    <SPLIT distance="100" swimtime="00:01:27.76" />
                    <SPLIT distance="150" swimtime="00:02:18.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" status="DNS" swimtime="00:00:00.00" resultid="2757" heatid="8039" lane="5" entrytime="00:01:23.00" />
                <RESULT eventid="1402" points="528" reactiontime="+97" swimtime="00:03:24.84" resultid="2758" heatid="8073" lane="4" entrytime="00:03:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.84" />
                    <SPLIT distance="100" swimtime="00:01:37.20" />
                    <SPLIT distance="150" swimtime="00:02:30.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="629" reactiontime="+76" swimtime="00:00:37.91" resultid="2759" heatid="8112" lane="3" entrytime="00:00:37.50" />
                <RESULT eventid="1569" points="457" reactiontime="+96" swimtime="00:01:34.57" resultid="2760" heatid="8128" lane="1" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1614" reactiontime="+85" swimtime="00:02:28.20" resultid="2761" heatid="8133" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.66" />
                    <SPLIT distance="100" swimtime="00:01:28.04" />
                    <SPLIT distance="150" swimtime="00:01:56.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2745" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="2740" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="2753" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="03001" nation="POL" region="DOL" clubid="3536" name="MUKP Just Swim Jelenia Góra">
          <CONTACT city="Jelenia Góra" email="marcin.binasiewicz@justswim.pl" name="Binasiewicz Marcin" phone="509071929" state="DOL" zip="58-506" />
          <ATHLETES>
            <ATHLETE birthdate="1987-09-16" firstname="Mariusz" gender="M" lastname="Winogrodzki" nation="POL" athleteid="3544">
              <RESULTS>
                <RESULT eventid="1228" points="893" reactiontime="+78" swimtime="00:00:30.42" resultid="3546" heatid="8010" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1402" points="891" reactiontime="+84" swimtime="00:02:32.11" resultid="3547" heatid="8077" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                    <SPLIT distance="100" swimtime="00:01:13.82" />
                    <SPLIT distance="150" swimtime="00:01:53.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="893" reactiontime="+73" swimtime="00:01:07.14" resultid="3548" heatid="8132" lane="5" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3269" name="niezrzeszony">
          <CONTACT name="Majcher Wiesław" />
          <ATHLETES>
            <ATHLETE birthdate="1950-09-19" firstname="Wiesław" gender="M" lastname="Majcher" nation="POL" athleteid="6017">
              <RESULTS>
                <RESULT eventid="1105" points="154" reactiontime="+86" swimtime="00:00:56.89" resultid="6018" heatid="7962" lane="9" />
                <RESULT eventid="1198" points="295" reactiontime="+116" swimtime="00:01:39.09" resultid="6019" heatid="7980" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="268" reactiontime="+108" swimtime="00:00:56.19" resultid="6020" heatid="8000" lane="9" />
                <RESULT comment="G8 - Ukończenie wyścigu nie w położeniu na plecach" eventid="1342" reactiontime="+75" status="DSQ" swimtime="00:02:12.93" resultid="6021" heatid="8036" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="326" reactiontime="+100" swimtime="00:00:41.80" resultid="6022" heatid="8051" lane="4" />
                <RESULT eventid="1539" points="172" reactiontime="+86" swimtime="00:01:00.16" resultid="6023" heatid="8108" lane="5" />
                <RESULT eventid="1569" points="227" reactiontime="+114" swimtime="00:02:14.85" resultid="6024" heatid="8124" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-04-21" firstname="Iwona" gender="F" lastname="Damljanović-Wacławik" nation="POL" athleteid="3285">
              <RESULTS>
                <RESULT eventid="1090" points="490" reactiontime="+90" swimtime="00:00:38.34" resultid="3286" heatid="7957" lane="2" entrytime="00:00:38.21" />
                <RESULT eventid="1120" points="433" reactiontime="+95" swimtime="00:13:37.49" resultid="3287" heatid="8137" lane="6" entrytime="00:13:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.01" />
                    <SPLIT distance="100" swimtime="00:01:32.50" />
                    <SPLIT distance="150" swimtime="00:02:23.12" />
                    <SPLIT distance="200" swimtime="00:03:14.56" />
                    <SPLIT distance="250" swimtime="00:04:05.72" />
                    <SPLIT distance="300" swimtime="00:04:57.61" />
                    <SPLIT distance="350" swimtime="00:05:49.24" />
                    <SPLIT distance="400" swimtime="00:06:41.75" />
                    <SPLIT distance="450" swimtime="00:07:33.28" />
                    <SPLIT distance="500" swimtime="00:08:25.88" />
                    <SPLIT distance="550" swimtime="00:09:17.87" />
                    <SPLIT distance="600" swimtime="00:10:10.73" />
                    <SPLIT distance="650" swimtime="00:11:02.79" />
                    <SPLIT distance="700" swimtime="00:11:55.30" />
                    <SPLIT distance="750" swimtime="00:12:47.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="457" reactiontime="+89" swimtime="00:01:23.32" resultid="3288" heatid="7975" lane="3" entrytime="00:01:22.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="406" reactiontime="+98" swimtime="00:06:32.90" resultid="3289" heatid="8148" lane="9" entrytime="00:06:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.24" />
                    <SPLIT distance="100" swimtime="00:01:29.86" />
                    <SPLIT distance="150" swimtime="00:02:19.68" />
                    <SPLIT distance="200" swimtime="00:03:10.47" />
                    <SPLIT distance="250" swimtime="00:04:01.38" />
                    <SPLIT distance="300" swimtime="00:04:52.23" />
                    <SPLIT distance="350" swimtime="00:05:43.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="327" reactiontime="+90" swimtime="00:01:43.63" resultid="3290" heatid="8079" lane="0" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="431" reactiontime="+90" swimtime="00:03:02.76" resultid="3291" heatid="8089" lane="2" entrytime="00:03:06.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.96" />
                    <SPLIT distance="100" swimtime="00:01:26.19" />
                    <SPLIT distance="150" swimtime="00:02:14.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-09-27" firstname="Weronika" gender="F" lastname="Kabut" nation="POL" athleteid="3549">
              <RESULTS>
                <RESULT eventid="1181" points="653" reactiontime="+77" swimtime="00:01:07.62" resultid="3550" heatid="7978" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="487" reactiontime="+86" swimtime="00:00:42.70" resultid="3551" heatid="7999" lane="7" entrytime="00:00:39.00" />
                <RESULT eventid="1357" points="635" reactiontime="+78" swimtime="00:00:30.96" resultid="3552" heatid="8050" lane="1" entrytime="00:00:29.00" />
                <RESULT eventid="1387" points="443" reactiontime="+97" swimtime="00:03:27.19" resultid="3553" heatid="8069" lane="1" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.52" />
                    <SPLIT distance="100" swimtime="00:01:39.97" />
                    <SPLIT distance="150" swimtime="00:02:34.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="551" reactiontime="+76" swimtime="00:02:36.31" resultid="3554" heatid="8091" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.97" />
                    <SPLIT distance="100" swimtime="00:01:13.06" />
                    <SPLIT distance="150" swimtime="00:01:55.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="458" reactiontime="+89" swimtime="00:01:36.00" resultid="3555" heatid="8122" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-02" firstname="Janusz" gender="M" lastname="Płonka" nation="POL" athleteid="4365">
              <RESULTS>
                <RESULT eventid="1075" points="173" reactiontime="+112" swimtime="00:04:57.26" resultid="4366" heatid="7945" lane="2" entrytime="00:04:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.20" />
                    <SPLIT distance="100" swimtime="00:02:28.00" />
                    <SPLIT distance="150" swimtime="00:03:56.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="229" reactiontime="+108" swimtime="00:00:49.88" resultid="4367" heatid="7962" lane="6" entrytime="00:00:54.00" />
                <RESULT eventid="1258" points="152" swimtime="00:05:29.74" resultid="4368" heatid="8013" lane="4" entrytime="00:05:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.48" />
                    <SPLIT distance="100" swimtime="00:02:27.52" />
                    <SPLIT distance="150" swimtime="00:04:01.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="180" reactiontime="+84" swimtime="00:04:44.88" resultid="4369" heatid="8023" lane="8" entrytime="00:04:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.63" />
                    <SPLIT distance="100" swimtime="00:02:22.50" />
                    <SPLIT distance="150" swimtime="00:03:39.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="227" reactiontime="+78" swimtime="00:02:00.96" resultid="4370" heatid="8037" lane="7" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="150" reactiontime="+93" swimtime="00:02:17.34" resultid="4371" heatid="8081" lane="5" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="213" reactiontime="+106" swimtime="00:04:11.85" resultid="4372" heatid="8093" lane="4" entrytime="00:04:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.54" />
                    <SPLIT distance="100" swimtime="00:02:03.05" />
                    <SPLIT distance="150" swimtime="00:03:11.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="196" reactiontime="+116" swimtime="00:10:49.08" resultid="4373" heatid="8167" lane="1" entrytime="00:10:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.52" />
                    <SPLIT distance="100" swimtime="00:02:29.68" />
                    <SPLIT distance="150" swimtime="00:04:09.62" />
                    <SPLIT distance="200" swimtime="00:05:33.51" />
                    <SPLIT distance="250" swimtime="00:07:06.24" />
                    <SPLIT distance="300" swimtime="00:08:40.12" />
                    <SPLIT distance="350" swimtime="00:09:45.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-06-07" firstname="Piotr" gender="M" lastname="Orłowski" nation="POL" athleteid="4319">
              <RESULTS>
                <RESULT eventid="1105" points="833" reactiontime="+72" swimtime="00:00:26.83" resultid="4320" heatid="7971" lane="2" entrytime="00:00:28.50" />
                <RESULT eventid="1258" points="743" reactiontime="+73" swimtime="00:02:19.13" resultid="4321" heatid="8017" lane="5" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                    <SPLIT distance="100" swimtime="00:01:05.92" />
                    <SPLIT distance="150" swimtime="00:01:42.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="861" reactiontime="+75" swimtime="00:00:59.34" resultid="4322" heatid="8086" lane="7" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-11-03" firstname="Zenon" gender="M" lastname="Mazur" nation="POL" athleteid="4186">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="4187" heatid="7946" lane="6" entrytime="00:03:55.00" />
                <RESULT eventid="1342" points="478" reactiontime="+79" swimtime="00:01:32.01" resultid="4190" heatid="8038" lane="0" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="377" reactiontime="+92" swimtime="00:03:49.16" resultid="4191" heatid="8072" lane="9" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.79" />
                    <SPLIT distance="100" swimtime="00:01:48.63" />
                    <SPLIT distance="150" swimtime="00:02:48.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="448" reactiontime="+71" swimtime="00:00:42.46" resultid="4192" heatid="8110" lane="5" entrytime="00:00:45.00" />
                <RESULT eventid="1569" points="337" reactiontime="+91" swimtime="00:01:44.68" resultid="4193" heatid="8125" lane="1" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-02-21" firstname="Michał" gender="M" lastname="Karczewski" nation="POL" athleteid="3564">
              <RESULTS>
                <RESULT eventid="1372" points="641" reactiontime="+77" swimtime="00:00:27.29" resultid="3565" heatid="8062" lane="8" entrytime="00:00:27.80" />
                <RESULT eventid="1539" status="DNS" swimtime="00:00:00.00" resultid="3566" heatid="8116" lane="7" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-06-29" firstname="Piotr" gender="M" lastname="Krzekotowski" nation="POL" athleteid="3611">
              <RESULTS>
                <RESULT eventid="1198" points="216" reactiontime="+102" swimtime="00:01:33.04" resultid="3612" heatid="7981" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="204" reactiontime="+106" swimtime="00:00:50.78" resultid="3613" heatid="8001" lane="8" entrytime="00:00:52.00" />
                <RESULT eventid="1372" points="244" reactiontime="+109" swimtime="00:00:40.21" resultid="3614" heatid="8052" lane="3" entrytime="00:00:45.00" />
                <RESULT eventid="1402" points="224" reactiontime="+111" swimtime="00:04:12.93" resultid="3615" heatid="8072" lane="8" entrytime="00:03:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.50" />
                    <SPLIT distance="100" swimtime="00:02:00.97" />
                    <SPLIT distance="150" swimtime="00:03:08.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-07-05" firstname="Sebastian" gender="M" lastname="Figarski" nation="POL" athleteid="3344">
              <RESULTS>
                <RESULT eventid="1288" points="746" reactiontime="+71" swimtime="00:02:25.43" resultid="3345" heatid="8028" lane="3" entrytime="00:02:19.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                    <SPLIT distance="100" swimtime="00:01:08.36" />
                    <SPLIT distance="150" swimtime="00:01:46.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="641" reactiontime="+70" swimtime="00:01:05.56" resultid="3346" heatid="8043" lane="6" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" status="DNS" swimtime="00:00:00.00" resultid="3347" heatid="8117" lane="0" entrytime="00:00:29.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-05-05" firstname="Bogdan" gender="M" lastname="Dubiński" nation="POL" athleteid="3270">
              <RESULTS>
                <RESULT eventid="1075" points="420" reactiontime="+93" swimtime="00:03:36.64" resultid="3271" heatid="7947" lane="8" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.94" />
                    <SPLIT distance="100" swimtime="00:01:48.10" />
                    <SPLIT distance="150" swimtime="00:02:52.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="511" reactiontime="+104" swimtime="00:13:22.68" resultid="3272" heatid="8140" lane="2" entrytime="00:13:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.49" />
                    <SPLIT distance="100" swimtime="00:01:26.55" />
                    <SPLIT distance="150" swimtime="00:02:16.06" />
                    <SPLIT distance="200" swimtime="00:03:06.44" />
                    <SPLIT distance="250" swimtime="00:03:57.21" />
                    <SPLIT distance="300" swimtime="00:04:48.79" />
                    <SPLIT distance="350" swimtime="00:05:40.56" />
                    <SPLIT distance="400" swimtime="00:06:33.03" />
                    <SPLIT distance="450" swimtime="00:07:24.98" />
                    <SPLIT distance="500" swimtime="00:08:17.14" />
                    <SPLIT distance="550" swimtime="00:09:08.55" />
                    <SPLIT distance="600" swimtime="00:09:59.86" />
                    <SPLIT distance="650" swimtime="00:10:51.85" />
                    <SPLIT distance="700" swimtime="00:11:43.36" />
                    <SPLIT distance="750" swimtime="00:12:34.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="344" reactiontime="+102" swimtime="00:04:02.14" resultid="3273" heatid="8015" lane="0" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.69" />
                    <SPLIT distance="100" swimtime="00:02:00.46" />
                    <SPLIT distance="150" swimtime="00:03:05.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="500" reactiontime="+97" swimtime="00:03:33.15" resultid="3274" heatid="8024" lane="1" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.12" />
                    <SPLIT distance="100" swimtime="00:01:44.10" />
                    <SPLIT distance="150" swimtime="00:02:38.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="551" reactiontime="+92" swimtime="00:00:33.32" resultid="3275" heatid="8056" lane="7" entrytime="00:00:32.00" />
                <RESULT eventid="1539" points="549" reactiontime="+83" swimtime="00:00:40.99" resultid="3277" heatid="8111" lane="3" entrytime="00:00:41.00" />
                <RESULT eventid="1599" points="456" reactiontime="+100" swimtime="00:07:38.21" resultid="3278" heatid="8166" lane="6" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.50" />
                    <SPLIT distance="100" swimtime="00:02:00.75" />
                    <SPLIT distance="150" swimtime="00:03:00.12" />
                    <SPLIT distance="200" swimtime="00:03:57.71" />
                    <SPLIT distance="250" swimtime="00:05:05.60" />
                    <SPLIT distance="300" swimtime="00:06:09.81" />
                    <SPLIT distance="350" swimtime="00:06:55.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="542" swimtime="00:06:19.65" resultid="8327" heatid="8325" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.91" />
                    <SPLIT distance="100" swimtime="00:01:26.75" />
                    <SPLIT distance="150" swimtime="00:02:15.83" />
                    <SPLIT distance="200" swimtime="00:03:06.20" />
                    <SPLIT distance="250" swimtime="00:03:56.71" />
                    <SPLIT distance="300" swimtime="00:04:46.95" />
                    <SPLIT distance="350" swimtime="00:05:36.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-02-08" firstname="Kazimierz" gender="M" lastname="Sinicki" nation="POL" athleteid="4475">
              <RESULTS>
                <RESULT eventid="1105" points="653" reactiontime="+88" swimtime="00:00:34.51" resultid="4476" heatid="7966" lane="0" entrytime="00:00:34.50" />
                <RESULT eventid="1198" points="699" reactiontime="+74" swimtime="00:01:08.75" resultid="4477" heatid="7987" lane="9" entrytime="00:01:07.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="725" reactiontime="+82" swimtime="00:00:30.42" resultid="4478" heatid="8058" lane="8" entrytime="00:00:29.75" />
                <RESULT eventid="1509" points="728" reactiontime="+87" swimtime="00:02:37.49" resultid="4479" heatid="8098" lane="6" entrytime="00:02:37.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                    <SPLIT distance="100" swimtime="00:01:18.72" />
                    <SPLIT distance="150" swimtime="00:01:58.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-05-03" firstname="Jakub" gender="M" lastname="Jankowski" nation="POL" athleteid="3514">
              <RESULTS>
                <RESULT eventid="1198" points="527" reactiontime="+112" swimtime="00:01:09.14" resultid="3515" heatid="7988" lane="6" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="566" reactiontime="+115" swimtime="00:00:30.41" resultid="3516" heatid="8059" lane="1" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-07-19" firstname="Wojciech" gender="M" lastname="Wyzga" nation="POL" athleteid="5182">
              <RESULTS>
                <RESULT eventid="1105" points="812" reactiontime="+84" swimtime="00:00:29.18" resultid="5183" heatid="7971" lane="7" entrytime="00:00:28.50" />
                <RESULT eventid="1198" points="656" reactiontime="+62" swimtime="00:01:04.25" resultid="5184" heatid="7991" lane="9" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-06-11" firstname="Marek" gender="M" lastname="Łukaszewicz" nation="POL" athleteid="3788">
              <RESULTS>
                <RESULT eventid="1075" points="560" reactiontime="+90" swimtime="00:03:20.85" resultid="3789" heatid="7946" lane="5" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.69" />
                    <SPLIT distance="100" swimtime="00:01:42.69" />
                    <SPLIT distance="150" swimtime="00:02:39.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="598" reactiontime="+88" swimtime="00:24:52.37" resultid="3790" heatid="8146" lane="4" entrytime="00:35:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.35" />
                    <SPLIT distance="100" swimtime="00:01:33.17" />
                    <SPLIT distance="150" swimtime="00:02:22.18" />
                    <SPLIT distance="200" swimtime="00:03:12.48" />
                    <SPLIT distance="250" swimtime="00:04:02.54" />
                    <SPLIT distance="300" swimtime="00:04:52.45" />
                    <SPLIT distance="350" swimtime="00:05:42.24" />
                    <SPLIT distance="400" swimtime="00:06:33.56" />
                    <SPLIT distance="450" swimtime="00:07:24.72" />
                    <SPLIT distance="500" swimtime="00:08:15.50" />
                    <SPLIT distance="550" swimtime="00:09:05.84" />
                    <SPLIT distance="600" swimtime="00:09:55.25" />
                    <SPLIT distance="650" swimtime="00:10:46.34" />
                    <SPLIT distance="700" swimtime="00:11:35.78" />
                    <SPLIT distance="750" swimtime="00:12:25.54" />
                    <SPLIT distance="800" swimtime="00:13:14.87" />
                    <SPLIT distance="850" swimtime="00:14:05.90" />
                    <SPLIT distance="900" swimtime="00:14:56.16" />
                    <SPLIT distance="950" swimtime="00:15:45.07" />
                    <SPLIT distance="1000" swimtime="00:16:34.75" />
                    <SPLIT distance="1050" swimtime="00:17:25.22" />
                    <SPLIT distance="1100" swimtime="00:18:15.79" />
                    <SPLIT distance="1150" swimtime="00:19:05.37" />
                    <SPLIT distance="1200" swimtime="00:19:56.27" />
                    <SPLIT distance="1250" swimtime="00:20:45.15" />
                    <SPLIT distance="1300" swimtime="00:21:34.75" />
                    <SPLIT distance="1350" swimtime="00:22:25.42" />
                    <SPLIT distance="1400" swimtime="00:23:16.63" />
                    <SPLIT distance="1450" swimtime="00:24:05.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="410" reactiontime="+89" swimtime="00:03:56.87" resultid="3791" heatid="8015" lane="7" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.10" />
                    <SPLIT distance="100" swimtime="00:01:48.12" />
                    <SPLIT distance="150" swimtime="00:02:51.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="614" reactiontime="+95" swimtime="00:06:18.09" resultid="3792" heatid="8155" lane="1" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.69" />
                    <SPLIT distance="100" swimtime="00:01:28.14" />
                    <SPLIT distance="150" swimtime="00:02:15.93" />
                    <SPLIT distance="200" swimtime="00:03:05.49" />
                    <SPLIT distance="250" swimtime="00:03:55.65" />
                    <SPLIT distance="300" swimtime="00:04:45.75" />
                    <SPLIT distance="350" swimtime="00:05:34.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="619" reactiontime="+87" swimtime="00:07:22.76" resultid="3793" heatid="8167" lane="6" entrytime="00:09:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.18" />
                    <SPLIT distance="100" swimtime="00:01:44.58" />
                    <SPLIT distance="150" swimtime="00:02:43.94" />
                    <SPLIT distance="200" swimtime="00:03:43.31" />
                    <SPLIT distance="250" swimtime="00:04:45.50" />
                    <SPLIT distance="300" swimtime="00:05:48.15" />
                    <SPLIT distance="350" swimtime="00:06:36.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-09-27" firstname="Wojciech" gender="M" lastname="Kossowski" nation="POL" athleteid="3567">
              <RESULTS>
                <RESULT eventid="1075" points="490" reactiontime="+129" swimtime="00:03:25.92" resultid="3568" heatid="7948" lane="8" entrytime="00:03:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.07" />
                    <SPLIT distance="100" swimtime="00:01:45.42" />
                    <SPLIT distance="150" swimtime="00:02:40.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="590" reactiontime="+114" swimtime="00:00:40.95" resultid="3569" heatid="8003" lane="7" entrytime="00:00:42.20" />
                <RESULT eventid="1402" points="624" reactiontime="+121" swimtime="00:03:29.33" resultid="3570" heatid="8074" lane="7" entrytime="00:03:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.18" />
                    <SPLIT distance="100" swimtime="00:01:40.26" />
                    <SPLIT distance="150" swimtime="00:02:35.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="645" reactiontime="+121" swimtime="00:01:31.77" resultid="3571" heatid="8128" lane="0" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-05-03" firstname="Joanna" gender="F" lastname="Stępień-Gielo" nation="POL" athleteid="4562">
              <RESULTS>
                <RESULT eventid="1150" points="509" reactiontime="+106" swimtime="00:27:31.45" resultid="4563" heatid="8142" lane="1" entrytime="00:30:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.11" />
                    <SPLIT distance="100" swimtime="00:01:36.56" />
                    <SPLIT distance="150" swimtime="00:02:28.63" />
                    <SPLIT distance="200" swimtime="00:03:22.51" />
                    <SPLIT distance="250" swimtime="00:04:17.08" />
                    <SPLIT distance="300" swimtime="00:05:12.08" />
                    <SPLIT distance="350" swimtime="00:06:07.59" />
                    <SPLIT distance="400" swimtime="00:07:03.66" />
                    <SPLIT distance="450" swimtime="00:07:59.22" />
                    <SPLIT distance="500" swimtime="00:08:54.81" />
                    <SPLIT distance="550" swimtime="00:09:51.00" />
                    <SPLIT distance="600" swimtime="00:10:47.26" />
                    <SPLIT distance="650" swimtime="00:11:43.04" />
                    <SPLIT distance="700" swimtime="00:12:38.77" />
                    <SPLIT distance="750" swimtime="00:13:34.95" />
                    <SPLIT distance="800" swimtime="00:14:31.16" />
                    <SPLIT distance="850" swimtime="00:15:27.24" />
                    <SPLIT distance="900" swimtime="00:16:22.68" />
                    <SPLIT distance="950" swimtime="00:17:19.03" />
                    <SPLIT distance="1000" swimtime="00:18:15.05" />
                    <SPLIT distance="1050" swimtime="00:19:10.54" />
                    <SPLIT distance="1100" swimtime="00:20:06.96" />
                    <SPLIT distance="1150" swimtime="00:21:02.81" />
                    <SPLIT distance="1200" swimtime="00:21:58.79" />
                    <SPLIT distance="1250" swimtime="00:22:55.27" />
                    <SPLIT distance="1300" swimtime="00:23:52.39" />
                    <SPLIT distance="1350" swimtime="00:24:47.63" />
                    <SPLIT distance="1400" swimtime="00:25:44.41" />
                    <SPLIT distance="1450" swimtime="00:26:39.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="624" reactiontime="+83" swimtime="00:00:44.17" resultid="4564" heatid="7997" lane="1" entrytime="00:00:43.52" />
                <RESULT eventid="1273" points="429" reactiontime="+78" swimtime="00:03:41.27" resultid="4565" heatid="8019" lane="8" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.06" />
                    <SPLIT distance="100" swimtime="00:01:47.93" />
                    <SPLIT distance="150" swimtime="00:02:46.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1387" points="582" reactiontime="+86" swimtime="00:03:39.45" resultid="4566" heatid="8068" lane="6" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.17" />
                    <SPLIT distance="100" swimtime="00:01:46.49" />
                    <SPLIT distance="150" swimtime="00:02:42.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="609" reactiontime="+89" swimtime="00:01:38.43" resultid="4567" heatid="8121" lane="1" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-02-06" firstname="Lech" gender="M" lastname="Orecki" nation="POL" athleteid="4315">
              <RESULTS>
                <RESULT eventid="1372" points="495" reactiontime="+87" swimtime="00:00:32.10" resultid="4316" heatid="8060" lane="9" entrytime="00:00:28.75" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-03-07" firstname="Jerzy" gender="M" lastname="Demetraki-Paleolog" nation="POL" athleteid="3517">
              <RESULTS>
                <RESULT eventid="1075" points="346" reactiontime="+111" swimtime="00:03:51.23" resultid="3518" heatid="7948" lane="7" entrytime="00:03:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.41" />
                    <SPLIT distance="100" swimtime="00:01:55.95" />
                    <SPLIT distance="150" swimtime="00:02:59.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="524" reactiontime="+105" swimtime="00:13:16.39" resultid="3519" heatid="8140" lane="7" entrytime="00:13:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.81" />
                    <SPLIT distance="100" swimtime="00:01:32.42" />
                    <SPLIT distance="150" swimtime="00:02:21.50" />
                    <SPLIT distance="200" swimtime="00:03:11.67" />
                    <SPLIT distance="250" swimtime="00:04:00.10" />
                    <SPLIT distance="300" swimtime="00:04:50.11" />
                    <SPLIT distance="350" swimtime="00:05:39.68" />
                    <SPLIT distance="400" swimtime="00:06:29.45" />
                    <SPLIT distance="450" swimtime="00:07:18.98" />
                    <SPLIT distance="500" swimtime="00:08:09.57" />
                    <SPLIT distance="550" swimtime="00:09:00.14" />
                    <SPLIT distance="600" swimtime="00:09:52.23" />
                    <SPLIT distance="650" swimtime="00:10:45.04" />
                    <SPLIT distance="700" swimtime="00:11:35.03" />
                    <SPLIT distance="750" swimtime="00:12:27.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="440" reactiontime="+109" swimtime="00:03:43.14" resultid="3520" heatid="8015" lane="2" entrytime="00:03:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.42" />
                    <SPLIT distance="100" swimtime="00:01:47.69" />
                    <SPLIT distance="150" swimtime="00:02:46.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="551" reactiontime="+106" swimtime="00:06:17.49" resultid="3521" heatid="8154" lane="8" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.76" />
                    <SPLIT distance="100" swimtime="00:01:31.88" />
                    <SPLIT distance="150" swimtime="00:02:21.08" />
                    <SPLIT distance="200" swimtime="00:03:09.97" />
                    <SPLIT distance="250" swimtime="00:03:58.62" />
                    <SPLIT distance="300" swimtime="00:04:45.95" />
                    <SPLIT distance="350" swimtime="00:05:34.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="454" reactiontime="+114" swimtime="00:01:33.13" resultid="3522" heatid="8083" lane="8" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" status="DNS" swimtime="00:00:00.00" resultid="3523" heatid="8097" lane="9" entrytime="00:02:50.00" />
                <RESULT eventid="1599" status="DNS" swimtime="00:00:00.00" resultid="3524" heatid="8166" lane="5" entrytime="00:07:28.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="BLR" clubid="4379" name="niezrzeszony">
          <CONTACT email="yauhenipuzan@gmail.com" name="Puzan Aliaksandr" />
          <ATHLETES>
            <ATHLETE birthdate="1972-01-02" firstname="Aliaksandr" gender="M" lastname="Puzan" nation="BLR" athleteid="4380">
              <RESULTS>
                <RESULT eventid="1105" points="468" reactiontime="+76" swimtime="00:00:33.34" resultid="4381" heatid="7969" lane="3" entrytime="00:00:30.00" />
                <RESULT eventid="1198" points="500" reactiontime="+81" swimtime="00:01:08.43" resultid="4382" heatid="7985" lane="6" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="578" reactiontime="+82" swimtime="00:00:29.50" resultid="4383" heatid="8057" lane="1" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-06-05" firstname="Yauheni" gender="M" lastname="Puzan" nation="BLR" athleteid="4384">
              <RESULTS>
                <RESULT eventid="1105" points="942" reactiontime="+71" swimtime="00:00:25.75" resultid="4385" heatid="7972" lane="3" entrytime="00:00:25.50" />
                <RESULT eventid="1198" points="646" reactiontime="+71" swimtime="00:00:59.80" resultid="4386" heatid="7992" lane="4" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="915" reactiontime="+71" swimtime="00:00:58.14" resultid="4387" heatid="8086" lane="4" entrytime="00:00:57.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3457" name="niezrzeszony Biała Podlaska">
          <CONTACT name="Gromisz Wilhelm" />
          <ATHLETES>
            <ATHLETE birthdate="1981-11-29" firstname="Iga" gender="F" lastname="Olszanowska" nation="POL" athleteid="3469">
              <RESULTS>
                <RESULT eventid="1090" points="721" reactiontime="+85" swimtime="00:00:32.67" resultid="3470" heatid="7960" lane="8" entrytime="00:00:33.00" />
                <RESULT eventid="1243" points="492" reactiontime="+95" swimtime="00:03:05.81" resultid="3471" heatid="8012" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.73" />
                    <SPLIT distance="100" swimtime="00:01:24.27" />
                    <SPLIT distance="150" swimtime="00:02:14.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="618" reactiontime="+84" swimtime="00:01:16.88" resultid="3472" heatid="8080" lane="6" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-03" firstname="Wilhelm" gender="M" lastname="Gromisz" nation="POL" athleteid="3463">
              <RESULTS>
                <RESULT eventid="1105" points="778" reactiontime="+101" swimtime="00:00:27.74" resultid="3464" heatid="7971" lane="6" entrytime="00:00:28.00" />
                <RESULT eventid="1288" points="640" reactiontime="+80" swimtime="00:02:34.94" resultid="3465" heatid="8028" lane="1" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="100" swimtime="00:01:12.55" />
                    <SPLIT distance="150" swimtime="00:01:52.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="751" reactiontime="+74" swimtime="00:01:08.23" resultid="3466" heatid="8043" lane="8" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="781" reactiontime="+101" swimtime="00:01:03.21" resultid="3467" heatid="8086" lane="1" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="842" reactiontime="+74" swimtime="00:00:29.86" resultid="3468" heatid="8117" lane="1" entrytime="00:00:29.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5467" name="Niezrzeszony Białystok">
          <CONTACT email="wzmasters@wp.pl" name="Żmiejko" phone="797309140" />
          <ATHLETES>
            <ATHLETE birthdate="1963-01-01" firstname="Wojciech" gender="M" lastname="Żmiejko" nation="POL" athleteid="5476">
              <RESULTS>
                <RESULT eventid="1075" points="714" reactiontime="+81" swimtime="00:02:41.33" resultid="5477" heatid="7951" lane="3" entrytime="00:02:42.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.03" />
                    <SPLIT distance="100" swimtime="00:01:14.06" />
                    <SPLIT distance="150" swimtime="00:02:02.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="746" reactiontime="+81" swimtime="00:00:30.64" resultid="5478" heatid="7969" lane="1" entrytime="00:00:30.85" />
                <RESULT eventid="1198" points="755" reactiontime="+76" swimtime="00:01:03.34" resultid="5479" heatid="7989" lane="4" entrytime="00:01:02.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="711" reactiontime="+75" swimtime="00:00:28.45" resultid="5480" heatid="8059" lane="3" entrytime="00:00:28.95" />
                <RESULT eventid="1462" points="716" reactiontime="+79" swimtime="00:01:11.17" resultid="5481" heatid="8085" lane="9" entrytime="00:01:11.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="692" reactiontime="+79" swimtime="00:02:26.13" resultid="5482" heatid="8100" lane="8" entrytime="00:02:24.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                    <SPLIT distance="100" swimtime="00:01:09.86" />
                    <SPLIT distance="150" swimtime="00:01:47.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="615" reactiontime="+78" swimtime="00:01:25.23" resultid="5483" heatid="8129" lane="7" entrytime="00:01:25.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="4392" name="niezrzeszony Kołobrzeg">
          <CONTACT name="ROGIŃSKI MARIUSZ" />
          <ATHLETES>
            <ATHLETE birthdate="1971-01-09" firstname="Mariusz" gender="M" lastname="Rogiński" nation="POL" athleteid="4393">
              <RESULTS>
                <RESULT eventid="1105" points="553" reactiontime="+74" swimtime="00:00:31.54" resultid="4394" heatid="7965" lane="6" entrytime="00:00:35.00" />
                <RESULT eventid="1198" points="497" reactiontime="+78" swimtime="00:01:08.56" resultid="4395" heatid="7986" lane="8" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="586" reactiontime="+78" swimtime="00:00:29.36" resultid="4396" heatid="8058" lane="6" entrytime="00:00:29.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAL" nation="POL" region="MAL" clubid="6026" name="Niezrzeszony Kraków">
          <CONTACT email="piotr_urbanczyk@onet.pl" name="URBAŃCZYK PIOTR" phone="608172201" />
          <ATHLETES>
            <ATHLETE birthdate="1984-03-16" firstname="Piotr" gender="M" lastname="Urbańczyk" nation="POL" athleteid="6027">
              <RESULTS>
                <RESULT eventid="1288" points="767" reactiontime="+71" swimtime="00:02:24.07" resultid="6028" heatid="8028" lane="5" entrytime="00:02:18.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                    <SPLIT distance="100" swimtime="00:01:08.27" />
                    <SPLIT distance="150" swimtime="00:01:45.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="690" reactiontime="+71" swimtime="00:01:03.97" resultid="6029" heatid="8043" lane="5" entrytime="00:01:01.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="682" reactiontime="+70" swimtime="00:00:29.56" resultid="6030" heatid="8117" lane="6" entrytime="00:00:28.97" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3794" name="niezrzeszony Nowogard">
          <CONTACT name="Marcel Futoma" />
          <ATHLETES>
            <ATHLETE birthdate="1995-05-18" firstname="Marcel" gender="M" lastname="Futoma" nation="POL" athleteid="3795">
              <RESULTS>
                <RESULT eventid="1198" points="585" reactiontime="+88" swimtime="00:01:01.83" resultid="3796" heatid="7991" lane="0" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="587" reactiontime="+81" swimtime="00:00:27.50" resultid="3797" heatid="8057" lane="7" entrytime="00:00:30.00" />
                <RESULT eventid="1432" points="426" reactiontime="+86" swimtime="00:05:17.43" resultid="3798" heatid="8153" lane="4" entrytime="00:05:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                    <SPLIT distance="100" swimtime="00:01:08.98" />
                    <SPLIT distance="150" swimtime="00:01:48.53" />
                    <SPLIT distance="200" swimtime="00:02:29.69" />
                    <SPLIT distance="250" swimtime="00:03:11.72" />
                    <SPLIT distance="300" swimtime="00:03:54.44" />
                    <SPLIT distance="350" swimtime="00:04:37.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2217" name="Niezrzeszony_AW">
          <CONTACT name="Ryszard Sielski" />
          <ATHLETES>
            <ATHLETE birthdate="1940-11-09" firstname="Alina" gender="F" lastname="Wieczorkiewicz" nation="POL" athleteid="2225">
              <RESULTS>
                <RESULT eventid="1090" points="87" reactiontime="+115" swimtime="00:01:50.30" resultid="2226" heatid="7954" lane="4" entrytime="00:01:55.00" />
                <RESULT eventid="1213" points="83" reactiontime="+126" swimtime="00:01:48.94" resultid="2227" heatid="7994" lane="7" entrytime="00:01:45.00" />
                <RESULT eventid="1273" points="195" reactiontime="+99" swimtime="00:06:54.86" resultid="2228" heatid="8018" lane="2" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:37.38" />
                    <SPLIT distance="100" swimtime="00:03:22.87" />
                    <SPLIT distance="150" swimtime="00:05:10.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="174" reactiontime="+92" swimtime="00:03:14.35" resultid="2229" heatid="8032" lane="6" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:34.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="78" reactiontime="+115" swimtime="00:01:33.08" resultid="2230" heatid="8044" lane="2" entrytime="00:01:25.00" />
                <RESULT eventid="1524" points="150" reactiontime="+89" swimtime="00:01:26.53" resultid="2231" heatid="8103" lane="5" entrytime="00:01:30.00" />
                <RESULT eventid="1554" points="125" reactiontime="+117" swimtime="00:03:48.21" resultid="2232" heatid="8118" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:49.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="3504" name="Niezrzeszony_JK">
          <CONTACT name="JAHNZ KAROLINA" />
          <ATHLETES>
            <ATHLETE birthdate="1984-12-12" firstname="Karolina" gender="F" lastname="Jahnz" nation="POL" athleteid="3505">
              <RESULTS>
                <RESULT eventid="1058" points="451" reactiontime="+72" swimtime="00:03:11.15" resultid="3506" heatid="7943" lane="2" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.42" />
                    <SPLIT distance="100" swimtime="00:01:31.10" />
                    <SPLIT distance="150" swimtime="00:02:27.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="424" reactiontime="+68" swimtime="00:12:42.82" resultid="3507" heatid="8137" lane="3" entrytime="00:13:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.46" />
                    <SPLIT distance="100" swimtime="00:01:25.65" />
                    <SPLIT distance="150" swimtime="00:02:12.82" />
                    <SPLIT distance="200" swimtime="00:03:01.26" />
                    <SPLIT distance="250" swimtime="00:03:50.58" />
                    <SPLIT distance="300" swimtime="00:04:39.48" />
                    <SPLIT distance="350" swimtime="00:05:28.48" />
                    <SPLIT distance="400" swimtime="00:06:17.57" />
                    <SPLIT distance="450" swimtime="00:07:06.10" />
                    <SPLIT distance="500" swimtime="00:07:55.32" />
                    <SPLIT distance="550" swimtime="00:08:43.82" />
                    <SPLIT distance="600" swimtime="00:09:32.75" />
                    <SPLIT distance="650" swimtime="00:10:21.54" />
                    <SPLIT distance="700" swimtime="00:11:09.96" />
                    <SPLIT distance="750" swimtime="00:11:57.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="424" reactiontime="+78" swimtime="00:01:18.42" resultid="3508" heatid="7977" lane="7" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="425" reactiontime="+73" swimtime="00:03:10.76" resultid="3509" heatid="8020" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.44" />
                    <SPLIT distance="100" swimtime="00:01:33.01" />
                    <SPLIT distance="150" swimtime="00:02:22.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="473" reactiontime="+69" swimtime="00:01:28.73" resultid="3510" heatid="8033" lane="6" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1387" points="422" reactiontime="+75" swimtime="00:03:33.76" resultid="3511" heatid="8069" lane="7" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.92" />
                    <SPLIT distance="100" swimtime="00:01:43.50" />
                    <SPLIT distance="150" swimtime="00:02:38.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="419" reactiontime="+64" swimtime="00:02:50.84" resultid="3512" heatid="8091" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                    <SPLIT distance="100" swimtime="00:01:20.09" />
                    <SPLIT distance="150" swimtime="00:02:05.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="384" reactiontime="+78" swimtime="00:01:40.61" resultid="3513" heatid="8121" lane="7" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2123" name="Niezrzeszony_MW">
          <CONTACT name="Wojtakajtis" phone="609481279" />
          <ATHLETES>
            <ATHLETE birthdate="1983-01-12" firstname="Maciej" gender="M" lastname="Wojtakajtis" nation="POL" athleteid="2124">
              <RESULTS>
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="2125" heatid="7993" lane="2" entrytime="00:00:57.00" />
                <RESULT eventid="1372" status="DNS" swimtime="00:00:00.00" resultid="2126" heatid="8065" lane="9" entrytime="00:00:26.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="4721" name="niezrzeszony_NT">
          <CONTACT name="TCHORZEWSKI NORBERT" />
          <ATHLETES>
            <ATHLETE birthdate="1965-03-04" firstname="Norbert" gender="M" lastname="Tchorzewski" nation="POL" athleteid="4722">
              <RESULTS>
                <RESULT eventid="1075" points="470" reactiontime="+87" swimtime="00:03:05.47" resultid="4723" heatid="7949" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.71" />
                    <SPLIT distance="100" swimtime="00:01:23.59" />
                    <SPLIT distance="150" swimtime="00:02:22.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="445" reactiontime="+112" swimtime="00:23:45.37" resultid="4724" heatid="8146" lane="0" entrytime="00:22:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.61" />
                    <SPLIT distance="100" swimtime="00:01:20.27" />
                    <SPLIT distance="150" swimtime="00:02:06.16" />
                    <SPLIT distance="200" swimtime="00:02:53.32" />
                    <SPLIT distance="250" swimtime="00:03:40.68" />
                    <SPLIT distance="300" swimtime="00:04:28.77" />
                    <SPLIT distance="350" swimtime="00:05:16.71" />
                    <SPLIT distance="400" swimtime="00:06:05.45" />
                    <SPLIT distance="450" swimtime="00:06:53.45" />
                    <SPLIT distance="500" swimtime="00:07:42.91" />
                    <SPLIT distance="550" swimtime="00:08:30.82" />
                    <SPLIT distance="600" swimtime="00:09:20.00" />
                    <SPLIT distance="650" swimtime="00:10:08.01" />
                    <SPLIT distance="700" swimtime="00:10:56.11" />
                    <SPLIT distance="750" swimtime="00:11:44.31" />
                    <SPLIT distance="800" swimtime="00:12:33.13" />
                    <SPLIT distance="850" swimtime="00:13:22.10" />
                    <SPLIT distance="900" swimtime="00:14:10.05" />
                    <SPLIT distance="950" swimtime="00:14:57.98" />
                    <SPLIT distance="1000" swimtime="00:15:46.50" />
                    <SPLIT distance="1050" swimtime="00:16:34.68" />
                    <SPLIT distance="1100" swimtime="00:17:23.22" />
                    <SPLIT distance="1150" swimtime="00:18:10.98" />
                    <SPLIT distance="1200" swimtime="00:19:00.64" />
                    <SPLIT distance="1250" swimtime="00:19:48.75" />
                    <SPLIT distance="1300" swimtime="00:20:37.50" />
                    <SPLIT distance="1350" swimtime="00:21:25.42" />
                    <SPLIT distance="1400" swimtime="00:22:14.13" />
                    <SPLIT distance="1450" swimtime="00:23:01.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="590" reactiontime="+83" swimtime="00:01:08.77" resultid="4725" heatid="7987" lane="6" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="383" reactiontime="+102" swimtime="00:03:28.64" resultid="4726" heatid="8015" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.85" />
                    <SPLIT distance="100" swimtime="00:01:29.11" />
                    <SPLIT distance="150" swimtime="00:02:24.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="456" reactiontime="+105" swimtime="00:05:53.97" resultid="4727" heatid="8154" lane="5" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.90" />
                    <SPLIT distance="100" swimtime="00:01:19.02" />
                    <SPLIT distance="150" swimtime="00:02:03.52" />
                    <SPLIT distance="200" swimtime="00:02:49.20" />
                    <SPLIT distance="250" swimtime="00:03:35.50" />
                    <SPLIT distance="300" swimtime="00:04:23.37" />
                    <SPLIT distance="350" swimtime="00:05:10.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="421" reactiontime="+98" swimtime="00:01:24.94" resultid="4728" heatid="8084" lane="2" entrytime="00:01:18.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="550" reactiontime="+103" swimtime="00:02:37.78" resultid="4729" heatid="8098" lane="8" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.63" />
                    <SPLIT distance="100" swimtime="00:01:15.15" />
                    <SPLIT distance="150" swimtime="00:01:57.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="452" reactiontime="+107" swimtime="00:06:54.95" resultid="4730" heatid="8164" lane="8" entrytime="00:06:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.80" />
                    <SPLIT distance="100" swimtime="00:01:35.88" />
                    <SPLIT distance="150" swimtime="00:02:31.91" />
                    <SPLIT distance="200" swimtime="00:03:31.19" />
                    <SPLIT distance="250" swimtime="00:04:31.78" />
                    <SPLIT distance="300" swimtime="00:05:30.85" />
                    <SPLIT distance="350" swimtime="00:06:13.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5320" name="Niezrzeszony_PL">
          <CONTACT name="ZIELEZIŃSKI WŁODZIMIERZ" />
          <ATHLETES>
            <ATHLETE birthdate="1953-04-24" firstname="Włodzimierz" gender="M" lastname="Zielieziński" nation="POL" athleteid="5321">
              <RESULTS>
                <RESULT eventid="1165" points="427" reactiontime="+141" swimtime="00:27:12.62" resultid="5322" heatid="8145" lane="6" entrytime="00:27:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.11" />
                    <SPLIT distance="100" swimtime="00:01:29.68" />
                    <SPLIT distance="150" swimtime="00:02:22.36" />
                    <SPLIT distance="200" swimtime="00:03:15.68" />
                    <SPLIT distance="250" swimtime="00:04:10.92" />
                    <SPLIT distance="300" swimtime="00:05:06.10" />
                    <SPLIT distance="350" swimtime="00:06:01.42" />
                    <SPLIT distance="400" swimtime="00:06:57.13" />
                    <SPLIT distance="450" swimtime="00:07:53.42" />
                    <SPLIT distance="500" swimtime="00:08:48.82" />
                    <SPLIT distance="550" swimtime="00:09:44.75" />
                    <SPLIT distance="600" swimtime="00:10:39.60" />
                    <SPLIT distance="650" swimtime="00:11:35.31" />
                    <SPLIT distance="700" swimtime="00:12:30.33" />
                    <SPLIT distance="750" swimtime="00:13:25.46" />
                    <SPLIT distance="800" swimtime="00:14:20.50" />
                    <SPLIT distance="850" swimtime="00:15:16.16" />
                    <SPLIT distance="900" swimtime="00:16:11.48" />
                    <SPLIT distance="950" swimtime="00:17:07.85" />
                    <SPLIT distance="1000" swimtime="00:18:03.04" />
                    <SPLIT distance="1050" swimtime="00:18:58.11" />
                    <SPLIT distance="1100" swimtime="00:19:53.38" />
                    <SPLIT distance="1150" swimtime="00:20:49.45" />
                    <SPLIT distance="1200" swimtime="00:21:45.36" />
                    <SPLIT distance="1250" swimtime="00:22:41.40" />
                    <SPLIT distance="1300" swimtime="00:23:36.43" />
                    <SPLIT distance="1350" swimtime="00:24:31.11" />
                    <SPLIT distance="1400" swimtime="00:25:25.56" />
                    <SPLIT distance="1450" swimtime="00:26:20.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="5323" heatid="7983" lane="6" entrytime="00:01:20.00" />
                <RESULT eventid="1288" points="491" reactiontime="+88" swimtime="00:03:34.41" resultid="5324" heatid="8024" lane="6" entrytime="00:03:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.42" />
                    <SPLIT distance="100" swimtime="00:01:42.13" />
                    <SPLIT distance="150" swimtime="00:02:39.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="421" reactiontime="+86" swimtime="00:01:39.51" resultid="5325" heatid="8038" lane="5" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" status="DNS" swimtime="00:00:00.00" resultid="5326" heatid="8154" lane="0" entrytime="00:06:15.00" />
                <RESULT eventid="1539" points="549" reactiontime="+75" swimtime="00:00:41.00" resultid="5328" heatid="8111" lane="2" entrytime="00:00:41.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="4374" name="Niezrzeszony_PP">
          <CONTACT name="Poniatowski" />
          <ATHLETES>
            <ATHLETE birthdate="1990-06-15" firstname="Patryk" gender="M" lastname="Poniatowski" nation="POL" athleteid="4375">
              <RESULTS>
                <RESULT eventid="1198" points="819" reactiontime="+74" swimtime="00:00:55.25" resultid="4376" heatid="7993" lane="4" entrytime="00:00:53.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="811" reactiontime="+69" swimtime="00:00:24.82" resultid="4377" heatid="8065" lane="4" entrytime="00:00:23.85" />
                <RESULT eventid="1539" points="813" reactiontime="+70" swimtime="00:00:28.69" resultid="4378" heatid="8117" lane="4" entrytime="00:00:27.90" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="2097" name="Niezrzeszony_ZL">
          <CONTACT name="Lewandowski" />
          <ATHLETES>
            <ATHLETE birthdate="1937-09-19" firstname="Zygmunt" gender="M" lastname="Lewandowski" nation="POL" athleteid="2098">
              <RESULTS>
                <RESULT eventid="1165" points="464" reactiontime="+91" swimtime="00:30:22.64" resultid="2099" heatid="8145" lane="0" entrytime="00:32:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.27" />
                    <SPLIT distance="100" swimtime="00:01:47.36" />
                    <SPLIT distance="150" swimtime="00:02:45.40" />
                    <SPLIT distance="200" swimtime="00:03:45.18" />
                    <SPLIT distance="250" swimtime="00:04:46.08" />
                    <SPLIT distance="300" swimtime="00:05:46.69" />
                    <SPLIT distance="350" swimtime="00:06:46.87" />
                    <SPLIT distance="400" swimtime="00:07:48.01" />
                    <SPLIT distance="450" swimtime="00:08:49.80" />
                    <SPLIT distance="500" swimtime="00:09:51.59" />
                    <SPLIT distance="550" swimtime="00:10:53.72" />
                    <SPLIT distance="600" swimtime="00:11:54.69" />
                    <SPLIT distance="650" swimtime="00:12:56.37" />
                    <SPLIT distance="700" swimtime="00:13:58.37" />
                    <SPLIT distance="750" swimtime="00:14:59.97" />
                    <SPLIT distance="800" swimtime="00:16:01.77" />
                    <SPLIT distance="850" swimtime="00:17:03.36" />
                    <SPLIT distance="900" swimtime="00:18:03.89" />
                    <SPLIT distance="950" swimtime="00:19:05.14" />
                    <SPLIT distance="1000" swimtime="00:20:07.07" />
                    <SPLIT distance="1050" swimtime="00:21:08.27" />
                    <SPLIT distance="1100" swimtime="00:22:09.80" />
                    <SPLIT distance="1150" swimtime="00:23:11.81" />
                    <SPLIT distance="1200" swimtime="00:24:14.70" />
                    <SPLIT distance="1250" swimtime="00:25:17.46" />
                    <SPLIT distance="1300" swimtime="00:26:18.89" />
                    <SPLIT distance="1350" swimtime="00:27:22.25" />
                    <SPLIT distance="1400" swimtime="00:28:24.63" />
                    <SPLIT distance="1450" swimtime="00:29:26.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="465" reactiontime="+105" swimtime="00:01:33.91" resultid="2100" heatid="7982" lane="7" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="433" reactiontime="+100" swimtime="00:00:41.57" resultid="2101" heatid="8053" lane="8" entrytime="00:00:40.00" />
                <RESULT eventid="1432" points="417" reactiontime="+108" swimtime="00:07:40.32" resultid="2102" heatid="8155" lane="0" entrytime="00:07:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.22" />
                    <SPLIT distance="100" swimtime="00:01:46.50" />
                    <SPLIT distance="150" swimtime="00:02:45.31" />
                    <SPLIT distance="200" swimtime="00:03:45.25" />
                    <SPLIT distance="250" swimtime="00:04:44.56" />
                    <SPLIT distance="300" swimtime="00:05:45.33" />
                    <SPLIT distance="350" swimtime="00:06:44.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="409" reactiontime="+103" swimtime="00:03:35.26" resultid="2103" heatid="8094" lane="5" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.51" />
                    <SPLIT distance="100" swimtime="00:01:44.10" />
                    <SPLIT distance="150" swimtime="00:02:40.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="DOL" clubid="4302" name="Niezrzezony">
          <CONTACT email="lorkowska@wp.pl" name="Musialik Marcin" />
          <ATHLETES>
            <ATHLETE birthdate="1994-07-07" firstname="Marcin" gender="M" lastname="Musialik" nation="POL" athleteid="4306">
              <RESULTS>
                <RESULT eventid="1075" points="629" reactiontime="+86" swimtime="00:02:31.25" resultid="4307" heatid="7952" lane="1" entrytime="00:02:38.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.20" />
                    <SPLIT distance="100" swimtime="00:01:10.69" />
                    <SPLIT distance="150" swimtime="00:01:56.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="562" reactiontime="+90" swimtime="00:19:35.77" resultid="4308" heatid="8143" lane="3" entrytime="00:19:30.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                    <SPLIT distance="100" swimtime="00:01:10.00" />
                    <SPLIT distance="150" swimtime="00:01:47.68" />
                    <SPLIT distance="200" swimtime="00:02:26.21" />
                    <SPLIT distance="250" swimtime="00:03:05.00" />
                    <SPLIT distance="300" swimtime="00:03:44.15" />
                    <SPLIT distance="350" swimtime="00:04:23.13" />
                    <SPLIT distance="400" swimtime="00:05:02.35" />
                    <SPLIT distance="450" swimtime="00:05:41.54" />
                    <SPLIT distance="500" swimtime="00:06:21.40" />
                    <SPLIT distance="550" swimtime="00:07:00.79" />
                    <SPLIT distance="600" swimtime="00:07:40.66" />
                    <SPLIT distance="650" swimtime="00:08:20.26" />
                    <SPLIT distance="700" swimtime="00:09:00.10" />
                    <SPLIT distance="750" swimtime="00:09:39.65" />
                    <SPLIT distance="800" swimtime="00:10:19.30" />
                    <SPLIT distance="850" swimtime="00:10:58.79" />
                    <SPLIT distance="900" swimtime="00:11:38.67" />
                    <SPLIT distance="950" swimtime="00:12:18.42" />
                    <SPLIT distance="1000" swimtime="00:12:58.35" />
                    <SPLIT distance="1050" swimtime="00:13:38.21" />
                    <SPLIT distance="1100" swimtime="00:14:17.83" />
                    <SPLIT distance="1150" swimtime="00:14:57.60" />
                    <SPLIT distance="1200" swimtime="00:15:37.62" />
                    <SPLIT distance="1250" swimtime="00:16:17.51" />
                    <SPLIT distance="1300" swimtime="00:16:57.47" />
                    <SPLIT distance="1350" swimtime="00:17:37.30" />
                    <SPLIT distance="1400" swimtime="00:18:17.06" />
                    <SPLIT distance="1450" swimtime="00:18:56.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="562" reactiontime="+85" swimtime="00:02:32.70" resultid="4309" heatid="8017" lane="9" entrytime="00:02:45.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.17" />
                    <SPLIT distance="100" swimtime="00:01:13.30" />
                    <SPLIT distance="150" swimtime="00:01:53.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="604" reactiontime="+74" swimtime="00:02:30.28" resultid="4310" heatid="8027" lane="1" entrytime="00:02:44.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.31" />
                    <SPLIT distance="100" swimtime="00:01:14.68" />
                    <SPLIT distance="150" swimtime="00:01:52.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="533" reactiontime="+71" swimtime="00:01:11.95" resultid="4311" heatid="8041" lane="1" entrytime="00:01:15.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="612" reactiontime="+82" swimtime="00:04:41.25" resultid="4312" heatid="8151" lane="2" entrytime="00:04:45.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                    <SPLIT distance="100" swimtime="00:01:06.38" />
                    <SPLIT distance="150" swimtime="00:01:41.98" />
                    <SPLIT distance="200" swimtime="00:02:18.23" />
                    <SPLIT distance="250" swimtime="00:02:54.19" />
                    <SPLIT distance="300" swimtime="00:03:30.73" />
                    <SPLIT distance="350" swimtime="00:04:06.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="654" reactiontime="+86" swimtime="00:02:13.17" resultid="4313" heatid="8100" lane="4" entrytime="00:02:20.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.97" />
                    <SPLIT distance="100" swimtime="00:01:04.55" />
                    <SPLIT distance="150" swimtime="00:01:39.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="661" reactiontime="+89" swimtime="00:05:21.19" resultid="4314" heatid="8162" lane="8" entrytime="00:05:39.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                    <SPLIT distance="100" swimtime="00:01:13.37" />
                    <SPLIT distance="150" swimtime="00:01:54.08" />
                    <SPLIT distance="200" swimtime="00:02:34.38" />
                    <SPLIT distance="250" swimtime="00:03:21.86" />
                    <SPLIT distance="300" swimtime="00:04:10.12" />
                    <SPLIT distance="350" swimtime="00:04:46.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ORS OPOLE" nation="POL" region="OPO" clubid="4323" name="ORS Opole">
          <CONTACT email="wkania62@gmail.com" name="Kania" />
          <ATHLETES>
            <ATHLETE birthdate="1962-01-01" firstname="Waldemar" gender="M" lastname="Kania" nation="POL" athleteid="4333">
              <RESULTS>
                <RESULT eventid="1165" points="467" reactiontime="+104" swimtime="00:23:22.80" resultid="4334" heatid="8144" lane="6" entrytime="00:22:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.42" />
                    <SPLIT distance="100" swimtime="00:01:25.90" />
                    <SPLIT distance="150" swimtime="00:02:12.00" />
                    <SPLIT distance="200" swimtime="00:02:58.56" />
                    <SPLIT distance="250" swimtime="00:03:44.83" />
                    <SPLIT distance="300" swimtime="00:04:30.55" />
                    <SPLIT distance="350" swimtime="00:05:17.33" />
                    <SPLIT distance="400" swimtime="00:06:03.68" />
                    <SPLIT distance="450" swimtime="00:06:50.15" />
                    <SPLIT distance="500" swimtime="00:07:36.73" />
                    <SPLIT distance="550" swimtime="00:08:23.83" />
                    <SPLIT distance="600" swimtime="00:09:11.01" />
                    <SPLIT distance="650" swimtime="00:09:58.10" />
                    <SPLIT distance="700" swimtime="00:10:45.28" />
                    <SPLIT distance="750" swimtime="00:11:32.58" />
                    <SPLIT distance="800" swimtime="00:12:19.58" />
                    <SPLIT distance="850" swimtime="00:13:07.07" />
                    <SPLIT distance="900" swimtime="00:13:54.67" />
                    <SPLIT distance="950" swimtime="00:14:42.22" />
                    <SPLIT distance="1000" swimtime="00:15:29.90" />
                    <SPLIT distance="1050" swimtime="00:16:17.70" />
                    <SPLIT distance="1100" swimtime="00:17:05.29" />
                    <SPLIT distance="1150" swimtime="00:17:53.17" />
                    <SPLIT distance="1200" swimtime="00:18:41.01" />
                    <SPLIT distance="1250" swimtime="00:19:28.97" />
                    <SPLIT distance="1300" swimtime="00:20:16.22" />
                    <SPLIT distance="1350" swimtime="00:21:03.55" />
                    <SPLIT distance="1400" swimtime="00:21:50.54" />
                    <SPLIT distance="1450" swimtime="00:22:37.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="4335" heatid="8024" lane="2" entrytime="00:03:30.00" />
                <RESULT eventid="1509" status="DNS" swimtime="00:00:00.00" resultid="4337" heatid="8097" lane="4" entrytime="00:02:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-01" firstname="Agnieszka" gender="F" lastname="Bartnikowska" nation="POL" athleteid="4324">
              <RESULTS>
                <RESULT eventid="1058" points="618" reactiontime="+89" swimtime="00:02:50.58" resultid="4325" heatid="7944" lane="7" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                    <SPLIT distance="100" swimtime="00:01:18.98" />
                    <SPLIT distance="150" swimtime="00:02:09.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="601" reactiontime="+90" swimtime="00:00:33.53" resultid="4326" heatid="7959" lane="7" entrytime="00:00:35.00" />
                <RESULT eventid="1181" status="DNS" swimtime="00:00:00.00" resultid="4327" heatid="7978" lane="6" entrytime="00:01:10.00" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="4328" heatid="8020" lane="3" entrytime="00:02:55.00" />
                <RESULT eventid="1326" status="DNS" swimtime="00:00:00.00" resultid="4329" heatid="8035" lane="9" entrytime="00:01:20.00" />
                <RESULT eventid="1447" status="DNS" swimtime="00:00:00.00" resultid="4330" heatid="8080" lane="0" entrytime="00:01:20.00" />
                <RESULT eventid="1493" status="DNS" swimtime="00:00:00.00" resultid="4331" heatid="8091" lane="2" entrytime="00:02:36.00" />
                <RESULT eventid="1584" status="DNS" swimtime="00:00:00.00" resultid="4332" heatid="8160" lane="4" entrytime="00:06:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="SVK" clubid="6031" name="PSK Žilina, Słowacja">
          <CONTACT name="Ratislav Pavlik" />
          <ATHLETES>
            <ATHLETE birthdate="1960-01-01" firstname="Ratislav" gender="M" lastname="Pavlik" nation="SVK" athleteid="6032">
              <RESULTS>
                <RESULT eventid="1228" points="761" reactiontime="+84" swimtime="00:00:34.00" resultid="6033" heatid="8008" lane="7" entrytime="00:00:34.50" />
                <RESULT eventid="1342" points="1107" reactiontime="+71" swimtime="00:01:09.59" resultid="6034" heatid="8042" lane="5" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="1009" reactiontime="+70" swimtime="00:00:32.39" resultid="6035" heatid="8115" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1569" points="788" reactiontime="+84" swimtime="00:01:18.85" resultid="6036" heatid="8131" lane="7" entrytime="00:01:16.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="RMKS RYBNI" nation="POL" region="SLA" clubid="3964" name="RMKS Rybnik">
          <CONTACT city="Rybnik" email="aniaduda0511@tlen.pl" internet="http://www.rmks.rybnik.pl/" name="Tymusz Rafał" phone="601861688" state="SLA" street="powstancow slaskich 40/42" zip="44-200" />
          <ATHLETES>
            <ATHLETE birthdate="1990-02-28" firstname="Monika" gender="F" lastname="Nowak" nation="POL" athleteid="3977">
              <RESULTS>
                <RESULT eventid="1090" points="495" reactiontime="+72" swimtime="00:00:35.76" resultid="3978" heatid="7958" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="1213" points="480" reactiontime="+77" swimtime="00:00:41.70" resultid="3979" heatid="7997" lane="4" entrytime="00:00:42.00" />
                <RESULT eventid="1447" points="471" reactiontime="+84" swimtime="00:01:22.42" resultid="3980" heatid="8080" lane="1" entrytime="00:01:16.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1584" points="457" reactiontime="+81" swimtime="00:06:44.53" resultid="3981" heatid="8160" lane="5" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                    <SPLIT distance="100" swimtime="00:01:25.75" />
                    <SPLIT distance="150" swimtime="00:02:25.09" />
                    <SPLIT distance="200" swimtime="00:03:20.90" />
                    <SPLIT distance="250" swimtime="00:04:15.38" />
                    <SPLIT distance="300" swimtime="00:05:10.54" />
                    <SPLIT distance="350" swimtime="00:05:59.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-11-07" firstname="Iwona" gender="F" lastname="Cymerman" nation="POL" athleteid="3972">
              <RESULTS>
                <RESULT eventid="1090" points="708" reactiontime="+65" swimtime="00:00:32.86" resultid="3973" heatid="7959" lane="6" entrytime="00:00:34.50" />
                <RESULT eventid="1213" points="510" reactiontime="+78" swimtime="00:00:40.87" resultid="3974" heatid="7999" lane="1" entrytime="00:00:39.00" />
                <RESULT eventid="1387" points="525" reactiontime="+73" swimtime="00:03:18.80" resultid="3975" heatid="8069" lane="3" entrytime="00:03:20.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.67" />
                    <SPLIT distance="100" swimtime="00:01:35.49" />
                    <SPLIT distance="150" swimtime="00:02:27.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="562" reactiontime="+74" swimtime="00:01:28.60" resultid="3976" heatid="8123" lane="2" entrytime="00:01:26.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-15" firstname="Anna" gender="F" lastname="Duda" nation="POL" athleteid="3965">
              <RESULTS>
                <RESULT eventid="1090" points="898" reactiontime="+67" swimtime="00:00:30.36" resultid="3966" heatid="7960" lane="5" entrytime="00:00:30.40" />
                <RESULT eventid="1181" points="708" reactiontime="+80" swimtime="00:01:06.14" resultid="3967" heatid="7978" lane="4" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.25" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1243" points="633" reactiontime="+85" swimtime="00:02:50.88" resultid="3968" heatid="8012" lane="3" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                    <SPLIT distance="100" swimtime="00:01:16.00" />
                    <SPLIT distance="150" swimtime="00:02:02.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="777" reactiontime="+78" swimtime="00:00:29.53" resultid="3969" heatid="8049" lane="5" entrytime="00:00:29.50" />
                <RESULT eventid="1447" points="777" reactiontime="+83" swimtime="00:01:11.22" resultid="3970" heatid="8080" lane="5" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1584" points="640" reactiontime="+91" swimtime="00:05:59.65" resultid="3971" heatid="8159" lane="8" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                    <SPLIT distance="100" swimtime="00:01:15.41" />
                    <SPLIT distance="150" swimtime="00:02:06.32" />
                    <SPLIT distance="200" swimtime="00:02:54.36" />
                    <SPLIT distance="250" swimtime="00:03:48.25" />
                    <SPLIT distance="300" swimtime="00:04:41.50" />
                    <SPLIT distance="350" swimtime="00:05:21.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-03" firstname="Agnieszka" gender="F" lastname="Bieniak" nation="POL" athleteid="3982">
              <RESULTS>
                <RESULT eventid="1058" points="601" reactiontime="+82" swimtime="00:02:52.17" resultid="3983" heatid="7944" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                    <SPLIT distance="100" swimtime="00:01:18.31" />
                    <SPLIT distance="150" swimtime="00:02:09.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="603" reactiontime="+80" swimtime="00:00:33.48" resultid="3984" heatid="7959" lane="4" entrytime="00:00:34.00" />
                <RESULT eventid="1213" points="574" swimtime="00:00:39.28" resultid="3985" heatid="7998" lane="0" entrytime="00:00:42.00" />
                <RESULT eventid="1326" points="662" swimtime="00:01:17.76" resultid="3986" heatid="8035" lane="8" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="703" reactiontime="+83" swimtime="00:00:30.41" resultid="3987" heatid="8048" lane="5" entrytime="00:00:32.00" />
                <RESULT eventid="1524" points="650" reactiontime="+73" swimtime="00:00:35.89" resultid="3988" heatid="8107" lane="1" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1303" reactiontime="+73" swimtime="00:04:35.45" resultid="3989" heatid="8029" lane="6" entrytime="00:04:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.83" />
                    <SPLIT distance="100" swimtime="00:01:08.44" />
                    <SPLIT distance="150" swimtime="00:01:43.68" />
                    <SPLIT distance="200" swimtime="00:02:23.17" />
                    <SPLIT distance="250" swimtime="00:02:54.07" />
                    <SPLIT distance="300" swimtime="00:03:30.24" />
                    <SPLIT distance="350" swimtime="00:04:00.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3972" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="3977" number="2" reactiontime="+75" />
                    <RELAYPOSITION athleteid="3982" number="3" reactiontime="+67" />
                    <RELAYPOSITION athleteid="3965" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="4397" name="Rydultowska.AAS 60+">
          <CONTACT city="wodzisla sl`" email="otelom.080966@interia.pl" name="otlik marian" phone="692112775" street="wodzisla sl" zip="44-300" />
          <ATHLETES>
            <ATHLETE birthdate="1953-11-24" firstname="Jerzy" gender="M" lastname="Ciecior" nation="POL" athleteid="4407">
              <RESULTS>
                <RESULT eventid="1075" points="531" reactiontime="+96" swimtime="00:03:20.41" resultid="4408" heatid="7948" lane="6" entrytime="00:03:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.70" />
                    <SPLIT distance="100" swimtime="00:01:31.76" />
                    <SPLIT distance="150" swimtime="00:02:35.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="528" swimtime="00:25:20.87" resultid="4409" heatid="8144" lane="9" entrytime="00:24:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.10" />
                    <SPLIT distance="100" swimtime="00:01:31.21" />
                    <SPLIT distance="150" swimtime="00:02:20.83" />
                    <SPLIT distance="200" swimtime="00:03:11.68" />
                    <SPLIT distance="250" swimtime="00:04:02.74" />
                    <SPLIT distance="300" swimtime="00:04:53.77" />
                    <SPLIT distance="350" swimtime="00:05:44.56" />
                    <SPLIT distance="400" swimtime="00:06:35.43" />
                    <SPLIT distance="450" swimtime="00:07:26.35" />
                    <SPLIT distance="500" swimtime="00:08:17.60" />
                    <SPLIT distance="550" swimtime="00:09:08.40" />
                    <SPLIT distance="600" swimtime="00:10:00.19" />
                    <SPLIT distance="650" swimtime="00:10:51.32" />
                    <SPLIT distance="700" swimtime="00:11:43.00" />
                    <SPLIT distance="750" swimtime="00:12:34.35" />
                    <SPLIT distance="800" swimtime="00:13:25.02" />
                    <SPLIT distance="850" swimtime="00:14:16.40" />
                    <SPLIT distance="900" swimtime="00:15:07.66" />
                    <SPLIT distance="950" swimtime="00:15:59.06" />
                    <SPLIT distance="1000" swimtime="00:16:50.98" />
                    <SPLIT distance="1050" swimtime="00:17:42.41" />
                    <SPLIT distance="1100" swimtime="00:18:33.61" />
                    <SPLIT distance="1150" swimtime="00:19:25.39" />
                    <SPLIT distance="1200" swimtime="00:20:16.85" />
                    <SPLIT distance="1250" swimtime="00:21:08.34" />
                    <SPLIT distance="1300" swimtime="00:22:00.40" />
                    <SPLIT distance="1350" swimtime="00:22:51.98" />
                    <SPLIT distance="1400" swimtime="00:23:43.10" />
                    <SPLIT distance="1450" swimtime="00:24:32.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="538" reactiontime="+81" swimtime="00:03:28.03" resultid="4410" heatid="8028" lane="4" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.66" />
                    <SPLIT distance="100" swimtime="00:01:40.02" />
                    <SPLIT distance="150" swimtime="00:02:34.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="477" reactiontime="+85" swimtime="00:01:35.51" resultid="4411" heatid="8039" lane="1" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="469" reactiontime="+89" swimtime="00:01:32.13" resultid="4412" heatid="8083" lane="2" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="516" reactiontime="+76" swimtime="00:00:41.86" resultid="4413" heatid="8112" lane="0" entrytime="00:00:40.00" />
                <RESULT eventid="1599" points="487" reactiontime="+97" swimtime="00:07:28.35" resultid="4414" heatid="8165" lane="1" entrytime="00:07:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.86" />
                    <SPLIT distance="100" swimtime="00:01:43.61" />
                    <SPLIT distance="150" swimtime="00:02:43.00" />
                    <SPLIT distance="200" swimtime="00:03:41.28" />
                    <SPLIT distance="250" swimtime="00:04:47.32" />
                    <SPLIT distance="300" swimtime="00:05:52.39" />
                    <SPLIT distance="350" swimtime="00:06:40.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-05-16" firstname="Rudolf" gender="M" lastname="Bugla" nation="POL" athleteid="4424">
              <RESULTS>
                <RESULT eventid="1075" points="348" reactiontime="+119" swimtime="00:04:26.06" resultid="4425" heatid="7945" lane="6" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.58" />
                    <SPLIT distance="100" swimtime="00:02:08.95" />
                    <SPLIT distance="150" swimtime="00:03:23.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="256" reactiontime="+102" swimtime="00:00:57.78" resultid="4426" heatid="7962" lane="7" entrytime="00:01:02.00" />
                <RESULT eventid="1228" points="339" reactiontime="+96" swimtime="00:00:56.75" resultid="4427" heatid="8000" lane="3" entrytime="00:01:01.00" />
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1258" points="317" reactiontime="+98" swimtime="00:05:10.52" resultid="4428" heatid="8014" lane="7" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.10" />
                    <SPLIT distance="100" swimtime="00:02:29.63" />
                    <SPLIT distance="150" swimtime="00:03:52.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="373" reactiontime="+99" swimtime="00:04:43.30" resultid="4429" heatid="8071" lane="3" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.56" />
                    <SPLIT distance="100" swimtime="00:02:17.72" />
                    <SPLIT distance="150" swimtime="00:03:31.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="256" reactiontime="+99" swimtime="00:02:19.56" resultid="4430" heatid="8081" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="335" reactiontime="+88" swimtime="00:02:09.39" resultid="4431" heatid="8125" lane="7" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="378" reactiontime="+88" swimtime="00:10:05.62" resultid="4432" heatid="8167" lane="2" entrytime="00:09:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.91" />
                    <SPLIT distance="100" swimtime="00:02:32.46" />
                    <SPLIT distance="150" swimtime="00:03:49.78" />
                    <SPLIT distance="200" swimtime="00:05:06.69" />
                    <SPLIT distance="250" swimtime="00:06:28.29" />
                    <SPLIT distance="300" swimtime="00:07:48.63" />
                    <SPLIT distance="350" swimtime="00:08:56.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-09-07" firstname="Leon" gender="M" lastname="Irczyk" nation="POL" athleteid="4398">
              <RESULTS>
                <RESULT eventid="1075" points="260" reactiontime="+134" swimtime="00:04:14.31" resultid="4399" heatid="7946" lane="3" entrytime="00:03:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.24" />
                    <SPLIT distance="100" swimtime="00:02:20.22" />
                    <SPLIT distance="150" swimtime="00:03:16.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="318" swimtime="00:15:40.44" resultid="4400" heatid="8141" lane="4" entrytime="00:15:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.66" />
                    <SPLIT distance="100" swimtime="00:01:49.23" />
                    <SPLIT distance="150" swimtime="00:02:49.37" />
                    <SPLIT distance="200" swimtime="00:03:48.77" />
                    <SPLIT distance="250" swimtime="00:04:48.29" />
                    <SPLIT distance="300" swimtime="00:05:48.29" />
                    <SPLIT distance="350" swimtime="00:06:48.39" />
                    <SPLIT distance="400" swimtime="00:07:48.10" />
                    <SPLIT distance="450" swimtime="00:08:47.84" />
                    <SPLIT distance="500" swimtime="00:09:46.93" />
                    <SPLIT distance="550" swimtime="00:10:46.25" />
                    <SPLIT distance="600" swimtime="00:11:45.80" />
                    <SPLIT distance="650" swimtime="00:12:45.07" />
                    <SPLIT distance="700" swimtime="00:13:43.64" />
                    <SPLIT distance="750" swimtime="00:14:42.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="349" reactiontime="+106" swimtime="00:00:48.75" resultid="4401" heatid="8001" lane="5" entrytime="00:00:48.47" />
                <RESULT eventid="1258" points="224" reactiontime="+122" swimtime="00:04:39.49" resultid="4402" heatid="8014" lane="3" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.18" />
                    <SPLIT distance="100" swimtime="00:02:16.71" />
                    <SPLIT distance="150" swimtime="00:03:28.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="502" reactiontime="+121" swimtime="00:03:45.12" resultid="4403" heatid="8072" lane="4" entrytime="00:03:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.89" />
                    <SPLIT distance="100" swimtime="00:01:49.47" />
                    <SPLIT distance="150" swimtime="00:02:48.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="313" reactiontime="+112" swimtime="00:07:35.71" resultid="4404" heatid="8155" lane="8" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.66" />
                    <SPLIT distance="100" swimtime="00:01:51.50" />
                    <SPLIT distance="150" swimtime="00:02:50.13" />
                    <SPLIT distance="200" swimtime="00:03:49.62" />
                    <SPLIT distance="250" swimtime="00:04:48.91" />
                    <SPLIT distance="300" swimtime="00:05:46.52" />
                    <SPLIT distance="350" swimtime="00:06:43.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="418" reactiontime="+110" swimtime="00:01:46.01" resultid="4405" heatid="8126" lane="3" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="277" reactiontime="+108" swimtime="00:09:00.60" resultid="4406" heatid="8166" lane="0" entrytime="00:08:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.55" />
                    <SPLIT distance="100" swimtime="00:02:08.97" />
                    <SPLIT distance="150" swimtime="00:03:31.41" />
                    <SPLIT distance="200" swimtime="00:04:53.66" />
                    <SPLIT distance="250" swimtime="00:05:57.11" />
                    <SPLIT distance="300" swimtime="00:07:00.36" />
                    <SPLIT distance="350" swimtime="00:08:01.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-09-08" firstname="Marian" gender="M" lastname="Otlik" nation="POL" athleteid="4415">
              <RESULTS>
                <RESULT eventid="1075" points="435" reactiontime="+71" swimtime="00:03:12.43" resultid="4416" heatid="7948" lane="3" entrytime="00:03:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                    <SPLIT distance="100" swimtime="00:01:31.64" />
                    <SPLIT distance="150" swimtime="00:02:29.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="412" reactiontime="+65" swimtime="00:00:36.57" resultid="4417" heatid="7965" lane="5" entrytime="00:00:35.00" />
                <RESULT eventid="1198" points="529" reactiontime="+60" swimtime="00:01:09.04" resultid="4418" heatid="7985" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="286" reactiontime="+68" swimtime="00:00:45.33" resultid="4419" heatid="8002" lane="3" entrytime="00:00:45.00" />
                <RESULT eventid="1372" points="584" reactiontime="+61" swimtime="00:00:30.09" resultid="4420" heatid="8057" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="1432" points="328" reactiontime="+75" swimtime="00:06:11.18" resultid="4421" heatid="8154" lane="3" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.40" />
                    <SPLIT distance="100" swimtime="00:01:22.32" />
                    <SPLIT distance="150" swimtime="00:02:08.74" />
                    <SPLIT distance="200" swimtime="00:02:57.80" />
                    <SPLIT distance="250" swimtime="00:03:47.18" />
                    <SPLIT distance="300" swimtime="00:04:36.25" />
                    <SPLIT distance="350" swimtime="00:05:25.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="365" reactiontime="+68" swimtime="00:02:46.91" resultid="4422" heatid="8097" lane="7" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                    <SPLIT distance="100" swimtime="00:01:17.22" />
                    <SPLIT distance="150" swimtime="00:02:02.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="367" reactiontime="+82" swimtime="00:07:16.11" resultid="4423" heatid="8165" lane="7" entrytime="00:07:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.56" />
                    <SPLIT distance="100" swimtime="00:01:37.28" />
                    <SPLIT distance="150" swimtime="00:02:37.02" />
                    <SPLIT distance="200" swimtime="00:03:36.37" />
                    <SPLIT distance="250" swimtime="00:04:37.65" />
                    <SPLIT distance="300" swimtime="00:05:40.27" />
                    <SPLIT distance="350" swimtime="00:06:30.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="4443" name="Sikret Gliwice">
          <CONTACT city="GLIWICE" email="joannaeco@tlen.pl" name="JOANNA ZAGAŁA" phone="601427257" state="ŚL" street="JAGIELOŃSKA 21" zip="44-100" />
          <ATHLETES>
            <ATHLETE birthdate="1959-06-24" firstname="Joanna" gender="F" lastname="Zagała" nation="POL" athleteid="4452">
              <RESULTS>
                <RESULT eventid="1058" points="408" reactiontime="+76" swimtime="00:03:54.08" resultid="4453" heatid="7941" lane="4" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.16" />
                    <SPLIT distance="100" swimtime="00:01:54.38" />
                    <SPLIT distance="150" swimtime="00:02:58.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="499" reactiontime="+72" swimtime="00:14:57.69" resultid="4454" heatid="8137" lane="9" entrytime="00:15:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.74" />
                    <SPLIT distance="100" swimtime="00:01:44.67" />
                    <SPLIT distance="150" swimtime="00:02:41.97" />
                    <SPLIT distance="200" swimtime="00:03:39.11" />
                    <SPLIT distance="250" swimtime="00:04:36.58" />
                    <SPLIT distance="300" swimtime="00:05:34.36" />
                    <SPLIT distance="350" swimtime="00:06:32.24" />
                    <SPLIT distance="400" swimtime="00:07:30.96" />
                    <SPLIT distance="450" swimtime="00:08:28.01" />
                    <SPLIT distance="500" swimtime="00:09:25.26" />
                    <SPLIT distance="550" swimtime="00:10:21.73" />
                    <SPLIT distance="600" swimtime="00:11:18.29" />
                    <SPLIT distance="650" swimtime="00:12:15.67" />
                    <SPLIT distance="700" swimtime="00:13:11.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="415" reactiontime="+75" swimtime="00:00:51.37" resultid="4455" heatid="7995" lane="1" entrytime="00:01:00.00" />
                <RESULT eventid="1273" points="426" reactiontime="+87" swimtime="00:03:51.85" resultid="4456" heatid="8018" lane="4" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.53" />
                    <SPLIT distance="100" swimtime="00:01:58.39" />
                    <SPLIT distance="150" swimtime="00:02:58.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="505" reactiontime="+77" swimtime="00:00:38.77" resultid="4457" heatid="8044" lane="3" entrytime="00:01:00.00" />
                <RESULT eventid="1387" points="462" reactiontime="+77" swimtime="00:04:08.34" resultid="4458" heatid="8067" lane="1" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.45" />
                    <SPLIT distance="100" swimtime="00:02:01.07" />
                    <SPLIT distance="150" swimtime="00:03:05.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="483" reactiontime="+73" swimtime="00:03:19.89" resultid="4459" heatid="8087" lane="5" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.19" />
                    <SPLIT distance="100" swimtime="00:01:40.17" />
                    <SPLIT distance="150" swimtime="00:02:32.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="413" reactiontime="+75" swimtime="00:01:54.69" resultid="4460" heatid="8119" lane="6" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-02-05" firstname="Zofia" gender="F" lastname="Dąbrowska" nation="POL" athleteid="4444">
              <RESULTS>
                <RESULT eventid="1090" points="263" reactiontime="+72" swimtime="00:00:53.99" resultid="4445" heatid="7955" lane="6" entrytime="00:00:52.00" />
                <RESULT eventid="1213" points="395" reactiontime="+77" swimtime="00:00:52.24" resultid="4446" heatid="7995" lane="4" entrytime="00:00:51.00" />
                <RESULT eventid="1243" points="315" reactiontime="+89" swimtime="00:04:45.62" resultid="4447" heatid="8011" lane="5" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.87" />
                    <SPLIT distance="100" swimtime="00:02:16.38" />
                    <SPLIT distance="150" swimtime="00:03:33.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1387" points="435" reactiontime="+76" swimtime="00:04:13.42" resultid="4448" heatid="8067" lane="2" entrytime="00:04:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.25" />
                    <SPLIT distance="100" swimtime="00:02:05.22" />
                    <SPLIT distance="150" swimtime="00:03:12.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="250" reactiontime="+83" swimtime="00:02:05.79" resultid="4449" heatid="8078" lane="8" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="283" reactiontime="+96" swimtime="00:02:10.11" resultid="4450" heatid="8119" lane="5" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1584" points="305" reactiontime="+88" swimtime="00:09:15.91" resultid="4451" heatid="8161" lane="3" entrytime="00:09:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.46" />
                    <SPLIT distance="100" swimtime="00:02:13.85" />
                    <SPLIT distance="150" swimtime="00:03:40.48" />
                    <SPLIT distance="200" swimtime="00:05:02.72" />
                    <SPLIT distance="250" swimtime="00:06:09.72" />
                    <SPLIT distance="300" swimtime="00:07:17.16" />
                    <SPLIT distance="350" swimtime="00:08:19.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-10-06" firstname="Arkadiusz" gender="M" lastname="Bednarek" nation="POL" athleteid="4469">
              <RESULTS>
                <RESULT eventid="1105" points="257" reactiontime="+94" swimtime="00:00:40.71" resultid="4470" heatid="7964" lane="8" entrytime="00:00:38.00" />
                <RESULT eventid="1198" points="283" reactiontime="+88" swimtime="00:01:22.73" resultid="4471" heatid="7983" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="307" reactiontime="+87" swimtime="00:00:36.43" resultid="4472" heatid="8054" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="1509" points="234" reactiontime="+89" swimtime="00:03:12.24" resultid="4473" heatid="8095" lane="6" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.07" />
                    <SPLIT distance="100" swimtime="00:01:30.86" />
                    <SPLIT distance="150" swimtime="00:02:23.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1614" status="DNS" swimtime="00:00:00.00" resultid="4474" heatid="8133" lane="6" entrytime="00:02:55.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" />
                    <RELAYPOSITION athleteid="4444" number="2" />
                    <RELAYPOSITION athleteid="4469" number="3" />
                    <RELAYPOSITION athleteid="4452" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SOPMAST" nation="POL" region="POM" clubid="4488" name="Sopot Masters">
          <CONTACT city="SOPOT" email="sopotmasters@o2.pl" internet="www.sopotmasters.pl" name="Gorbaczow Mirosław" phone="696 258 185" state="POMOR" street="ul. Haffnera 57" zip="81-715" />
          <ATHLETES>
            <ATHLETE birthdate="1979-04-20" firstname="Piotr" gender="M" lastname="Suwara" nation="POL" athleteid="4502">
              <RESULTS>
                <RESULT eventid="1135" points="561" reactiontime="+92" swimtime="00:10:49.31" resultid="4503" heatid="8139" lane="3" entrytime="00:10:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                    <SPLIT distance="100" swimtime="00:01:16.02" />
                    <SPLIT distance="150" swimtime="00:01:56.89" />
                    <SPLIT distance="200" swimtime="00:02:38.38" />
                    <SPLIT distance="250" swimtime="00:03:20.22" />
                    <SPLIT distance="300" swimtime="00:04:02.48" />
                    <SPLIT distance="350" swimtime="00:04:44.02" />
                    <SPLIT distance="400" swimtime="00:05:26.02" />
                    <SPLIT distance="450" swimtime="00:06:07.73" />
                    <SPLIT distance="500" swimtime="00:06:49.20" />
                    <SPLIT distance="550" swimtime="00:07:30.66" />
                    <SPLIT distance="600" swimtime="00:08:11.69" />
                    <SPLIT distance="650" swimtime="00:08:53.05" />
                    <SPLIT distance="700" swimtime="00:09:33.58" />
                    <SPLIT distance="750" swimtime="00:10:12.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="571" reactiontime="+86" swimtime="00:01:02.63" resultid="4504" heatid="7990" lane="7" entrytime="00:01:02.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="504" reactiontime="+91" swimtime="00:02:47.78" resultid="4505" heatid="8026" lane="2" entrytime="00:02:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.98" />
                    <SPLIT distance="100" swimtime="00:01:21.28" />
                    <SPLIT distance="150" swimtime="00:02:05.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" status="DNS" swimtime="00:00:00.00" resultid="4506" heatid="8040" lane="2" entrytime="00:01:19.00" entrycourse="LCM" />
                <RESULT eventid="1432" points="562" reactiontime="+90" swimtime="00:05:10.77" resultid="4507" heatid="8152" lane="3" entrytime="00:05:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                    <SPLIT distance="100" swimtime="00:01:11.33" />
                    <SPLIT distance="150" swimtime="00:01:51.31" />
                    <SPLIT distance="200" swimtime="00:02:32.05" />
                    <SPLIT distance="250" swimtime="00:03:12.36" />
                    <SPLIT distance="300" swimtime="00:03:53.37" />
                    <SPLIT distance="350" swimtime="00:04:33.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="515" reactiontime="+91" swimtime="00:02:24.24" resultid="4508" heatid="8100" lane="5" entrytime="00:02:21.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                    <SPLIT distance="100" swimtime="00:01:07.96" />
                    <SPLIT distance="150" swimtime="00:01:45.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-12-28" firstname="Dariusz" gender="M" lastname="Gorbaczow" nation="POL" athleteid="4489">
              <RESULTS>
                <RESULT eventid="1105" points="782" reactiontime="+77" swimtime="00:00:30.96" resultid="4490" heatid="7968" lane="8" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="1198" points="709" reactiontime="+86" swimtime="00:01:08.13" resultid="4491" heatid="7987" lane="2" entrytime="00:01:06.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="733" reactiontime="+106" swimtime="00:01:19.83" resultid="4492" heatid="8039" lane="7" entrytime="00:01:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="718" reactiontime="+79" swimtime="00:00:29.71" resultid="4493" heatid="8057" lane="2" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT eventid="1539" points="815" reactiontime="+84" swimtime="00:00:34.78" resultid="4494" heatid="8113" lane="2" entrytime="00:00:35.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-02-08" firstname="Anna" gender="F" lastname="Maciejowska" nation="POL" athleteid="4495">
              <RESULTS>
                <RESULT eventid="1090" points="562" reactiontime="+88" swimtime="00:00:41.95" resultid="4496" heatid="7957" lane="0" entrytime="00:00:41.00" entrycourse="LCM" />
                <RESULT eventid="1120" points="642" reactiontime="+96" swimtime="00:13:45.53" resultid="4497" heatid="8137" lane="2" entrytime="00:13:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.58" />
                    <SPLIT distance="100" swimtime="00:01:34.08" />
                    <SPLIT distance="150" swimtime="00:02:26.21" />
                    <SPLIT distance="200" swimtime="00:03:18.36" />
                    <SPLIT distance="250" swimtime="00:04:09.64" />
                    <SPLIT distance="300" swimtime="00:05:02.62" />
                    <SPLIT distance="350" swimtime="00:05:55.32" />
                    <SPLIT distance="400" swimtime="00:06:48.48" />
                    <SPLIT distance="450" swimtime="00:07:41.00" />
                    <SPLIT distance="500" swimtime="00:08:33.52" />
                    <SPLIT distance="550" swimtime="00:09:26.75" />
                    <SPLIT distance="600" swimtime="00:10:19.17" />
                    <SPLIT distance="650" swimtime="00:11:12.44" />
                    <SPLIT distance="700" swimtime="00:12:04.30" />
                    <SPLIT distance="750" swimtime="00:12:54.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="578" reactiontime="+90" swimtime="00:01:22.98" resultid="4498" heatid="7976" lane="0" entrytime="00:01:21.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="642" reactiontime="+79" swimtime="00:00:35.78" resultid="4499" heatid="8046" lane="6" entrytime="00:00:36.00" entrycourse="LCM" />
                <RESULT eventid="1417" points="700" reactiontime="+94" swimtime="00:06:28.85" resultid="4500" heatid="8149" lane="4" entrytime="00:06:35.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.88" />
                    <SPLIT distance="100" swimtime="00:01:30.02" />
                    <SPLIT distance="150" swimtime="00:02:19.44" />
                    <SPLIT distance="200" swimtime="00:03:10.00" />
                    <SPLIT distance="250" swimtime="00:03:59.80" />
                    <SPLIT distance="300" swimtime="00:04:50.19" />
                    <SPLIT distance="350" swimtime="00:05:40.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="618" reactiontime="+86" swimtime="00:03:04.11" resultid="4501" heatid="8089" lane="4" entrytime="00:03:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.98" />
                    <SPLIT distance="100" swimtime="00:01:28.16" />
                    <SPLIT distance="150" swimtime="00:02:16.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="07514" nation="POL" region="WAR" clubid="4509" name="Squatina Ostrołęka">
          <CONTACT city="Ostrołęka" email="biezunskamaja@gmail.com" name="Bieżuńska Maja" phone="666353028" state="MAZ" street="Łęczysk 10/14 m.26" zip="07-410" />
          <ATHLETES>
            <ATHLETE birthdate="1979-06-26" firstname="Maja" gender="F" lastname="Bieżuńska" nation="POL" athleteid="4510">
              <RESULTS>
                <RESULT eventid="1213" points="588" reactiontime="+91" swimtime="00:00:40.14" resultid="4511" heatid="7999" lane="9" entrytime="00:00:40.05" />
                <RESULT eventid="1387" points="578" reactiontime="+95" swimtime="00:03:20.65" resultid="4512" heatid="8069" lane="6" entrytime="00:03:21.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.66" />
                    <SPLIT distance="100" swimtime="00:01:34.80" />
                    <SPLIT distance="150" swimtime="00:02:27.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="563" reactiontime="+92" swimtime="00:01:31.23" resultid="4513" heatid="8123" lane="9" entrytime="00:01:29.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="WIE" clubid="4514" name="Start Poznań">
          <CONTACT city="Poznań" email="robert.beym@gmail.com" name="Beym Robert" phone="512111513" street="os. Batorego 8/67" zip="60-687" />
          <ATHLETES>
            <ATHLETE birthdate="1967-06-06" firstname="Piotr" gender="M" lastname="Monczak" nation="POL" athleteid="4523">
              <RESULTS>
                <RESULT eventid="1075" points="895" reactiontime="+72" swimtime="00:02:31.33" resultid="4524" heatid="7952" lane="5" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                    <SPLIT distance="100" swimtime="00:01:12.22" />
                    <SPLIT distance="150" swimtime="00:01:57.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="896" reactiontime="+74" swimtime="00:00:57.93" resultid="4525" heatid="7992" lane="7" entrytime="00:00:58.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="820" reactiontime="+79" swimtime="00:00:26.88" resultid="4526" heatid="8062" lane="3" entrytime="00:00:27.20" />
                <RESULT eventid="1432" points="689" reactiontime="+82" swimtime="00:04:50.06" resultid="4527" heatid="8151" lane="8" entrytime="00:04:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                    <SPLIT distance="100" swimtime="00:01:10.80" />
                    <SPLIT distance="150" swimtime="00:01:48.87" />
                    <SPLIT distance="200" swimtime="00:02:26.62" />
                    <SPLIT distance="250" swimtime="00:03:03.86" />
                    <SPLIT distance="300" swimtime="00:03:40.98" />
                    <SPLIT distance="350" swimtime="00:04:16.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="750" reactiontime="+77" swimtime="00:02:11.34" resultid="4528" heatid="8102" lane="8" entrytime="00:02:10.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.16" />
                    <SPLIT distance="100" swimtime="00:01:05.46" />
                    <SPLIT distance="150" swimtime="00:01:38.83" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1599" points="831" reactiontime="+85" swimtime="00:05:32.19" resultid="4529" heatid="8162" lane="7" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                    <SPLIT distance="100" swimtime="00:01:15.15" />
                    <SPLIT distance="150" swimtime="00:01:59.70" />
                    <SPLIT distance="200" swimtime="00:02:43.37" />
                    <SPLIT distance="250" swimtime="00:03:31.92" />
                    <SPLIT distance="300" swimtime="00:04:21.02" />
                    <SPLIT distance="350" swimtime="00:04:57.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-06-06" firstname="Joanna" gender="F" lastname="Kostencka" nation="POL" athleteid="4530">
              <RESULTS>
                <RESULT eventid="1058" points="542" reactiontime="+89" swimtime="00:02:58.24" resultid="4531" heatid="7944" lane="1" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.82" />
                    <SPLIT distance="100" swimtime="00:01:21.98" />
                    <SPLIT distance="150" swimtime="00:02:16.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="567" swimtime="00:01:10.95" resultid="4532" heatid="7978" lane="9" entrytime="00:01:12.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="644" reactiontime="+85" swimtime="00:02:50.06" resultid="4533" heatid="8021" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.14" />
                    <SPLIT distance="100" swimtime="00:01:21.11" />
                    <SPLIT distance="150" swimtime="00:02:05.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="643" reactiontime="+78" swimtime="00:01:18.51" resultid="4534" heatid="8035" lane="2" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="577" reactiontime="+83" swimtime="00:00:32.48" resultid="4535" heatid="8048" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1524" points="600" reactiontime="+79" swimtime="00:00:36.86" resultid="4536" heatid="8107" lane="0" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-06-06" firstname="Aneta" gender="F" lastname="Maduzia" nation="POL" athleteid="4537">
              <RESULTS>
                <RESULT eventid="1058" points="385" reactiontime="+91" swimtime="00:03:21.41" resultid="4538" heatid="7942" lane="3" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.88" />
                    <SPLIT distance="100" swimtime="00:01:33.49" />
                    <SPLIT distance="150" swimtime="00:02:34.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="434" reactiontime="+91" swimtime="00:01:17.84" resultid="4539" heatid="7975" lane="4" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="482" reactiontime="+86" swimtime="00:00:34.61" resultid="4540" heatid="8047" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="1417" points="421" reactiontime="+86" swimtime="00:06:05.43" resultid="4541" heatid="8148" lane="8" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.44" />
                    <SPLIT distance="100" swimtime="00:01:27.02" />
                    <SPLIT distance="150" swimtime="00:02:13.10" />
                    <SPLIT distance="200" swimtime="00:03:00.00" />
                    <SPLIT distance="250" swimtime="00:03:47.17" />
                    <SPLIT distance="300" swimtime="00:04:34.20" />
                    <SPLIT distance="350" swimtime="00:05:20.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="413" reactiontime="+85" swimtime="00:02:51.69" resultid="4542" heatid="8090" lane="9" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.82" />
                    <SPLIT distance="100" swimtime="00:01:22.06" />
                    <SPLIT distance="150" swimtime="00:02:07.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="364" reactiontime="+88" swimtime="00:01:42.39" resultid="4543" heatid="8120" lane="7" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-06-06" firstname="Robert" gender="M" lastname="Beym" nation="POL" athleteid="4515">
              <RESULTS>
                <RESULT eventid="1075" points="873" reactiontime="+80" swimtime="00:02:32.57" resultid="4516" heatid="7951" lane="9" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                    <SPLIT distance="100" swimtime="00:01:09.87" />
                    <SPLIT distance="150" swimtime="00:01:55.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="4517" heatid="7990" lane="2" entrytime="00:01:02.00" />
                <RESULT eventid="1288" points="787" reactiontime="+66" swimtime="00:02:33.38" resultid="4518" heatid="8027" lane="7" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.52" />
                    <SPLIT distance="100" swimtime="00:01:13.78" />
                    <SPLIT distance="150" swimtime="00:01:53.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="762" reactiontime="+68" swimtime="00:01:09.96" resultid="4519" heatid="8039" lane="9" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="788" reactiontime="+82" swimtime="00:00:27.24" resultid="4520" heatid="8062" lane="0" entrytime="00:00:27.90" />
                <RESULT eventid="1539" points="734" reactiontime="+62" swimtime="00:00:32.41" resultid="4521" heatid="8115" lane="7" entrytime="00:00:33.00" />
                <RESULT eventid="1599" status="DNS" swimtime="00:00:00.00" resultid="4522" heatid="8163" lane="2" entrytime="00:06:00.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="STEEF" nation="POL" region="DOL" clubid="4544" name="STEEF Wrocław">
          <CONTACT city="Wrocław" email="ste1@wp.pl" name="Skrzypek Stefan" phone="500388374" street="Edyty Stein 6/1" zip="50-322" />
          <ATHLETES>
            <ATHLETE birthdate="1956-09-02" firstname="Stefan" gender="M" lastname="Skrzypek" nation="POL" athleteid="4554">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="4555" heatid="7948" lane="4" entrytime="00:03:15.00" />
                <RESULT eventid="1165" points="473" reactiontime="+100" swimtime="00:25:19.07" resultid="4556" heatid="8144" lane="0" entrytime="00:24:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.20" />
                    <SPLIT distance="100" swimtime="00:01:33.31" />
                    <SPLIT distance="150" swimtime="00:02:24.07" />
                    <SPLIT distance="200" swimtime="00:03:14.76" />
                    <SPLIT distance="250" swimtime="00:04:04.72" />
                    <SPLIT distance="300" swimtime="00:04:56.43" />
                    <SPLIT distance="350" swimtime="00:05:47.04" />
                    <SPLIT distance="400" swimtime="00:06:37.65" />
                    <SPLIT distance="450" swimtime="00:07:28.28" />
                    <SPLIT distance="500" swimtime="00:08:20.56" />
                    <SPLIT distance="550" swimtime="00:09:11.25" />
                    <SPLIT distance="600" swimtime="00:10:02.88" />
                    <SPLIT distance="650" swimtime="00:10:53.01" />
                    <SPLIT distance="700" swimtime="00:11:43.34" />
                    <SPLIT distance="750" swimtime="00:12:34.00" />
                    <SPLIT distance="800" swimtime="00:13:24.78" />
                    <SPLIT distance="850" swimtime="00:14:15.90" />
                    <SPLIT distance="900" swimtime="00:15:08.11" />
                    <SPLIT distance="950" swimtime="00:15:59.38" />
                    <SPLIT distance="1000" swimtime="00:16:51.73" />
                    <SPLIT distance="1050" swimtime="00:17:41.60" />
                    <SPLIT distance="1100" swimtime="00:18:33.08" />
                    <SPLIT distance="1150" swimtime="00:19:23.35" />
                    <SPLIT distance="1200" swimtime="00:20:14.86" />
                    <SPLIT distance="1250" swimtime="00:21:06.07" />
                    <SPLIT distance="1300" swimtime="00:21:57.94" />
                    <SPLIT distance="1350" swimtime="00:22:49.53" />
                    <SPLIT distance="1400" swimtime="00:23:42.26" />
                    <SPLIT distance="1450" swimtime="00:24:31.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" status="DNS" swimtime="00:00:00.00" resultid="4557" heatid="8015" lane="5" entrytime="00:03:20.00" />
                <RESULT eventid="1432" points="523" reactiontime="+98" swimtime="00:06:06.15" resultid="4558" heatid="8154" lane="6" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.36" />
                    <SPLIT distance="100" swimtime="00:01:30.68" />
                    <SPLIT distance="150" swimtime="00:02:18.67" />
                    <SPLIT distance="200" swimtime="00:03:06.12" />
                    <SPLIT distance="250" swimtime="00:03:51.96" />
                    <SPLIT distance="300" swimtime="00:04:37.29" />
                    <SPLIT distance="350" swimtime="00:05:22.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" status="DNS" swimtime="00:00:00.00" resultid="4559" heatid="8083" lane="7" entrytime="00:01:30.00" />
                <RESULT eventid="1509" points="512" reactiontime="+98" swimtime="00:02:50.13" resultid="4560" heatid="8097" lane="8" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.99" />
                    <SPLIT distance="100" swimtime="00:01:23.39" />
                    <SPLIT distance="150" swimtime="00:02:06.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" status="DNS" swimtime="00:00:00.00" resultid="4561" heatid="8165" lane="6" entrytime="00:07:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-03-19" firstname="Ewa" gender="F" lastname="Szała" nation="POL" athleteid="4545">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1058" points="847" reactiontime="+89" swimtime="00:03:03.57" resultid="4546" heatid="7943" lane="6" entrytime="00:03:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.33" />
                    <SPLIT distance="100" swimtime="00:01:26.34" />
                    <SPLIT distance="150" swimtime="00:02:20.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="874" reactiontime="+97" swimtime="00:12:24.97" resultid="4547" heatid="8136" lane="0" entrytime="00:12:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.33" />
                    <SPLIT distance="100" swimtime="00:01:25.96" />
                    <SPLIT distance="150" swimtime="00:02:12.52" />
                    <SPLIT distance="200" swimtime="00:02:59.51" />
                    <SPLIT distance="250" swimtime="00:03:46.79" />
                    <SPLIT distance="300" swimtime="00:04:34.15" />
                    <SPLIT distance="350" swimtime="00:05:21.27" />
                    <SPLIT distance="400" swimtime="00:06:08.20" />
                    <SPLIT distance="450" swimtime="00:06:54.83" />
                    <SPLIT distance="500" swimtime="00:07:42.28" />
                    <SPLIT distance="550" swimtime="00:08:29.19" />
                    <SPLIT distance="600" swimtime="00:09:16.49" />
                    <SPLIT distance="650" swimtime="00:10:03.25" />
                    <SPLIT distance="700" swimtime="00:10:50.89" />
                    <SPLIT distance="750" swimtime="00:11:37.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="575" reactiontime="+94" swimtime="00:01:23.12" resultid="4548" heatid="7977" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.49" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1273" points="855" reactiontime="+92" swimtime="00:03:03.88" resultid="4549" heatid="8020" lane="1" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.00" />
                    <SPLIT distance="100" swimtime="00:01:31.06" />
                    <SPLIT distance="150" swimtime="00:02:17.91" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1326" points="803" reactiontime="+91" swimtime="00:01:26.98" resultid="4550" heatid="8034" lane="7" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.16" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1447" points="671" reactiontime="+92" swimtime="00:01:30.53" resultid="4551" heatid="8079" lane="1" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="706" reactiontime="+87" swimtime="00:00:40.91" resultid="4552" heatid="8105" lane="6" entrytime="00:00:41.00" />
                <RESULT eventid="1584" points="871" reactiontime="+95" swimtime="00:06:31.99" resultid="4553" heatid="8160" lane="6" entrytime="00:06:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.47" />
                    <SPLIT distance="100" swimtime="00:01:34.75" />
                    <SPLIT distance="150" swimtime="00:02:24.74" />
                    <SPLIT distance="200" swimtime="00:03:13.61" />
                    <SPLIT distance="250" swimtime="00:04:08.41" />
                    <SPLIT distance="300" swimtime="00:05:03.17" />
                    <SPLIT distance="350" swimtime="00:05:48.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="POL" nation="POL" region="LOD" clubid="4433" name="Stowarzyszenie Przyjaciół Pływania" shortname="Stowarzyszenie Przyjaciół Pływ">
          <CONTACT city="Bełchatów" email="piotreksiewiera@wp.pl" internet="www.wejdzdowody.pl" name="Siewiera" phone="667923503" state="ŁÓDZK" street="ul Słoneczna 57" zip="97-400" />
          <ATHLETES>
            <ATHLETE birthdate="1994-06-07" firstname="Piotr" gender="M" lastname="Siewiera" nation="POL" license="AFD082521" athleteid="4434">
              <RESULTS>
                <RESULT eventid="1105" points="421" reactiontime="+92" swimtime="00:00:33.69" resultid="4435" heatid="7961" lane="3" />
                <RESULT eventid="1135" points="410" swimtime="00:11:23.36" resultid="4436" heatid="8141" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.37" />
                    <SPLIT distance="100" swimtime="00:01:13.75" />
                    <SPLIT distance="150" swimtime="00:01:55.56" />
                    <SPLIT distance="200" swimtime="00:02:38.89" />
                    <SPLIT distance="250" swimtime="00:03:22.44" />
                    <SPLIT distance="300" swimtime="00:04:06.72" />
                    <SPLIT distance="350" swimtime="00:04:51.11" />
                    <SPLIT distance="400" swimtime="00:05:35.94" />
                    <SPLIT distance="450" swimtime="00:06:19.40" />
                    <SPLIT distance="500" swimtime="00:07:03.16" />
                    <SPLIT distance="550" swimtime="00:07:47.94" />
                    <SPLIT distance="600" swimtime="00:08:31.88" />
                    <SPLIT distance="650" swimtime="00:09:16.86" />
                    <SPLIT distance="700" swimtime="00:10:00.50" />
                    <SPLIT distance="750" swimtime="00:10:42.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="635" reactiontime="+89" swimtime="00:01:00.16" resultid="4437" heatid="7991" lane="8" entrytime="00:01:00.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="500" reactiontime="+77" swimtime="00:02:40.08" resultid="4438" heatid="8022" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.52" />
                    <SPLIT distance="100" swimtime="00:01:17.92" />
                    <SPLIT distance="150" swimtime="00:01:59.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="511" reactiontime="+79" swimtime="00:01:12.99" resultid="4439" heatid="8042" lane="0" entrytime="00:01:10.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="614" reactiontime="+99" swimtime="00:00:27.09" resultid="4440" heatid="8064" lane="2" entrytime="00:00:26.06" entrycourse="SCM" />
                <RESULT eventid="1509" points="512" reactiontime="+108" swimtime="00:02:24.51" resultid="4441" heatid="8093" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.55" />
                    <SPLIT distance="100" swimtime="00:01:06.25" />
                    <SPLIT distance="150" swimtime="00:01:47.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="546" reactiontime="+76" swimtime="00:00:33.33" resultid="4442" heatid="8108" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SMMK" nation="POL" region="MAL" clubid="3953" name="Straż Miejska Miasta Kraków">
          <CONTACT city="Kraków" name="Jawień Krzysztof" phone="500677133" state="MAŁ" />
          <ATHLETES>
            <ATHLETE birthdate="1971-06-11" firstname="Krzysztof" gender="M" lastname="Jawień" nation="POL" athleteid="3955">
              <RESULTS>
                <RESULT eventid="1075" points="524" reactiontime="+80" swimtime="00:02:44.20" resultid="3956" heatid="7946" lane="1" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                    <SPLIT distance="100" swimtime="00:01:15.98" />
                    <SPLIT distance="150" swimtime="00:02:02.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="391" reactiontime="+82" swimtime="00:11:59.94" resultid="3957" heatid="8139" lane="2" entrytime="00:10:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                    <SPLIT distance="100" swimtime="00:01:18.15" />
                    <SPLIT distance="150" swimtime="00:02:01.96" />
                    <SPLIT distance="200" swimtime="00:02:47.63" />
                    <SPLIT distance="250" swimtime="00:03:34.27" />
                    <SPLIT distance="300" swimtime="00:04:20.92" />
                    <SPLIT distance="350" swimtime="00:05:07.69" />
                    <SPLIT distance="400" swimtime="00:05:54.43" />
                    <SPLIT distance="450" swimtime="00:06:41.10" />
                    <SPLIT distance="500" swimtime="00:07:27.18" />
                    <SPLIT distance="550" swimtime="00:08:13.22" />
                    <SPLIT distance="600" swimtime="00:08:58.89" />
                    <SPLIT distance="650" swimtime="00:09:44.93" />
                    <SPLIT distance="700" swimtime="00:10:30.87" />
                    <SPLIT distance="750" swimtime="00:11:15.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="623" reactiontime="+76" swimtime="00:00:35.72" resultid="3958" heatid="8002" lane="2" entrytime="00:00:45.00" />
                <RESULT eventid="1288" points="503" reactiontime="+71" swimtime="00:02:50.47" resultid="3959" heatid="8025" lane="5" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.04" />
                    <SPLIT distance="100" swimtime="00:01:22.95" />
                    <SPLIT distance="150" swimtime="00:02:07.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="542" reactiontime="+67" swimtime="00:01:17.17" resultid="3960" heatid="8036" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="612" reactiontime="+74" swimtime="00:02:57.62" resultid="3961" heatid="8076" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.01" />
                    <SPLIT distance="100" swimtime="00:01:25.29" />
                    <SPLIT distance="150" swimtime="00:02:11.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="618" reactiontime="+79" swimtime="00:01:20.65" resultid="3962" heatid="8124" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="479" reactiontime="+82" swimtime="00:06:01.57" resultid="3963" heatid="8163" lane="3" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                    <SPLIT distance="100" swimtime="00:01:17.63" />
                    <SPLIT distance="150" swimtime="00:02:09.00" />
                    <SPLIT distance="200" swimtime="00:02:58.90" />
                    <SPLIT distance="250" swimtime="00:03:47.97" />
                    <SPLIT distance="300" swimtime="00:04:37.58" />
                    <SPLIT distance="350" swimtime="00:05:19.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="MAZ" clubid="4568" name="Swimmerst Stowarzyszenie Pływackie" shortname="Swimmerst Stowarzyszenie Pływa">
          <CONTACT city="WARSZAWA" email="INFO@SWIMMERSTEAM.PL" name="REMIGIUSZ GOŁĘBIOWSKI" phone="601333782" state="MAZ" street="GŁADKA 18" zip="02-172" />
          <ATHLETES>
            <ATHLETE birthdate="1982-11-04" firstname="Napora" gender="M" lastname="Grzegorz" nation="POL" athleteid="4573">
              <RESULTS>
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="4574" heatid="7992" lane="9" entrytime="00:00:59.00" />
                <RESULT eventid="1372" status="DNS" swimtime="00:00:00.00" resultid="4575" heatid="8063" lane="6" entrytime="00:00:26.50" />
                <RESULT eventid="1509" status="DNS" swimtime="00:00:00.00" resultid="4576" heatid="8102" lane="6" entrytime="00:02:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-03-03" firstname="Katarzyna" gender="F" lastname="Napora" nation="POL" athleteid="4585">
              <RESULTS>
                <RESULT eventid="1090" status="DNS" swimtime="00:00:00.00" resultid="4586" heatid="7956" lane="5" entrytime="00:00:41.11" />
                <RESULT eventid="1181" points="486" reactiontime="+67" swimtime="00:01:14.96" resultid="4587" heatid="7977" lane="4" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="585" reactiontime="+66" swimtime="00:00:32.45" resultid="4588" heatid="8049" lane="8" entrytime="00:00:31.87" />
                <RESULT eventid="1417" points="396" swimtime="00:06:12.89" resultid="4589" heatid="8147" lane="9" entrytime="00:05:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.20" />
                    <SPLIT distance="100" swimtime="00:01:20.93" />
                    <SPLIT distance="150" swimtime="00:02:08.05" />
                    <SPLIT distance="200" swimtime="00:02:57.64" />
                    <SPLIT distance="250" swimtime="00:03:46.81" />
                    <SPLIT distance="300" swimtime="00:04:36.80" />
                    <SPLIT distance="350" swimtime="00:05:25.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" status="DNS" swimtime="00:00:00.00" resultid="4590" heatid="8091" lane="0" entrytime="00:02:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-12-11" firstname="Mikołaj" gender="M" lastname="Tusiński" nation="POL" athleteid="4591">
              <RESULTS>
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="4592" heatid="7966" lane="3" entrytime="00:00:33.00" />
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="4593" heatid="7991" lane="5" entrytime="00:00:59.00" />
                <RESULT eventid="1372" status="DNS" swimtime="00:00:00.00" resultid="4594" heatid="8062" lane="5" entrytime="00:00:27.00" />
                <RESULT eventid="1462" status="DNS" swimtime="00:00:00.00" resultid="4595" heatid="8085" lane="7" entrytime="00:01:09.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-12-20" firstname="Arkadiusz" gender="M" lastname="Aptewicz" nation="POL" athleteid="4580">
              <RESULTS>
                <RESULT eventid="1075" points="792" reactiontime="+71" swimtime="00:02:20.03" resultid="4581" heatid="7953" lane="3" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.39" />
                    <SPLIT distance="100" swimtime="00:01:07.17" />
                    <SPLIT distance="150" swimtime="00:01:45.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="826" reactiontime="+66" swimtime="00:00:31.12" resultid="4582" heatid="8010" lane="3" entrytime="00:00:31.40" />
                <RESULT eventid="1402" points="891" reactiontime="+70" swimtime="00:02:29.87" resultid="4583" heatid="8077" lane="5" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.87" />
                    <SPLIT distance="100" swimtime="00:01:12.83" />
                    <SPLIT distance="150" swimtime="00:01:51.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="883" reactiontime="+72" swimtime="00:01:09.19" resultid="4584" heatid="8132" lane="2" entrytime="00:01:09.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-28" firstname="Marek" gender="M" lastname="Brożyna" nation="POL" athleteid="4569">
              <RESULTS>
                <RESULT eventid="1288" points="514" reactiontime="+66" swimtime="00:02:46.68" resultid="4570" heatid="8027" lane="8" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                    <SPLIT distance="100" swimtime="00:01:17.90" />
                    <SPLIT distance="150" swimtime="00:02:01.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="581" reactiontime="+71" swimtime="00:01:14.33" resultid="4571" heatid="8041" lane="5" entrytime="00:01:12.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" status="DNS" swimtime="00:00:00.00" resultid="4572" heatid="8114" lane="6" entrytime="00:00:33.88" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-07-01" firstname="Katarzyna" gender="F" lastname="Koba" nation="POL" athleteid="4596">
              <RESULTS>
                <RESULT eventid="1090" points="494" reactiontime="+77" swimtime="00:00:35.78" resultid="4597" heatid="7958" lane="7" entrytime="00:00:37.00" />
                <RESULT eventid="1181" points="559" reactiontime="+81" swimtime="00:01:11.28" resultid="4598" heatid="7977" lane="6" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="644" reactiontime="+87" swimtime="00:00:31.31" resultid="4599" heatid="8049" lane="7" entrytime="00:00:31.50" />
                <RESULT eventid="1493" points="473" reactiontime="+80" swimtime="00:02:45.40" resultid="4600" heatid="8090" lane="4" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.73" />
                    <SPLIT distance="100" swimtime="00:01:19.59" />
                    <SPLIT distance="150" swimtime="00:02:02.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-07-07" firstname="Remigiusz" gender="M" lastname="Gołębiowski" nation="POL" athleteid="4577">
              <RESULTS>
                <RESULT eventid="1105" points="673" reactiontime="+89" swimtime="00:00:29.11" resultid="4578" heatid="7971" lane="0" entrytime="00:00:29.00" />
                <RESULT eventid="1372" points="611" reactiontime="+78" swimtime="00:00:27.72" resultid="4579" heatid="8061" lane="7" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="4601" heatid="8031" lane="7" entrytime="00:04:10.00" />
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1614" status="DNS" swimtime="00:00:00.00" resultid="4602" heatid="8135" lane="6" entrytime="00:02:10.00" />
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="4603" name="Swimming Masters Team Szczecin" shortname="SMT Szczecin">
          <CONTACT city="Szczecin" email="teczowy.dyndol@gmail.com" name="Brodacki Maciej" phone="608396939" street="Szafera 110/1" zip="71-245" />
          <ATHLETES>
            <ATHLETE birthdate="1974-08-12" firstname="Marek" gender="M" lastname="Zienkiewicz" nation="POL" athleteid="4653">
              <RESULTS>
                <RESULT eventid="1105" points="400" reactiontime="+75" swimtime="00:00:35.14" resultid="4654" heatid="7964" lane="3" entrytime="00:00:36.00" entrycourse="LCM" />
                <RESULT eventid="1198" points="359" reactiontime="+76" swimtime="00:01:16.43" resultid="4655" heatid="7983" lane="2" entrytime="00:01:22.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="490" reactiontime="+77" swimtime="00:00:31.17" resultid="4656" heatid="8056" lane="6" entrytime="00:00:31.28" entrycourse="LCM" />
                <RESULT eventid="1462" points="301" reactiontime="+84" swimtime="00:01:27.55" resultid="4657" heatid="8083" lane="0" entrytime="00:01:32.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="282" reactiontime="+78" swimtime="00:03:00.63" resultid="4658" heatid="8095" lane="8" entrytime="00:03:19.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                    <SPLIT distance="100" swimtime="00:01:25.10" />
                    <SPLIT distance="150" swimtime="00:02:12.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-11-03" firstname="Agnieszka" gender="F" lastname="Suwiczak" nation="POL" athleteid="4659">
              <RESULTS>
                <RESULT eventid="1090" points="551" reactiontime="+84" swimtime="00:00:34.50" resultid="4660" heatid="7959" lane="8" entrytime="00:00:35.00" entrycourse="LCM" />
                <RESULT eventid="1181" points="645" reactiontime="+87" swimtime="00:01:07.97" resultid="4661" heatid="7979" lane="0" entrytime="00:01:05.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="496" reactiontime="+76" swimtime="00:00:41.24" resultid="4662" heatid="7997" lane="8" entrytime="00:00:45.57" entrycourse="LCM" />
                <RESULT eventid="1357" points="725" reactiontime="+78" swimtime="00:00:30.10" resultid="4663" heatid="8049" lane="3" entrytime="00:00:29.99" entrycourse="LCM" />
                <RESULT eventid="1493" status="DNS" swimtime="00:00:00.00" resultid="4664" heatid="8092" lane="9" entrytime="00:02:30.00" entrycourse="LCM" />
                <RESULT eventid="1524" points="657" reactiontime="+73" swimtime="00:00:35.76" resultid="4665" heatid="8107" lane="8" entrytime="00:00:35.60" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1995-07-21" firstname="Wiktoria" gender="F" lastname="Podkowińska" nation="POL" athleteid="4612">
              <RESULTS>
                <RESULT eventid="1058" points="572" reactiontime="+70" swimtime="00:02:56.46" resultid="4613" heatid="7943" lane="4" entrytime="00:02:59.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.62" />
                    <SPLIT distance="100" swimtime="00:01:24.51" />
                    <SPLIT distance="150" swimtime="00:02:16.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="511" reactiontime="+71" swimtime="00:00:34.87" resultid="4614" heatid="7958" lane="3" entrytime="00:00:36.00" entrycourse="LCM" />
                <RESULT eventid="1181" points="592" reactiontime="+73" swimtime="00:01:09.88" resultid="4615" heatid="7977" lane="3" entrytime="00:01:13.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="540" reactiontime="+69" swimtime="00:00:32.68" resultid="4616" heatid="8049" lane="0" entrytime="00:00:31.98" entrycourse="LCM" />
                <RESULT eventid="1447" points="395" reactiontime="+66" swimtime="00:01:26.37" resultid="4617" heatid="8080" lane="9" entrytime="00:01:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1584" points="475" reactiontime="+79" swimtime="00:06:23.86" resultid="4618" heatid="8160" lane="7" entrytime="00:06:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.17" />
                    <SPLIT distance="100" swimtime="00:01:30.19" />
                    <SPLIT distance="150" swimtime="00:02:23.70" />
                    <SPLIT distance="200" swimtime="00:03:14.38" />
                    <SPLIT distance="250" swimtime="00:04:07.60" />
                    <SPLIT distance="300" swimtime="00:05:01.83" />
                    <SPLIT distance="350" swimtime="00:05:44.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-20" firstname="Agnieszka" gender="F" lastname="Krzyżostaniak" nation="POL" athleteid="4619">
              <RESULTS>
                <RESULT eventid="1120" points="764" reactiontime="+75" swimtime="00:10:13.13" resultid="4620" heatid="8136" lane="4" entrytime="00:10:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.53" />
                    <SPLIT distance="100" swimtime="00:01:08.93" />
                    <SPLIT distance="150" swimtime="00:01:46.49" />
                    <SPLIT distance="200" swimtime="00:02:24.61" />
                    <SPLIT distance="250" swimtime="00:03:03.12" />
                    <SPLIT distance="300" swimtime="00:03:41.74" />
                    <SPLIT distance="350" swimtime="00:04:20.32" />
                    <SPLIT distance="400" swimtime="00:04:59.52" />
                    <SPLIT distance="450" swimtime="00:05:38.71" />
                    <SPLIT distance="500" swimtime="00:06:17.63" />
                    <SPLIT distance="550" swimtime="00:06:56.58" />
                    <SPLIT distance="600" swimtime="00:07:36.45" />
                    <SPLIT distance="650" swimtime="00:08:15.77" />
                    <SPLIT distance="700" swimtime="00:08:56.37" />
                    <SPLIT distance="750" swimtime="00:09:35.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="760" reactiontime="+77" swimtime="00:00:29.16" resultid="4621" heatid="8049" lane="6" entrytime="00:00:30.00" entrycourse="LCM" />
                <RESULT eventid="1417" points="750" reactiontime="+80" swimtime="00:04:55.56" resultid="4622" heatid="8147" lane="3" entrytime="00:05:05.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.00" />
                    <SPLIT distance="100" swimtime="00:01:11.71" />
                    <SPLIT distance="150" swimtime="00:01:48.91" />
                    <SPLIT distance="200" swimtime="00:02:26.44" />
                    <SPLIT distance="250" swimtime="00:03:03.64" />
                    <SPLIT distance="300" swimtime="00:03:41.08" />
                    <SPLIT distance="350" swimtime="00:04:19.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="879" reactiontime="+70" swimtime="00:00:32.55" resultid="4623" heatid="8107" lane="5" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="1584" points="662" reactiontime="+83" swimtime="00:05:43.76" resultid="4624" heatid="8159" lane="6" entrytime="00:06:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                    <SPLIT distance="100" swimtime="00:01:23.48" />
                    <SPLIT distance="150" swimtime="00:02:06.53" />
                    <SPLIT distance="200" swimtime="00:02:48.72" />
                    <SPLIT distance="250" swimtime="00:03:38.25" />
                    <SPLIT distance="300" swimtime="00:04:28.08" />
                    <SPLIT distance="350" swimtime="00:05:06.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-06-14" firstname="Kinga" gender="F" lastname="Maciupa" nation="POL" athleteid="4666">
              <RESULTS>
                <RESULT eventid="1090" points="609" reactiontime="+66" swimtime="00:00:32.89" resultid="4667" heatid="7960" lane="2" entrytime="00:00:31.80" entrycourse="LCM" />
                <RESULT eventid="1273" points="732" reactiontime="+65" swimtime="00:02:40.77" resultid="4668" heatid="8021" lane="4" entrytime="00:02:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                    <SPLIT distance="100" swimtime="00:01:16.51" />
                    <SPLIT distance="150" swimtime="00:01:58.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="777" reactiontime="+69" swimtime="00:01:13.45" resultid="4669" heatid="8035" lane="4" entrytime="00:01:08.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="519" reactiontime="+65" swimtime="00:00:33.12" resultid="4670" heatid="8049" lane="4" entrytime="00:00:29.50" entrycourse="LCM" />
                <RESULT eventid="1524" points="760" reactiontime="+65" swimtime="00:00:34.17" resultid="4671" heatid="8107" lane="3" entrytime="00:00:32.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-02-24" firstname="Maciej" gender="M" lastname="Brodacki" nation="POL" athleteid="4637">
              <RESULTS>
                <RESULT eventid="1075" points="723" reactiontime="+76" swimtime="00:02:26.61" resultid="4638" heatid="7952" lane="6" entrytime="00:02:36.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.72" />
                    <SPLIT distance="100" swimtime="00:01:07.20" />
                    <SPLIT distance="150" swimtime="00:01:51.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="620" reactiontime="+70" swimtime="00:00:29.33" resultid="4639" heatid="7967" lane="9" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT eventid="1198" points="723" reactiontime="+78" swimtime="00:00:56.64" resultid="4640" heatid="7992" lane="2" entrytime="00:00:58.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="4641" heatid="8026" lane="8" entrytime="00:02:50.00" entrycourse="LCM" />
                <RESULT eventid="1372" points="727" reactiontime="+77" swimtime="00:00:25.85" resultid="4642" heatid="8063" lane="3" entrytime="00:00:26.50" entrycourse="LCM" />
                <RESULT eventid="1432" points="598" reactiontime="+87" swimtime="00:04:54.99" resultid="4643" heatid="8152" lane="7" entrytime="00:05:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                    <SPLIT distance="100" swimtime="00:01:09.81" />
                    <SPLIT distance="150" swimtime="00:01:47.71" />
                    <SPLIT distance="200" swimtime="00:02:25.90" />
                    <SPLIT distance="250" swimtime="00:03:04.16" />
                    <SPLIT distance="300" swimtime="00:03:41.53" />
                    <SPLIT distance="350" swimtime="00:04:19.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="650" reactiontime="+84" swimtime="00:02:13.53" resultid="4644" heatid="8101" lane="0" entrytime="00:02:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.96" />
                    <SPLIT distance="100" swimtime="00:01:03.47" />
                    <SPLIT distance="150" swimtime="00:01:38.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="574" reactiontime="+99" swimtime="00:05:29.48" resultid="4645" heatid="8162" lane="0" entrytime="00:05:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                    <SPLIT distance="100" swimtime="00:01:13.73" />
                    <SPLIT distance="150" swimtime="00:01:57.22" />
                    <SPLIT distance="200" swimtime="00:02:40.01" />
                    <SPLIT distance="250" swimtime="00:03:27.65" />
                    <SPLIT distance="300" swimtime="00:04:15.97" />
                    <SPLIT distance="350" swimtime="00:04:54.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-11-22" firstname="Michał" gender="M" lastname="Bałka" nation="POL" athleteid="4646">
              <RESULTS>
                <RESULT eventid="1075" points="468" reactiontime="+81" swimtime="00:02:42.22" resultid="4647" heatid="7951" lane="6" entrytime="00:02:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.69" />
                    <SPLIT distance="100" swimtime="00:01:11.34" />
                    <SPLIT distance="150" swimtime="00:02:00.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="562" reactiontime="+81" swimtime="00:00:30.37" resultid="4648" heatid="7966" lane="5" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT eventid="1258" points="511" reactiontime="+90" swimtime="00:02:40.30" resultid="4649" heatid="8017" lane="8" entrytime="00:02:35.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                    <SPLIT distance="100" swimtime="00:01:12.74" />
                    <SPLIT distance="150" swimtime="00:01:55.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="534" reactiontime="+69" swimtime="00:00:28.52" resultid="4650" heatid="8059" lane="8" entrytime="00:00:29.00" entrycourse="LCM" />
                <RESULT eventid="1462" points="545" reactiontime="+81" swimtime="00:01:09.58" resultid="4651" heatid="8085" lane="0" entrytime="00:01:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="523" reactiontime="+95" swimtime="00:05:54.02" resultid="4652" heatid="8163" lane="7" entrytime="00:06:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                    <SPLIT distance="100" swimtime="00:01:15.48" />
                    <SPLIT distance="150" swimtime="00:02:01.95" />
                    <SPLIT distance="200" swimtime="00:02:47.61" />
                    <SPLIT distance="250" swimtime="00:03:40.28" />
                    <SPLIT distance="300" swimtime="00:04:32.74" />
                    <SPLIT distance="350" swimtime="00:05:13.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-09" firstname="Helena" gender="F" lastname="Szulc" nation="POL" athleteid="4630">
              <RESULTS>
                <RESULT eventid="1058" points="527" reactiontime="+91" swimtime="00:02:59.87" resultid="4631" heatid="7944" lane="0" entrytime="00:02:56.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.39" />
                    <SPLIT distance="100" swimtime="00:01:24.34" />
                    <SPLIT distance="150" swimtime="00:02:17.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="450" reactiontime="+82" swimtime="00:00:36.92" resultid="4632" heatid="7958" lane="2" entrytime="00:00:37.00" entrycourse="LCM" />
                <RESULT eventid="1213" points="340" reactiontime="+78" swimtime="00:00:46.75" resultid="4633" heatid="7997" lane="9" entrytime="00:00:46.00" entrycourse="LCM" />
                <RESULT eventid="1243" points="375" reactiontime="+105" swimtime="00:03:23.16" resultid="4634" heatid="8012" lane="1" entrytime="00:03:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.59" />
                    <SPLIT distance="100" swimtime="00:01:35.89" />
                    <SPLIT distance="150" swimtime="00:02:29.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="383" reactiontime="+71" swimtime="00:01:28.30" resultid="4635" heatid="8079" lane="8" entrytime="00:01:28.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1584" points="516" reactiontime="+94" swimtime="00:06:28.68" resultid="4636" heatid="8159" lane="0" entrytime="00:06:19.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.32" />
                    <SPLIT distance="100" swimtime="00:01:33.82" />
                    <SPLIT distance="150" swimtime="00:02:22.96" />
                    <SPLIT distance="200" swimtime="00:03:11.55" />
                    <SPLIT distance="250" swimtime="00:04:05.19" />
                    <SPLIT distance="300" swimtime="00:05:00.07" />
                    <SPLIT distance="350" swimtime="00:05:45.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-04-21" firstname="Michał" gender="M" lastname="Krysiak" nation="POL" athleteid="4625">
              <RESULTS>
                <RESULT eventid="1198" points="485" reactiontime="+76" swimtime="00:01:05.80" resultid="4626" heatid="7991" lane="7" entrytime="00:01:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" status="DNS" swimtime="00:00:00.00" resultid="4627" heatid="8017" lane="1" entrytime="00:02:33.56" entrycourse="LCM" />
                <RESULT eventid="1372" points="565" reactiontime="+79" swimtime="00:00:27.99" resultid="4628" heatid="8062" lane="6" entrytime="00:00:27.54" entrycourse="LCM" />
                <RESULT eventid="1462" points="520" reactiontime="+76" swimtime="00:01:10.67" resultid="4629" heatid="8085" lane="5" entrytime="00:01:05.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-06-12" firstname="Kamila" gender="F" lastname="Gębka" nation="POL" athleteid="4606">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="4607" heatid="7944" lane="9" entrytime="00:02:57.00" entrycourse="LCM" />
                <RESULT eventid="1213" status="DNS" swimtime="00:00:00.00" resultid="4608" heatid="7997" lane="3" entrytime="00:00:43.00" entrycourse="LCM" />
                <RESULT eventid="1387" points="483" reactiontime="+84" swimtime="00:03:18.48" resultid="4609" heatid="8070" lane="1" entrytime="00:03:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.97" />
                    <SPLIT distance="100" swimtime="00:01:35.89" />
                    <SPLIT distance="150" swimtime="00:02:27.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="468" reactiontime="+94" swimtime="00:01:33.21" resultid="4610" heatid="8122" lane="7" entrytime="00:01:31.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1584" status="DNS" swimtime="00:00:00.00" resultid="4611" heatid="8160" lane="2" entrytime="00:06:45.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1303" reactiontime="+68" swimtime="00:04:47.00" resultid="6101" heatid="8029" lane="5" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.87" />
                    <SPLIT distance="100" swimtime="00:01:11.24" />
                    <SPLIT distance="150" swimtime="00:01:45.83" />
                    <SPLIT distance="200" swimtime="00:02:26.12" />
                    <SPLIT distance="250" swimtime="00:03:00.93" />
                    <SPLIT distance="300" swimtime="00:03:39.04" />
                    <SPLIT distance="350" swimtime="00:04:11.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4612" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="4630" number="2" reactiontime="+63" />
                    <RELAYPOSITION athleteid="4606" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="4659" number="4" reactiontime="+71" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1614" reactiontime="+76" swimtime="00:02:11.13" resultid="6099" heatid="8135" lane="3" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                    <SPLIT distance="100" swimtime="00:01:15.77" />
                    <SPLIT distance="150" swimtime="00:01:45.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4619" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="4606" number="2" />
                    <RELAYPOSITION athleteid="4646" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="4637" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1614" reactiontime="+73" swimtime="00:02:23.68" resultid="6100" heatid="8135" lane="8" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.88" />
                    <SPLIT distance="100" swimtime="00:01:22.71" />
                    <SPLIT distance="150" swimtime="00:01:52.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4659" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="4630" number="2" />
                    <RELAYPOSITION athleteid="4625" number="3" reactiontime="+76" />
                    <RELAYPOSITION athleteid="4653" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5150" name="Szkoła Pływania Goleniów">
          <CONTACT name="Wierzchoń" />
          <ATHLETES>
            <ATHLETE birthdate="1962-10-01" firstname="Aleksy" gender="M" lastname="Wierzchoń" nation="POL" athleteid="5151">
              <RESULTS>
                <RESULT eventid="1165" points="420" reactiontime="+101" swimtime="00:24:12.98" resultid="5152" heatid="8144" lane="1" entrytime="00:23:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.63" />
                    <SPLIT distance="100" swimtime="00:01:22.46" />
                    <SPLIT distance="150" swimtime="00:02:08.79" />
                    <SPLIT distance="200" swimtime="00:02:55.63" />
                    <SPLIT distance="250" swimtime="00:03:43.73" />
                    <SPLIT distance="300" swimtime="00:04:32.27" />
                    <SPLIT distance="350" swimtime="00:05:20.20" />
                    <SPLIT distance="400" swimtime="00:06:07.94" />
                    <SPLIT distance="450" swimtime="00:06:56.91" />
                    <SPLIT distance="500" swimtime="00:07:45.52" />
                    <SPLIT distance="550" swimtime="00:08:34.37" />
                    <SPLIT distance="600" swimtime="00:09:22.50" />
                    <SPLIT distance="650" swimtime="00:10:11.20" />
                    <SPLIT distance="700" swimtime="00:11:00.59" />
                    <SPLIT distance="750" swimtime="00:11:48.98" />
                    <SPLIT distance="800" swimtime="00:12:37.48" />
                    <SPLIT distance="850" swimtime="00:13:26.95" />
                    <SPLIT distance="900" swimtime="00:14:16.98" />
                    <SPLIT distance="950" swimtime="00:15:05.87" />
                    <SPLIT distance="1000" swimtime="00:15:55.65" />
                    <SPLIT distance="1050" swimtime="00:16:44.36" />
                    <SPLIT distance="1100" swimtime="00:17:34.93" />
                    <SPLIT distance="1150" swimtime="00:18:24.76" />
                    <SPLIT distance="1200" swimtime="00:19:14.78" />
                    <SPLIT distance="1250" swimtime="00:20:04.54" />
                    <SPLIT distance="1300" swimtime="00:20:54.01" />
                    <SPLIT distance="1350" swimtime="00:21:43.54" />
                    <SPLIT distance="1400" swimtime="00:22:33.53" />
                    <SPLIT distance="1450" swimtime="00:23:23.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="441" reactiontime="+99" swimtime="00:00:42.27" resultid="5153" heatid="8002" lane="5" entrytime="00:00:44.00" />
                <RESULT eventid="1432" points="426" reactiontime="+101" swimtime="00:06:02.09" resultid="5154" heatid="8154" lane="7" entrytime="00:06:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.35" />
                    <SPLIT distance="100" swimtime="00:01:24.75" />
                    <SPLIT distance="150" swimtime="00:02:11.42" />
                    <SPLIT distance="200" swimtime="00:02:59.21" />
                    <SPLIT distance="250" swimtime="00:03:47.04" />
                    <SPLIT distance="300" swimtime="00:04:34.81" />
                    <SPLIT distance="350" swimtime="00:05:21.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="486" reactiontime="+105" swimtime="00:02:44.43" resultid="5155" heatid="8096" lane="4" entrytime="00:02:53.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                    <SPLIT distance="100" swimtime="00:01:19.06" />
                    <SPLIT distance="150" swimtime="00:02:03.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="4859" name="T.P Skalar Słupsk">
          <CONTACT name="Zubel Beata" />
          <ATHLETES>
            <ATHLETE birthdate="1968-09-28" firstname="Beata" gender="F" lastname="Zubel" nation="POL" athleteid="4863">
              <RESULTS>
                <RESULT eventid="1120" points="560" reactiontime="+91" swimtime="00:11:44.18" resultid="4864" heatid="8136" lane="1" entrytime="00:11:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                    <SPLIT distance="100" swimtime="00:01:21.27" />
                    <SPLIT distance="150" swimtime="00:02:04.64" />
                    <SPLIT distance="200" swimtime="00:02:48.33" />
                    <SPLIT distance="250" swimtime="00:03:32.60" />
                    <SPLIT distance="300" swimtime="00:04:17.29" />
                    <SPLIT distance="350" swimtime="00:05:01.68" />
                    <SPLIT distance="400" swimtime="00:05:46.63" />
                    <SPLIT distance="450" swimtime="00:06:31.29" />
                    <SPLIT distance="500" swimtime="00:07:16.46" />
                    <SPLIT distance="550" swimtime="00:08:01.62" />
                    <SPLIT distance="600" swimtime="00:08:46.50" />
                    <SPLIT distance="650" swimtime="00:09:31.75" />
                    <SPLIT distance="700" swimtime="00:10:16.72" />
                    <SPLIT distance="750" swimtime="00:11:01.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="554" reactiontime="+91" swimtime="00:05:46.15" resultid="4865" heatid="8148" lane="5" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.74" />
                    <SPLIT distance="100" swimtime="00:01:22.93" />
                    <SPLIT distance="150" swimtime="00:02:06.89" />
                    <SPLIT distance="200" swimtime="00:02:50.86" />
                    <SPLIT distance="250" swimtime="00:03:34.63" />
                    <SPLIT distance="300" swimtime="00:04:19.36" />
                    <SPLIT distance="350" swimtime="00:05:03.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="613" reactiontime="+78" swimtime="00:00:39.05" resultid="4866" heatid="8106" lane="6" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="4836" name="T.P. Masters Opole">
          <CONTACT name="KRASNODĘBSKI" />
          <ATHLETES>
            <ATHLETE birthdate="1937-01-01" firstname="Tadeusz" gender="M" lastname="Witkowski" nation="POL" athleteid="4842">
              <RESULTS>
                <RESULT eventid="1198" points="417" reactiontime="+121" swimtime="00:01:37.34" resultid="4843" heatid="7982" lane="1" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="295" reactiontime="+100" swimtime="00:04:50.71" resultid="4844" heatid="8023" lane="3" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.58" />
                    <SPLIT distance="100" swimtime="00:02:19.90" />
                    <SPLIT distance="150" swimtime="00:03:36.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="221" reactiontime="+95" swimtime="00:02:27.76" resultid="4845" heatid="8037" lane="9" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="495" reactiontime="+112" swimtime="00:00:39.75" resultid="4846" heatid="8054" lane="9" entrytime="00:00:37.00" />
                <RESULT eventid="1509" points="220" reactiontime="+122" swimtime="00:04:24.47" resultid="4847" heatid="8094" lane="2" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.23" />
                    <SPLIT distance="100" swimtime="00:02:01.81" />
                    <SPLIT distance="150" swimtime="00:03:14.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="396" reactiontime="+93" swimtime="00:00:54.77" resultid="4848" heatid="8110" lane="1" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Jerzy" gender="M" lastname="Minkiewicz" nation="POL" athleteid="4837">
              <RESULTS>
                <RESULT eventid="1198" points="605" reactiontime="+97" swimtime="00:01:11.84" resultid="4838" heatid="7985" lane="2" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="436" reactiontime="+81" swimtime="00:01:34.87" resultid="4839" heatid="8038" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="609" reactiontime="+95" swimtime="00:00:31.39" resultid="4840" heatid="8056" lane="8" entrytime="00:00:32.00" />
                <RESULT eventid="1539" points="502" reactiontime="+77" swimtime="00:00:40.87" resultid="4841" heatid="8111" lane="5" entrytime="00:00:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Zbigniew" gender="M" lastname="Krasnodębski" nation="POL" athleteid="4855">
              <RESULTS>
                <RESULT eventid="1228" points="405" reactiontime="+72" swimtime="00:00:41.96" resultid="4856" heatid="8003" lane="2" entrytime="00:00:42.00" />
                <RESULT eventid="1569" points="425" reactiontime="+65" swimtime="00:01:36.83" resultid="4857" heatid="8128" lane="9" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-01" firstname="Zbigniew" gender="M" lastname="Januszkiewicz" nation="POL" athleteid="4849">
              <RESULTS>
                <RESULT eventid="1198" points="829" reactiontime="+82" swimtime="00:01:01.39" resultid="4850" heatid="7989" lane="3" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="913" reactiontime="+67" swimtime="00:02:33.15" resultid="4851" heatid="8027" lane="5" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.46" />
                    <SPLIT distance="100" swimtime="00:01:15.41" />
                    <SPLIT distance="150" swimtime="00:01:54.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="779" reactiontime="+73" swimtime="00:01:11.55" resultid="4852" heatid="8042" lane="7" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="764" reactiontime="+81" swimtime="00:00:27.78" resultid="4853" heatid="8061" lane="6" entrytime="00:00:28.00" />
                <RESULT eventid="1539" points="826" reactiontime="+66" swimtime="00:00:32.52" resultid="4854" heatid="8115" lane="0" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1318" reactiontime="+83" swimtime="00:05:39.46" resultid="4858" heatid="8030" lane="1" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                    <SPLIT distance="100" swimtime="00:01:06.43" />
                    <SPLIT distance="150" swimtime="00:01:45.15" />
                    <SPLIT distance="200" swimtime="00:02:32.37" />
                    <SPLIT distance="250" swimtime="00:03:22.84" />
                    <SPLIT distance="300" swimtime="00:04:24.22" />
                    <SPLIT distance="350" swimtime="00:04:59.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4849" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="4855" number="2" reactiontime="+63" />
                    <RELAYPOSITION athleteid="4842" number="3" reactiontime="+96" />
                    <RELAYPOSITION athleteid="4837" number="4" reactiontime="+82" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="4731" name="TKKF Koszalin Masters">
          <CONTACT email="jakubkielar3@gmail.com" name="Kielar" phone="693193137" />
          <ATHLETES>
            <ATHLETE birthdate="1972-12-06" firstname="Joanna" gender="F" lastname="Stankiewicz-Majkowska" nation="POL" athleteid="4732">
              <RESULTS>
                <RESULT eventid="1554" points="310" reactiontime="+98" swimtime="00:01:53.39" resultid="4733" heatid="8120" lane="5" entrytime="00:01:43.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1584" points="326" reactiontime="+99" swimtime="00:07:51.16" resultid="4734" heatid="8160" lane="9" entrytime="00:07:57.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.43" />
                    <SPLIT distance="100" swimtime="00:01:52.46" />
                    <SPLIT distance="150" swimtime="00:02:53.16" />
                    <SPLIT distance="200" swimtime="00:03:52.69" />
                    <SPLIT distance="250" swimtime="00:04:55.56" />
                    <SPLIT distance="300" swimtime="00:05:59.27" />
                    <SPLIT distance="350" swimtime="00:06:56.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-07-05" firstname="Krzysztof" gender="M" lastname="Stefański" nation="POL" athleteid="4742">
              <RESULTS>
                <RESULT eventid="1105" points="467" reactiontime="+92" swimtime="00:00:33.37" resultid="4743" heatid="7966" lane="4" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1198" points="565" reactiontime="+81" swimtime="00:01:05.67" resultid="4744" heatid="7988" lane="3" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="626" reactiontime="+76" swimtime="00:00:28.72" resultid="4745" heatid="8061" lane="0" entrytime="00:00:28.00" entrycourse="SCM" />
                <RESULT eventid="1509" points="405" reactiontime="+79" swimtime="00:02:40.09" resultid="4746" heatid="8097" lane="5" entrytime="00:02:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                    <SPLIT distance="100" swimtime="00:01:13.77" />
                    <SPLIT distance="150" swimtime="00:01:56.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" status="DNS" swimtime="00:00:00.00" resultid="4747" heatid="8132" lane="4" entrytime="00:01:00.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-23" firstname="Jarosław" gender="M" lastname="Winiarczyk" nation="POL" athleteid="4748">
              <RESULTS>
                <RESULT eventid="1198" points="566" reactiontime="+81" swimtime="00:01:05.65" resultid="4749" heatid="7988" lane="5" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="597" reactiontime="+75" swimtime="00:00:29.18" resultid="4750" heatid="8061" lane="8" entrytime="00:00:28.00" entrycourse="SCM" />
                <RESULT eventid="1509" points="443" reactiontime="+74" swimtime="00:02:35.39" resultid="4752" heatid="8098" lane="9" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                    <SPLIT distance="100" swimtime="00:01:14.63" />
                    <SPLIT distance="150" swimtime="00:01:55.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-03-02" firstname="Andrzej" gender="M" lastname="Michałkowski" nation="POL" athleteid="4735">
              <RESULTS>
                <RESULT eventid="1198" points="222" reactiontime="+95" swimtime="00:01:40.78" resultid="4736" heatid="7981" lane="5" entrytime="00:01:41.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="502" reactiontime="+101" swimtime="00:00:43.21" resultid="4737" heatid="8004" lane="0" entrytime="00:00:41.80" entrycourse="SCM" />
                <RESULT eventid="1372" points="292" reactiontime="+93" swimtime="00:00:41.15" resultid="4738" heatid="8053" lane="7" entrytime="00:00:39.00" entrycourse="SCM" />
                <RESULT eventid="1402" points="436" reactiontime="+101" swimtime="00:03:55.85" resultid="4739" heatid="8072" lane="6" entrytime="00:03:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.56" />
                    <SPLIT distance="100" swimtime="00:01:49.32" />
                    <SPLIT distance="150" swimtime="00:02:53.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="226" reactiontime="+92" swimtime="00:03:52.41" resultid="4740" heatid="8094" lane="6" entrytime="00:03:47.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.88" />
                    <SPLIT distance="100" swimtime="00:01:47.44" />
                    <SPLIT distance="150" swimtime="00:02:50.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="455" reactiontime="+98" swimtime="00:01:43.12" resultid="4741" heatid="8127" lane="1" entrytime="00:01:38.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02602" nation="POL" region="KUJ" clubid="4753" name="Toruń Multisport Team">
          <CONTACT city="Toruń" email="szufar@o2.pl" name="Szufarski Andrzej" phone="600898866" state="KUJ-P" street="Matejki 60/7" zip="87-100" />
          <ATHLETES>
            <ATHLETE birthdate="1978-03-02" firstname="Maciej" gender="M" lastname="Kuras" nation="POL" athleteid="4791">
              <RESULTS>
                <RESULT eventid="1075" points="472" reactiontime="+81" swimtime="00:02:53.44" resultid="4792" heatid="7950" lane="1" entrytime="00:02:55.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.17" />
                    <SPLIT distance="100" swimtime="00:01:19.87" />
                    <SPLIT distance="150" swimtime="00:02:09.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="512" reactiontime="+77" swimtime="00:00:31.89" resultid="4793" heatid="7967" lane="7" entrytime="00:00:32.55" />
                <RESULT eventid="1288" points="491" reactiontime="+85" swimtime="00:02:49.24" resultid="4794" heatid="8025" lane="3" entrytime="00:02:55.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.79" />
                    <SPLIT distance="100" swimtime="00:01:21.99" />
                    <SPLIT distance="150" swimtime="00:02:05.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="494" reactiontime="+77" swimtime="00:01:18.45" resultid="4795" heatid="8040" lane="3" entrytime="00:01:18.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="449" reactiontime="+82" swimtime="00:01:16.02" resultid="4796" heatid="8084" lane="6" entrytime="00:01:16.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="457" reactiontime="+73" swimtime="00:00:36.60" resultid="4797" heatid="8113" lane="1" entrytime="00:00:35.55" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-23" firstname="Marcin" gender="M" lastname="Mykowski" nation="POL" athleteid="4754">
              <RESULTS>
                <RESULT eventid="1105" points="547" reactiontime="+78" swimtime="00:00:31.19" resultid="4755" heatid="7965" lane="3" entrytime="00:00:35.00" />
                <RESULT eventid="1198" points="635" reactiontime="+80" swimtime="00:01:00.45" resultid="4756" heatid="7985" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="647" reactiontime="+79" swimtime="00:02:34.37" resultid="4757" heatid="8026" lane="6" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.07" />
                    <SPLIT distance="100" swimtime="00:01:17.34" />
                    <SPLIT distance="150" swimtime="00:01:56.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="714" reactiontime="+68" swimtime="00:01:09.39" resultid="4758" heatid="8040" lane="7" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="556" reactiontime="+75" swimtime="00:00:28.61" resultid="4759" heatid="8059" lane="9" entrytime="00:00:29.00" />
                <RESULT eventid="1539" points="707" reactiontime="+69" swimtime="00:00:31.65" resultid="4760" heatid="8113" lane="7" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-10-25" firstname="Katarzyna" gender="F" lastname="Walenta" nation="POL" athleteid="4818">
              <RESULTS>
                <RESULT eventid="1058" points="708" reactiontime="+83" swimtime="00:02:44.49" resultid="4819" heatid="7943" lane="5" entrytime="00:02:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                    <SPLIT distance="100" swimtime="00:01:17.17" />
                    <SPLIT distance="150" swimtime="00:02:04.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="642" reactiontime="+65" swimtime="00:00:33.95" resultid="4820" heatid="7959" lane="9" entrytime="00:00:35.80" />
                <RESULT eventid="1243" points="526" reactiontime="+72" swimtime="00:03:01.70" resultid="4821" heatid="8012" lane="8" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                    <SPLIT distance="100" swimtime="00:01:24.88" />
                    <SPLIT distance="150" swimtime="00:02:13.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1387" points="645" reactiontime="+84" swimtime="00:03:05.58" resultid="4822" heatid="8068" lane="3" entrytime="00:03:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.61" />
                    <SPLIT distance="100" swimtime="00:01:29.07" />
                    <SPLIT distance="150" swimtime="00:02:17.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="598" reactiontime="+85" swimtime="00:01:17.73" resultid="4823" heatid="8079" lane="5" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="619" reactiontime="+78" swimtime="00:01:25.80" resultid="4824" heatid="8122" lane="8" entrytime="00:01:31.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1584" points="628" reactiontime="+92" swimtime="00:06:01.81" resultid="4825" heatid="8159" lane="1" entrytime="00:06:12.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.37" />
                    <SPLIT distance="100" swimtime="00:01:24.43" />
                    <SPLIT distance="150" swimtime="00:02:11.30" />
                    <SPLIT distance="200" swimtime="00:02:56.95" />
                    <SPLIT distance="250" swimtime="00:03:46.04" />
                    <SPLIT distance="300" swimtime="00:04:36.52" />
                    <SPLIT distance="350" swimtime="00:05:20.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-08-24" firstname="Jan" gender="M" lastname="Bantkowski" nation="POL" athleteid="4798">
              <RESULTS>
                <RESULT eventid="1198" points="257" reactiontime="+117" swimtime="00:01:43.75" resultid="4799" heatid="7981" lane="2" entrytime="00:01:48.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="117" reactiontime="+110" swimtime="00:05:28.59" resultid="4800" heatid="8023" lane="0" entrytime="00:04:58.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.24" />
                    <SPLIT distance="100" swimtime="00:02:41.67" />
                    <SPLIT distance="150" swimtime="00:04:06.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="192" reactiontime="+134" swimtime="00:09:16.55" resultid="4801" heatid="8156" lane="3" entrytime="00:08:31.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.66" />
                    <SPLIT distance="100" swimtime="00:02:16.46" />
                    <SPLIT distance="150" swimtime="00:03:29.49" />
                    <SPLIT distance="200" swimtime="00:04:41.39" />
                    <SPLIT distance="250" swimtime="00:05:56.23" />
                    <SPLIT distance="300" swimtime="00:07:07.88" />
                    <SPLIT distance="350" swimtime="00:08:18.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="113" reactiontime="+135" swimtime="00:02:31.20" resultid="4802" heatid="8081" lane="3" entrytime="00:02:23.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="236" reactiontime="+138" swimtime="00:04:03.48" resultid="4803" heatid="8094" lane="1" entrytime="00:03:59.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.83" />
                    <SPLIT distance="100" swimtime="00:01:51.66" />
                    <SPLIT distance="150" swimtime="00:02:56.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="194" reactiontime="+135" swimtime="00:10:51.93" resultid="4804" heatid="8167" lane="8" entrytime="00:10:33.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.09" />
                    <SPLIT distance="100" swimtime="00:02:35.05" />
                    <SPLIT distance="150" swimtime="00:04:07.24" />
                    <SPLIT distance="200" swimtime="00:05:36.22" />
                    <SPLIT distance="250" swimtime="00:07:09.72" />
                    <SPLIT distance="300" swimtime="00:08:38.87" />
                    <SPLIT distance="350" swimtime="00:09:49.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-07-25" firstname="Sławomir" gender="M" lastname="Prędki" nation="POL" athleteid="4826">
              <RESULTS>
                <RESULT eventid="1075" points="882" reactiontime="+77" swimtime="00:02:20.89" resultid="4827" heatid="7946" lane="8" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.95" />
                    <SPLIT distance="100" swimtime="00:01:06.76" />
                    <SPLIT distance="150" swimtime="00:01:47.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="820" reactiontime="+61" swimtime="00:00:27.26" resultid="4828" heatid="7963" lane="9" entrytime="00:00:50.00" />
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1198" points="763" reactiontime="+80" swimtime="00:00:56.87" resultid="4829" heatid="7981" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="744" reactiontime="+71" swimtime="00:00:32.23" resultid="4830" heatid="8000" lane="5" entrytime="00:01:00.00" />
                <RESULT eventid="1402" points="812" reactiontime="+80" swimtime="00:02:42.20" resultid="4831" heatid="8072" lane="0" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.37" />
                    <SPLIT distance="100" swimtime="00:01:16.74" />
                    <SPLIT distance="150" swimtime="00:01:59.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="856" reactiontime="+76" swimtime="00:01:01.31" resultid="4832" heatid="8082" lane="8" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="751" reactiontime="+80" swimtime="00:02:07.24" resultid="4833" heatid="8094" lane="8" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.28" />
                    <SPLIT distance="100" swimtime="00:01:01.94" />
                    <SPLIT distance="150" swimtime="00:01:35.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="805" reactiontime="+78" swimtime="00:01:11.43" resultid="4834" heatid="8124" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-03-07" firstname="Grzegorz" gender="M" lastname="Arentewicz" nation="POL" athleteid="4783">
              <RESULTS>
                <RESULT eventid="1258" points="354" reactiontime="+98" swimtime="00:03:06.98" resultid="4786" heatid="8016" lane="0" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.11" />
                    <SPLIT distance="100" swimtime="00:01:26.15" />
                    <SPLIT distance="150" swimtime="00:02:17.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="425" reactiontime="+88" swimtime="00:01:15.35" resultid="4788" heatid="8083" lane="4" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="374" reactiontime="+85" swimtime="00:02:40.46" resultid="4789" heatid="8096" lane="3" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.82" />
                    <SPLIT distance="100" swimtime="00:01:18.95" />
                    <SPLIT distance="150" swimtime="00:02:00.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="318" reactiontime="+91" swimtime="00:06:40.93" resultid="4790" heatid="8165" lane="4" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.07" />
                    <SPLIT distance="100" swimtime="00:01:23.37" />
                    <SPLIT distance="150" swimtime="00:02:21.43" />
                    <SPLIT distance="200" swimtime="00:03:16.82" />
                    <SPLIT distance="250" swimtime="00:04:14.11" />
                    <SPLIT distance="300" swimtime="00:05:09.63" />
                    <SPLIT distance="350" swimtime="00:05:56.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-02-27" firstname="Magdalena" gender="F" lastname="Rogozińska" nation="POL" athleteid="4774">
              <RESULTS>
                <RESULT eventid="1058" points="464" reactiontime="+89" swimtime="00:03:12.67" resultid="4775" heatid="7942" lane="6" entrytime="00:03:30.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.06" />
                    <SPLIT distance="100" swimtime="00:01:31.05" />
                    <SPLIT distance="150" swimtime="00:02:27.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="401" reactiontime="+95" swimtime="00:00:40.28" resultid="4776" heatid="7956" lane="1" entrytime="00:00:46.10" />
                <RESULT eventid="1181" points="385" reactiontime="+97" swimtime="00:01:22.06" resultid="4777" heatid="7975" lane="8" entrytime="00:01:25.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="475" reactiontime="+87" swimtime="00:00:43.10" resultid="4778" heatid="7996" lane="5" entrytime="00:00:46.30" />
                <RESULT eventid="1357" points="460" reactiontime="+94" swimtime="00:00:35.55" resultid="4779" heatid="8045" lane="3" entrytime="00:00:40.50" />
                <RESULT eventid="1387" points="437" reactiontime="+93" swimtime="00:03:40.24" resultid="4780" heatid="8068" lane="2" entrytime="00:03:40.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.00" />
                    <SPLIT distance="100" swimtime="00:01:49.03" />
                    <SPLIT distance="150" swimtime="00:02:46.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="434" reactiontime="+69" swimtime="00:00:42.38" resultid="4781" heatid="8105" lane="0" entrytime="00:00:46.30" />
                <RESULT eventid="1554" points="424" reactiontime="+90" swimtime="00:01:40.27" resultid="4782" heatid="8121" lane="8" entrytime="00:01:40.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-05-05" firstname="Jarosław" gender="M" lastname="Wysocki" nation="POL" athleteid="4761">
              <RESULTS>
                <RESULT eventid="1075" points="409" reactiontime="+97" swimtime="00:03:38.70" resultid="4762" heatid="7945" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.11" />
                    <SPLIT distance="100" swimtime="00:01:45.50" />
                    <SPLIT distance="150" swimtime="00:02:44.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="391" swimtime="00:03:52.00" resultid="4763" heatid="8013" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.24" />
                    <SPLIT distance="100" swimtime="00:01:42.63" />
                    <SPLIT distance="150" swimtime="00:02:44.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="491" reactiontime="+92" swimtime="00:03:46.71" resultid="4764" heatid="8071" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.67" />
                    <SPLIT distance="100" swimtime="00:01:54.34" />
                    <SPLIT distance="150" swimtime="00:02:53.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="393" reactiontime="+98" swimtime="00:08:01.51" resultid="4765" heatid="8167" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.45" />
                    <SPLIT distance="100" swimtime="00:01:48.15" />
                    <SPLIT distance="150" swimtime="00:02:57.79" />
                    <SPLIT distance="200" swimtime="00:04:03.21" />
                    <SPLIT distance="250" swimtime="00:05:06.32" />
                    <SPLIT distance="300" swimtime="00:06:09.75" />
                    <SPLIT distance="350" swimtime="00:07:07.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-07-06" firstname="Andrzej" gender="M" lastname="Szufarski" nation="POL" athleteid="4812">
              <RESULTS>
                <RESULT eventid="1105" points="328" reactiontime="+100" swimtime="00:00:43.39" resultid="4813" heatid="7963" lane="5" entrytime="00:00:42.00" />
                <RESULT eventid="1228" points="331" reactiontime="+98" swimtime="00:00:49.63" resultid="4814" heatid="8001" lane="6" entrytime="00:00:49.00" />
                <RESULT eventid="1342" points="230" reactiontime="+104" swimtime="00:02:01.74" resultid="4815" heatid="8037" lane="2" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="250" reactiontime="+102" swimtime="00:00:53.24" resultid="4816" heatid="8109" lane="4" entrytime="00:00:49.00" />
                <RESULT eventid="1569" points="311" reactiontime="+101" swimtime="00:01:56.97" resultid="4817" heatid="8125" lane="4" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-04-23" firstname="Krzysztof" gender="M" lastname="Lietz" nation="POL" athleteid="4805">
              <RESULTS>
                <RESULT eventid="1075" points="521" reactiontime="+82" swimtime="00:03:21.73" resultid="4806" heatid="7949" lane="9" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.80" />
                    <SPLIT distance="100" swimtime="00:01:40.15" />
                    <SPLIT distance="150" swimtime="00:02:39.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="531" reactiontime="+86" swimtime="00:00:36.97" resultid="4807" heatid="7965" lane="0" entrytime="00:00:35.50" />
                <RESULT eventid="1198" points="593" reactiontime="+85" swimtime="00:01:12.64" resultid="4808" heatid="7985" lane="7" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="611" reactiontime="+77" swimtime="00:00:32.20" resultid="4809" heatid="8056" lane="2" entrytime="00:00:31.50" />
                <RESULT eventid="1462" points="429" reactiontime="+77" swimtime="00:01:34.89" resultid="4810" heatid="8083" lane="6" entrytime="00:01:27.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="562" reactiontime="+82" swimtime="00:02:51.74" resultid="4811" heatid="8097" lane="3" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.57" />
                    <SPLIT distance="100" swimtime="00:01:24.59" />
                    <SPLIT distance="150" swimtime="00:02:11.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-02-16" firstname="Agnieszka" gender="F" lastname="Kostyra" nation="POL" athleteid="4766">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="4767" heatid="7941" lane="6" />
                <RESULT eventid="1120" status="DNS" swimtime="00:00:00.00" resultid="4768" heatid="8138" lane="4" entrytime="00:13:00.00" />
                <RESULT eventid="1273" points="502" reactiontime="+46" swimtime="00:03:04.70" resultid="4769" heatid="8020" lane="0" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.50" />
                    <SPLIT distance="100" swimtime="00:01:30.80" />
                    <SPLIT distance="150" swimtime="00:02:18.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1387" points="415" reactiontime="+80" swimtime="00:03:28.82" resultid="4770" heatid="8069" lane="9" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.45" />
                    <SPLIT distance="100" swimtime="00:01:40.83" />
                    <SPLIT distance="150" swimtime="00:02:34.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="403" reactiontime="+81" swimtime="00:06:09.25" resultid="4771" heatid="8148" lane="7" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.74" />
                    <SPLIT distance="100" swimtime="00:01:26.37" />
                    <SPLIT distance="150" swimtime="00:02:13.25" />
                    <SPLIT distance="200" swimtime="00:03:01.60" />
                    <SPLIT distance="250" swimtime="00:03:49.88" />
                    <SPLIT distance="300" swimtime="00:04:38.17" />
                    <SPLIT distance="350" swimtime="00:05:26.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="395" reactiontime="+77" swimtime="00:01:38.63" resultid="4772" heatid="8118" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1584" points="431" reactiontime="+80" swimtime="00:06:52.60" resultid="4773" heatid="8160" lane="1" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.34" />
                    <SPLIT distance="100" swimtime="00:01:44.85" />
                    <SPLIT distance="150" swimtime="00:02:37.93" />
                    <SPLIT distance="200" swimtime="00:03:27.80" />
                    <SPLIT distance="250" swimtime="00:04:24.20" />
                    <SPLIT distance="300" swimtime="00:05:21.14" />
                    <SPLIT distance="350" swimtime="00:06:08.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1614" reactiontime="+63" swimtime="00:02:19.96" resultid="4835" heatid="8134" lane="2" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                    <SPLIT distance="100" swimtime="00:01:15.29" />
                    <SPLIT distance="150" swimtime="00:01:48.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4754" number="1" reactiontime="+63" />
                    <RELAYPOSITION athleteid="4774" number="2" />
                    <RELAYPOSITION athleteid="4818" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="4805" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="OLPOZ" nation="POL" region="WIE" clubid="5268" name="TS Olimpia Poznań">
          <CONTACT name="Pietraszewski" phone="501 648 415" />
          <ATHLETES>
            <ATHLETE birthdate="1951-01-01" firstname="Jerzy" gender="M" lastname="Boryski" nation="POL" athleteid="5287">
              <RESULTS>
                <RESULT eventid="1135" points="365" reactiontime="+93" swimtime="00:14:57.96" resultid="5288" heatid="8140" lane="9" entrytime="00:15:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.02" />
                    <SPLIT distance="100" swimtime="00:01:44.73" />
                    <SPLIT distance="150" swimtime="00:02:41.42" />
                    <SPLIT distance="200" swimtime="00:03:39.14" />
                    <SPLIT distance="250" swimtime="00:04:35.57" />
                    <SPLIT distance="300" swimtime="00:05:33.63" />
                    <SPLIT distance="350" swimtime="00:06:30.40" />
                    <SPLIT distance="400" swimtime="00:07:28.05" />
                    <SPLIT distance="450" swimtime="00:08:25.47" />
                    <SPLIT distance="500" swimtime="00:09:22.74" />
                    <SPLIT distance="550" swimtime="00:10:19.65" />
                    <SPLIT distance="600" swimtime="00:11:16.58" />
                    <SPLIT distance="650" swimtime="00:12:13.18" />
                    <SPLIT distance="700" swimtime="00:13:09.89" />
                    <SPLIT distance="750" swimtime="00:14:05.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="461" reactiontime="+78" swimtime="00:01:36.60" resultid="5289" heatid="8038" lane="7" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="537" reactiontime="+80" swimtime="00:00:41.31" resultid="5290" heatid="8111" lane="8" entrytime="00:00:43.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Grażyna" gender="F" lastname="Cabaj-Drela" nation="POL" athleteid="5277">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1090" points="738" reactiontime="+82" swimtime="00:00:38.31" resultid="5278" heatid="7956" lane="3" entrytime="00:00:43.00" />
                <RESULT eventid="1213" points="781" reactiontime="+81" swimtime="00:00:41.63" resultid="5279" heatid="7997" lane="6" entrytime="00:00:43.00" />
                <RESULT eventid="1387" points="774" reactiontime="+85" swimtime="00:03:29.11" resultid="5280" heatid="8069" lane="2" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.01" />
                    <SPLIT distance="100" swimtime="00:01:41.09" />
                    <SPLIT distance="150" swimtime="00:02:35.91" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1554" points="805" reactiontime="+82" swimtime="00:01:31.81" resultid="5281" heatid="8121" lane="5" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Sławomir" gender="M" lastname="Cybertowicz" nation="POL" athleteid="5308">
              <RESULTS>
                <RESULT eventid="1228" status="DNS" swimtime="00:00:00.00" resultid="5309" heatid="8006" lane="5" entrytime="00:00:37.00" />
                <RESULT eventid="1402" points="584" reactiontime="+79" swimtime="00:03:03.89" resultid="5310" heatid="8075" lane="3" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.28" />
                    <SPLIT distance="100" swimtime="00:01:28.36" />
                    <SPLIT distance="150" swimtime="00:02:16.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="587" reactiontime="+74" swimtime="00:01:22.30" resultid="5311" heatid="8130" lane="3" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Andrzej" gender="M" lastname="Sypniewski" nation="POL" athleteid="5299">
              <RESULTS>
                <RESULT eventid="1075" points="475" reactiontime="+110" swimtime="00:03:18.68" resultid="5300" heatid="7948" lane="0" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.55" />
                    <SPLIT distance="100" swimtime="00:01:36.61" />
                    <SPLIT distance="150" swimtime="00:02:31.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="443" reactiontime="+108" swimtime="00:00:37.42" resultid="5301" heatid="7964" lane="2" entrytime="00:00:36.80" />
                <RESULT eventid="1198" points="494" reactiontime="+88" swimtime="00:01:16.83" resultid="5302" heatid="7984" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="359" reactiontime="+83" swimtime="00:00:43.66" resultid="5303" heatid="8004" lane="6" entrytime="00:00:40.15" />
                <RESULT eventid="1342" points="409" reactiontime="+77" swimtime="00:01:36.94" resultid="5304" heatid="8038" lane="6" entrytime="00:01:32.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="514" reactiontime="+87" swimtime="00:00:33.20" resultid="5305" heatid="8055" lane="5" entrytime="00:00:32.16" />
                <RESULT eventid="1539" points="498" reactiontime="+86" swimtime="00:00:40.99" resultid="5306" heatid="8112" lane="9" entrytime="00:00:40.28" />
                <RESULT eventid="1569" points="445" reactiontime="+103" swimtime="00:01:35.37" resultid="5307" heatid="8128" lane="7" entrytime="00:01:30.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Zbigniew" gender="M" lastname="Pietraszewski" nation="POL" athleteid="5291">
              <RESULTS>
                <RESULT eventid="1075" points="597" reactiontime="+94" swimtime="00:03:12.78" resultid="5292" heatid="7949" lane="7" entrytime="00:03:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.39" />
                    <SPLIT distance="100" swimtime="00:01:35.66" />
                    <SPLIT distance="150" swimtime="00:02:28.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="565" reactiontime="+91" swimtime="00:00:41.53" resultid="5293" heatid="8003" lane="3" entrytime="00:00:42.00" />
                <RESULT eventid="1288" points="693" reactiontime="+77" swimtime="00:03:11.22" resultid="5294" heatid="8024" lane="4" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.60" />
                    <SPLIT distance="100" swimtime="00:01:32.33" />
                    <SPLIT distance="150" swimtime="00:02:22.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="575" reactiontime="+82" swimtime="00:01:29.73" resultid="5295" heatid="8039" lane="0" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="536" reactiontime="+94" swimtime="00:06:21.01" resultid="5296" heatid="8154" lane="1" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.31" />
                    <SPLIT distance="100" swimtime="00:01:29.77" />
                    <SPLIT distance="150" swimtime="00:02:18.88" />
                    <SPLIT distance="200" swimtime="00:03:08.24" />
                    <SPLIT distance="250" swimtime="00:03:57.34" />
                    <SPLIT distance="300" swimtime="00:04:46.54" />
                    <SPLIT distance="350" swimtime="00:05:34.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="504" reactiontime="+75" swimtime="00:00:42.17" resultid="5297" heatid="8111" lane="4" entrytime="00:00:41.00" />
                <RESULT eventid="1599" points="609" reactiontime="+88" swimtime="00:06:56.05" resultid="5298" heatid="8164" lane="9" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.13" />
                    <SPLIT distance="100" swimtime="00:01:46.98" />
                    <SPLIT distance="150" swimtime="00:02:38.59" />
                    <SPLIT distance="200" swimtime="00:03:30.44" />
                    <SPLIT distance="250" swimtime="00:04:25.97" />
                    <SPLIT distance="300" swimtime="00:05:22.37" />
                    <SPLIT distance="350" swimtime="00:06:11.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Anna" gender="F" lastname="Gano-Kosturkiewicz" nation="POL" athleteid="5282">
              <RESULTS>
                <RESULT eventid="1090" points="349" reactiontime="+118" swimtime="00:00:49.17" resultid="5283" heatid="7956" lane="0" entrytime="00:00:47.00" />
                <RESULT eventid="1181" points="274" reactiontime="+130" swimtime="00:01:46.40" resultid="5284" heatid="7974" lane="0" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="360" reactiontime="+108" swimtime="00:00:43.40" resultid="5285" heatid="8045" lane="2" entrytime="00:00:43.00" />
                <RESULT eventid="1524" points="263" reactiontime="+88" swimtime="00:00:56.80" resultid="5286" heatid="8104" lane="6" entrytime="00:00:53.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Maria" gender="F" lastname="Łutowicz" nation="POL" athleteid="5269">
              <RESULTS>
                <RESULT eventid="1090" points="376" reactiontime="+93" swimtime="00:00:49.52" resultid="5270" heatid="7955" lane="2" entrytime="00:00:53.00" />
                <RESULT eventid="1181" points="505" reactiontime="+98" swimtime="00:01:30.39" resultid="5271" heatid="7974" lane="2" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="533" reactiontime="+96" swimtime="00:00:51.18" resultid="5272" heatid="7995" lane="3" entrytime="00:00:53.00" />
                <RESULT eventid="1357" points="597" reactiontime="+88" swimtime="00:00:38.61" resultid="5273" heatid="8046" lane="9" entrytime="00:00:39.00" />
                <RESULT comment="Rekord Polski Masters" eventid="1417" points="580" reactiontime="+100" swimtime="00:07:12.35" resultid="5274" heatid="8149" lane="3" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.08" />
                    <SPLIT distance="100" swimtime="00:01:42.62" />
                    <SPLIT distance="150" swimtime="00:02:40.60" />
                    <SPLIT distance="200" swimtime="00:03:36.40" />
                    <SPLIT distance="250" swimtime="00:04:30.62" />
                    <SPLIT distance="300" swimtime="00:05:25.28" />
                    <SPLIT distance="350" swimtime="00:06:20.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="502" reactiontime="+84" swimtime="00:03:24.07" resultid="5275" heatid="8088" lane="1" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.81" />
                    <SPLIT distance="100" swimtime="00:01:37.09" />
                    <SPLIT distance="150" swimtime="00:02:32.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="543" reactiontime="+73" swimtime="00:00:49.81" resultid="5276" heatid="8104" lane="4" entrytime="00:00:49.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-01" firstname="Bartłomiej" gender="M" lastname="Zadorożny" nation="POL" athleteid="5312">
              <RESULTS>
                <RESULT eventid="1105" points="559" reactiontime="+74" swimtime="00:00:30.98" resultid="5313" heatid="7967" lane="2" entrytime="00:00:32.51" />
                <RESULT eventid="1198" points="499" reactiontime="+126" swimtime="00:01:05.53" resultid="5314" heatid="7989" lane="8" entrytime="00:01:04.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="552" swimtime="00:00:35.59" resultid="5315" heatid="8007" lane="5" entrytime="00:00:35.71" />
                <RESULT eventid="1372" points="586" reactiontime="+68" swimtime="00:00:28.11" resultid="5316" heatid="8059" lane="4" entrytime="00:00:28.82" />
                <RESULT eventid="1402" points="620" reactiontime="+88" swimtime="00:02:57.49" resultid="5317" heatid="8076" lane="8" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.86" />
                    <SPLIT distance="100" swimtime="00:01:25.12" />
                    <SPLIT distance="150" swimtime="00:02:11.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="586" reactiontime="+72" swimtime="00:01:19.40" resultid="5318" heatid="8130" lane="7" entrytime="00:01:21.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1614" reactiontime="+87" swimtime="00:02:29.60" resultid="5319" heatid="8133" lane="5" entrytime="00:02:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.32" />
                    <SPLIT distance="100" swimtime="00:01:18.22" />
                    <SPLIT distance="150" swimtime="00:01:50.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5277" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="5308" number="2" />
                    <RELAYPOSITION athleteid="5312" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="5269" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00408" nation="POL" region="RZ" clubid="4867" name="Uks Delfin Masters Tarnobrzeg">
          <CONTACT city="TARNOBRZEG" email="piotr.michalik@i-bs.pl" name="MICHALIK ANGELIKA" state="PODKA" street="SKALNA GÓRA 8/21" street2="TARNOBRZEG" zip="39-400" />
          <ATHLETES>
            <ATHLETE birthdate="1977-04-24" firstname="Renata" gender="F" lastname="Osmala" nation="POL" athleteid="4868">
              <RESULTS>
                <RESULT eventid="1120" points="687" reactiontime="+82" swimtime="00:10:59.18" resultid="4869" heatid="8136" lane="7" entrytime="00:11:27.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                    <SPLIT distance="100" swimtime="00:01:15.95" />
                    <SPLIT distance="150" swimtime="00:01:56.94" />
                    <SPLIT distance="200" swimtime="00:02:38.23" />
                    <SPLIT distance="250" swimtime="00:03:19.56" />
                    <SPLIT distance="300" swimtime="00:04:01.31" />
                    <SPLIT distance="350" swimtime="00:04:43.17" />
                    <SPLIT distance="400" swimtime="00:05:25.49" />
                    <SPLIT distance="450" swimtime="00:06:07.33" />
                    <SPLIT distance="500" swimtime="00:06:49.30" />
                    <SPLIT distance="550" swimtime="00:07:31.36" />
                    <SPLIT distance="600" swimtime="00:08:13.87" />
                    <SPLIT distance="650" swimtime="00:08:55.86" />
                    <SPLIT distance="700" swimtime="00:09:38.03" />
                    <SPLIT distance="750" swimtime="00:10:19.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="539" swimtime="00:00:41.32" resultid="4870" heatid="7998" lane="8" entrytime="00:00:41.50" />
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1273" points="667" reactiontime="+77" swimtime="00:02:50.41" resultid="4871" heatid="8020" lane="4" entrytime="00:02:54.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.29" />
                    <SPLIT distance="100" swimtime="00:01:23.14" />
                    <SPLIT distance="150" swimtime="00:02:06.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="636" reactiontime="+75" swimtime="00:01:21.22" resultid="4872" heatid="8034" lane="6" entrytime="00:01:24.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="696" reactiontime="+83" swimtime="00:05:20.79" resultid="4873" heatid="8147" lane="1" entrytime="00:05:25.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                    <SPLIT distance="100" swimtime="00:01:15.87" />
                    <SPLIT distance="150" swimtime="00:01:56.80" />
                    <SPLIT distance="200" swimtime="00:02:37.93" />
                    <SPLIT distance="250" swimtime="00:03:18.93" />
                    <SPLIT distance="300" swimtime="00:04:00.40" />
                    <SPLIT distance="350" swimtime="00:04:41.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="590" reactiontime="+74" swimtime="00:00:38.28" resultid="4874" heatid="8106" lane="8" entrytime="00:00:39.09" />
                <RESULT eventid="1554" points="562" reactiontime="+79" swimtime="00:01:31.30" resultid="4875" heatid="8122" lane="1" entrytime="00:01:31.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-23" firstname="Krzysztof" gender="M" lastname="Ślęczka" nation="POL" athleteid="4919">
              <RESULTS>
                <RESULT eventid="1105" points="647" reactiontime="+80" swimtime="00:00:29.94" resultid="4920" heatid="7967" lane="1" entrytime="00:00:32.68" />
                <RESULT eventid="1135" points="542" reactiontime="+88" swimtime="00:10:45.51" resultid="4921" heatid="8139" lane="8" entrytime="00:11:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                    <SPLIT distance="100" swimtime="00:01:12.33" />
                    <SPLIT distance="150" swimtime="00:01:52.56" />
                    <SPLIT distance="200" swimtime="00:02:33.55" />
                    <SPLIT distance="250" swimtime="00:03:14.60" />
                    <SPLIT distance="300" swimtime="00:03:56.08" />
                    <SPLIT distance="350" swimtime="00:04:37.61" />
                    <SPLIT distance="400" swimtime="00:05:18.73" />
                    <SPLIT distance="450" swimtime="00:06:00.54" />
                    <SPLIT distance="500" swimtime="00:06:42.39" />
                    <SPLIT distance="550" swimtime="00:07:24.34" />
                    <SPLIT distance="600" swimtime="00:08:05.91" />
                    <SPLIT distance="650" swimtime="00:08:47.45" />
                    <SPLIT distance="700" swimtime="00:09:29.30" />
                    <SPLIT distance="750" swimtime="00:10:09.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="767" reactiontime="+78" swimtime="00:00:59.32" resultid="4922" heatid="7990" lane="9" entrytime="00:01:02.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="701" swimtime="00:00:34.33" resultid="4923" heatid="8007" lane="8" entrytime="00:00:36.89" />
                <RESULT eventid="1372" points="751" reactiontime="+82" swimtime="00:00:27.04" resultid="4924" heatid="8059" lane="5" entrytime="00:00:28.84" />
                <RESULT eventid="1432" points="591" reactiontime="+83" swimtime="00:05:03.10" resultid="4925" heatid="8152" lane="6" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                    <SPLIT distance="100" swimtime="00:01:10.77" />
                    <SPLIT distance="150" swimtime="00:01:49.64" />
                    <SPLIT distance="200" swimtime="00:02:29.81" />
                    <SPLIT distance="250" swimtime="00:03:09.54" />
                    <SPLIT distance="300" swimtime="00:03:49.40" />
                    <SPLIT distance="350" swimtime="00:04:27.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="688" reactiontime="+79" swimtime="00:02:14.18" resultid="4926" heatid="8100" lane="2" entrytime="00:02:22.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.95" />
                    <SPLIT distance="100" swimtime="00:01:03.75" />
                    <SPLIT distance="150" swimtime="00:01:38.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="657" reactiontime="+82" swimtime="00:01:19.03" resultid="4927" heatid="8130" lane="8" entrytime="00:01:22.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-03-30" firstname="Angelika" gender="F" lastname="Rozmus" nation="POL" athleteid="4876">
              <RESULTS>
                <RESULT eventid="1058" points="538" reactiontime="+84" swimtime="00:03:03.40" resultid="4877" heatid="7942" lane="2" entrytime="00:03:30.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.40" />
                    <SPLIT distance="100" swimtime="00:01:27.74" />
                    <SPLIT distance="150" swimtime="00:02:20.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="487" reactiontime="+87" swimtime="00:00:37.74" resultid="4878" heatid="7957" lane="6" entrytime="00:00:38.20" />
                <RESULT eventid="1181" points="528" reactiontime="+80" swimtime="00:01:13.84" resultid="4879" heatid="7977" lane="5" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="464" swimtime="00:00:43.44" resultid="4880" heatid="7998" lane="3" entrytime="00:00:41.00" />
                <RESULT eventid="1357" points="546" reactiontime="+80" swimtime="00:00:33.57" resultid="4881" heatid="8047" lane="5" entrytime="00:00:33.50" />
                <RESULT eventid="1447" points="393" reactiontime="+84" swimtime="00:01:30.97" resultid="4882" heatid="8079" lane="2" entrytime="00:01:27.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="492" reactiontime="+83" swimtime="00:00:40.65" resultid="4883" heatid="8106" lane="9" entrytime="00:00:39.30" />
                <RESULT eventid="1554" points="494" reactiontime="+76" swimtime="00:01:35.29" resultid="4884" heatid="8121" lane="4" entrytime="00:01:33.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-04-09" firstname="Zbigniew" gender="M" lastname="Ramos" nation="POL" athleteid="4899">
              <RESULTS>
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="4900" heatid="7967" lane="0" entrytime="00:00:33.00" />
                <RESULT eventid="1198" points="541" reactiontime="+85" swimtime="00:01:08.53" resultid="4901" heatid="7986" lane="1" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="469" reactiontime="+85" swimtime="00:00:38.47" resultid="4902" heatid="8005" lane="4" entrytime="00:00:38.00" />
                <RESULT eventid="1372" status="DNS" swimtime="00:00:00.00" resultid="4903" heatid="8057" lane="8" entrytime="00:00:30.00" />
                <RESULT eventid="1402" points="473" reactiontime="+97" swimtime="00:03:17.25" resultid="4904" heatid="8074" lane="6" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.73" />
                    <SPLIT distance="100" swimtime="00:01:34.54" />
                    <SPLIT distance="150" swimtime="00:02:27.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="526" reactiontime="+87" swimtime="00:01:25.33" resultid="4905" heatid="8129" lane="5" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-17" firstname="Sławomir" gender="M" lastname="Kowalski" nation="POL" athleteid="4912">
              <RESULTS>
                <RESULT eventid="1075" points="569" reactiontime="+79" swimtime="00:02:39.78" resultid="4913" heatid="7951" lane="1" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                    <SPLIT distance="100" swimtime="00:01:17.10" />
                    <SPLIT distance="150" swimtime="00:02:01.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="565" reactiontime="+73" swimtime="00:00:31.32" resultid="4914" heatid="7966" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="1228" points="676" reactiontime="+72" swimtime="00:00:34.75" resultid="4915" heatid="8008" lane="6" entrytime="00:00:34.00" />
                <RESULT eventid="1372" points="435" reactiontime="+78" swimtime="00:00:32.42" resultid="4916" heatid="8055" lane="1" entrytime="00:00:33.00" />
                <RESULT eventid="1402" points="618" reactiontime="+72" swimtime="00:02:57.11" resultid="4917" heatid="8076" lane="0" entrytime="00:02:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                    <SPLIT distance="100" swimtime="00:01:24.99" />
                    <SPLIT distance="150" swimtime="00:02:11.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="670" reactiontime="+65" swimtime="00:01:18.53" resultid="4918" heatid="8131" lane="9" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-12" firstname="Maciej" gender="M" lastname="Płaneta" nation="POL" athleteid="4885">
              <RESULTS>
                <RESULT eventid="1105" points="411" reactiontime="+73" swimtime="00:00:34.82" resultid="4886" heatid="7966" lane="7" entrytime="00:00:34.00" />
                <RESULT eventid="1165" points="398" reactiontime="+80" swimtime="00:22:46.77" resultid="4887" heatid="8144" lane="3" entrytime="00:22:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.37" />
                    <SPLIT distance="100" swimtime="00:01:22.41" />
                    <SPLIT distance="150" swimtime="00:02:07.24" />
                    <SPLIT distance="200" swimtime="00:02:52.34" />
                    <SPLIT distance="250" swimtime="00:03:37.42" />
                    <SPLIT distance="300" swimtime="00:04:23.15" />
                    <SPLIT distance="350" swimtime="00:05:08.61" />
                    <SPLIT distance="400" swimtime="00:05:54.36" />
                    <SPLIT distance="450" swimtime="00:06:40.25" />
                    <SPLIT distance="500" swimtime="00:07:26.21" />
                    <SPLIT distance="550" swimtime="00:08:11.67" />
                    <SPLIT distance="600" swimtime="00:08:57.56" />
                    <SPLIT distance="650" swimtime="00:09:43.48" />
                    <SPLIT distance="700" swimtime="00:10:29.14" />
                    <SPLIT distance="750" swimtime="00:11:15.21" />
                    <SPLIT distance="800" swimtime="00:12:01.14" />
                    <SPLIT distance="850" swimtime="00:12:47.33" />
                    <SPLIT distance="900" swimtime="00:13:33.20" />
                    <SPLIT distance="950" swimtime="00:14:19.63" />
                    <SPLIT distance="1000" swimtime="00:15:05.03" />
                    <SPLIT distance="1050" swimtime="00:15:50.58" />
                    <SPLIT distance="1100" swimtime="00:16:36.30" />
                    <SPLIT distance="1150" swimtime="00:17:22.83" />
                    <SPLIT distance="1200" swimtime="00:18:09.57" />
                    <SPLIT distance="1250" swimtime="00:18:56.48" />
                    <SPLIT distance="1300" swimtime="00:19:43.19" />
                    <SPLIT distance="1350" swimtime="00:20:30.59" />
                    <SPLIT distance="1400" swimtime="00:21:18.01" />
                    <SPLIT distance="1450" swimtime="00:22:04.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="476" reactiontime="+81" swimtime="00:01:09.57" resultid="4888" heatid="7987" lane="1" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="504" reactiontime="+79" swimtime="00:00:30.88" resultid="4889" heatid="8057" lane="4" entrytime="00:00:30.00" />
                <RESULT eventid="1432" points="420" reactiontime="+70" swimtime="00:05:39.47" resultid="4890" heatid="8152" lane="9" entrytime="00:05:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.19" />
                    <SPLIT distance="100" swimtime="00:01:16.77" />
                    <SPLIT distance="150" swimtime="00:02:00.47" />
                    <SPLIT distance="200" swimtime="00:02:44.70" />
                    <SPLIT distance="250" swimtime="00:03:29.75" />
                    <SPLIT distance="300" swimtime="00:04:14.26" />
                    <SPLIT distance="350" swimtime="00:04:58.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="448" reactiontime="+79" swimtime="00:02:34.80" resultid="4891" heatid="8099" lane="5" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                    <SPLIT distance="100" swimtime="00:01:11.82" />
                    <SPLIT distance="150" swimtime="00:01:52.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="360" reactiontime="+82" swimtime="00:06:37.56" resultid="4892" heatid="8163" lane="1" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.29" />
                    <SPLIT distance="100" swimtime="00:01:32.11" />
                    <SPLIT distance="150" swimtime="00:02:26.93" />
                    <SPLIT distance="200" swimtime="00:03:19.22" />
                    <SPLIT distance="250" swimtime="00:04:16.67" />
                    <SPLIT distance="300" swimtime="00:05:13.48" />
                    <SPLIT distance="350" swimtime="00:05:56.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-25" firstname="Artur" gender="M" lastname="Szklarz" nation="POL" athleteid="4893">
              <RESULTS>
                <RESULT eventid="1105" points="475" reactiontime="+75" swimtime="00:00:33.19" resultid="4894" heatid="7967" lane="6" entrytime="00:00:32.50" />
                <RESULT eventid="1228" points="520" reactiontime="+77" swimtime="00:00:37.94" resultid="4895" heatid="8006" lane="6" entrytime="00:00:37.00" />
                <RESULT eventid="1372" points="542" reactiontime="+74" swimtime="00:00:30.13" resultid="4896" heatid="8058" lane="2" entrytime="00:00:29.50" />
                <RESULT eventid="1462" points="364" reactiontime="+78" swimtime="00:01:22.13" resultid="4897" heatid="8084" lane="5" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="455" reactiontime="+68" swimtime="00:00:37.04" resultid="4898" heatid="8113" lane="9" entrytime="00:00:36.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-03-28" firstname="Agata" gender="F" lastname="Meksuła" nation="POL" athleteid="4906">
              <RESULTS>
                <RESULT eventid="1090" points="533" reactiontime="+63" swimtime="00:00:36.64" resultid="4907" heatid="7958" lane="8" entrytime="00:00:37.15" />
                <RESULT eventid="1181" points="559" reactiontime="+88" swimtime="00:01:12.45" resultid="4908" heatid="7978" lane="7" entrytime="00:01:10.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="619" reactiontime="+90" swimtime="00:00:32.20" resultid="4909" heatid="8048" lane="7" entrytime="00:00:32.05" />
                <RESULT eventid="1493" points="541" reactiontime="+84" swimtime="00:02:42.47" resultid="4910" heatid="8091" lane="8" entrytime="00:02:40.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                    <SPLIT distance="100" swimtime="00:01:19.34" />
                    <SPLIT distance="150" swimtime="00:02:01.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="523" reactiontime="+70" swimtime="00:00:39.84" resultid="4911" heatid="8106" lane="1" entrytime="00:00:39.06" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1318" status="DNS" swimtime="00:00:00.00" resultid="4929" heatid="8031" lane="0" entrytime="00:04:12.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4919" number="1" />
                    <RELAYPOSITION athleteid="4912" number="2" />
                    <RELAYPOSITION athleteid="4893" number="3" />
                    <RELAYPOSITION athleteid="4899" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1318" reactiontime="+81" swimtime="00:04:15.43" resultid="6171" heatid="8031" lane="1" entrytime="00:04:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.82" />
                    <SPLIT distance="100" swimtime="00:00:59.38" />
                    <SPLIT distance="150" swimtime="00:01:29.10" />
                    <SPLIT distance="200" swimtime="00:02:03.74" />
                    <SPLIT distance="250" swimtime="00:02:34.32" />
                    <SPLIT distance="300" swimtime="00:03:08.69" />
                    <SPLIT distance="350" swimtime="00:03:39.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4919" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="4912" number="2" reactiontime="+24" />
                    <RELAYPOSITION athleteid="4893" number="3" reactiontime="+32" />
                    <RELAYPOSITION athleteid="4899" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1614" reactiontime="+79" swimtime="00:02:14.21" resultid="6170" heatid="8134" lane="4" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                    <SPLIT distance="100" swimtime="00:01:13.48" />
                    <SPLIT distance="150" swimtime="00:01:42.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4868" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="4912" number="2" />
                    <RELAYPOSITION athleteid="4919" number="3" reactiontime="+60" />
                    <RELAYPOSITION athleteid="4906" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="00501" nation="POL" region="DOL" clubid="4967" name="UKS Energetyk Zgorzelec">
          <CONTACT city="Zgorzelec" email="biuro@plywanie-zgorzelec.pl" internet="www. plywanie-zgorzelec.pl" name="Daszyński" phone="607151541" state="DOL" zip="59-900" />
          <ATHLETES>
            <ATHLETE birthdate="1948-11-29" firstname="Andrzej" gender="M" lastname="Daszyński" nation="POL" athleteid="4968">
              <RESULTS>
                <RESULT eventid="1075" points="287" reactiontime="+88" swimtime="00:04:10.96" resultid="4969" heatid="7946" lane="7" entrytime="00:03:59.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.89" />
                    <SPLIT distance="100" swimtime="00:02:01.03" />
                    <SPLIT distance="150" swimtime="00:03:16.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="308" swimtime="00:16:10.58" resultid="4970" heatid="8141" lane="5" entrytime="00:17:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.57" />
                    <SPLIT distance="100" swimtime="00:01:52.08" />
                    <SPLIT distance="150" swimtime="00:02:54.50" />
                    <SPLIT distance="200" swimtime="00:03:56.22" />
                    <SPLIT distance="250" swimtime="00:04:59.32" />
                    <SPLIT distance="300" swimtime="00:06:02.41" />
                    <SPLIT distance="350" swimtime="00:07:05.90" />
                    <SPLIT distance="400" swimtime="00:08:07.89" />
                    <SPLIT distance="450" swimtime="00:09:08.01" />
                    <SPLIT distance="500" swimtime="00:10:09.36" />
                    <SPLIT distance="550" swimtime="00:11:10.84" />
                    <SPLIT distance="600" swimtime="00:12:13.78" />
                    <SPLIT distance="650" swimtime="00:13:13.54" />
                    <SPLIT distance="700" swimtime="00:14:14.73" />
                    <SPLIT distance="750" swimtime="00:15:15.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="235" reactiontime="+90" swimtime="00:04:44.85" resultid="4971" heatid="8014" lane="2" entrytime="00:04:36.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.46" />
                    <SPLIT distance="100" swimtime="00:02:17.80" />
                    <SPLIT distance="150" swimtime="00:03:32.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="304" reactiontime="+74" swimtime="00:03:59.13" resultid="4972" heatid="8024" lane="8" entrytime="00:03:55.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.39" />
                    <SPLIT distance="100" swimtime="00:01:59.02" />
                    <SPLIT distance="150" swimtime="00:03:01.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="275" reactiontime="+73" swimtime="00:01:53.41" resultid="4973" heatid="8038" lane="9" entrytime="00:01:50.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="191" swimtime="00:02:06.76" resultid="4974" heatid="8082" lane="9" entrytime="00:02:02.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="302" reactiontime="+76" swimtime="00:00:49.93" resultid="4975" heatid="8109" lane="5" entrytime="00:00:49.00" />
                <RESULT eventid="1599" points="368" reactiontime="+89" swimtime="00:08:46.28" resultid="4976" heatid="8167" lane="5" entrytime="00:08:42.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.83" />
                    <SPLIT distance="100" swimtime="00:02:10.32" />
                    <SPLIT distance="150" swimtime="00:03:18.01" />
                    <SPLIT distance="200" swimtime="00:04:21.56" />
                    <SPLIT distance="250" swimtime="00:05:38.66" />
                    <SPLIT distance="300" swimtime="00:06:51.85" />
                    <SPLIT distance="350" swimtime="00:07:48.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="02214" nation="POL" clubid="4930" name="UKS JAGIELLONKA Warszawa">
          <CONTACT email="klipson@op.pl" name="Klepko" />
          <ATHLETES>
            <ATHLETE birthdate="1982-06-03" firstname="Piotr" gender="M" lastname="Fuliński" nation="POL" athleteid="4933">
              <RESULTS>
                <RESULT eventid="1198" points="654" reactiontime="+83" swimtime="00:00:58.56" resultid="4934" heatid="7993" lane="1" entrytime="00:00:57.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="671" reactiontime="+83" swimtime="00:00:26.55" resultid="4935" heatid="8064" lane="1" entrytime="00:00:26.10" />
                <RESULT eventid="1509" points="614" reactiontime="+87" swimtime="00:02:16.10" resultid="4936" heatid="8102" lane="7" entrytime="00:02:10.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.51" />
                    <SPLIT distance="100" swimtime="00:01:05.60" />
                    <SPLIT distance="150" swimtime="00:01:41.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WODKAT" nation="POL" region="SLA" clubid="4937" name="UKS Wodnik 29 Katowice">
          <CONTACT email="skoczyt@gmail.com" name="Skoczylas Tomasz" phone="662297707" />
          <ATHLETES>
            <ATHLETE birthdate="1940-07-09" firstname="Krystyna" gender="F" lastname="Nicpoń" nation="POL" athleteid="4953">
              <RESULTS>
                <RESULT eventid="1090" points="177" reactiontime="+98" swimtime="00:01:27.20" resultid="4954" heatid="7955" lane="9" entrytime="00:01:45.00" />
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1120" points="441" swimtime="00:18:20.93" resultid="4955" heatid="8138" lane="3" entrytime="00:20:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.55" />
                    <SPLIT distance="100" swimtime="00:02:03.59" />
                    <SPLIT distance="150" swimtime="00:03:11.51" />
                    <SPLIT distance="200" swimtime="00:04:19.93" />
                    <SPLIT distance="250" swimtime="00:05:29.42" />
                    <SPLIT distance="300" swimtime="00:06:40.27" />
                    <SPLIT distance="350" swimtime="00:07:50.17" />
                    <SPLIT distance="400" swimtime="00:08:58.31" />
                    <SPLIT distance="450" swimtime="00:10:09.69" />
                    <SPLIT distance="500" swimtime="00:11:20.53" />
                    <SPLIT distance="550" swimtime="00:12:31.92" />
                    <SPLIT distance="600" swimtime="00:13:42.39" />
                    <SPLIT distance="650" swimtime="00:14:53.57" />
                    <SPLIT distance="700" swimtime="00:16:03.22" />
                    <SPLIT distance="750" swimtime="00:17:12.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="495" reactiontime="+102" swimtime="00:01:55.94" resultid="4956" heatid="7973" lane="3" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.41" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1273" points="884" reactiontime="+77" swimtime="00:04:10.82" resultid="4957" heatid="8018" lane="5" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.27" />
                    <SPLIT distance="100" swimtime="00:02:00.03" />
                    <SPLIT distance="150" swimtime="00:03:05.86" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1326" points="719" reactiontime="+84" swimtime="00:02:01.08" resultid="4958" heatid="8032" lane="5" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.91" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1417" points="460" reactiontime="+79" swimtime="00:08:46.41" resultid="4959" heatid="8150" lane="5" entrytime="00:10:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.76" />
                    <SPLIT distance="100" swimtime="00:02:00.80" />
                    <SPLIT distance="150" swimtime="00:03:08.68" />
                    <SPLIT distance="200" swimtime="00:04:17.37" />
                    <SPLIT distance="250" swimtime="00:05:25.75" />
                    <SPLIT distance="300" swimtime="00:06:33.20" />
                    <SPLIT distance="350" swimtime="00:07:41.19" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1524" points="659" reactiontime="+84" swimtime="00:00:52.86" resultid="4960" heatid="8104" lane="0" entrytime="00:01:00.00" />
                <RESULT comment="Rekord Polski Masters" eventid="1584" points="442" reactiontime="+93" swimtime="00:10:41.27" resultid="4961" heatid="8161" lane="6" entrytime="00:15:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:33.97" />
                    <SPLIT distance="100" swimtime="00:03:23.23" />
                    <SPLIT distance="150" swimtime="00:04:25.86" />
                    <SPLIT distance="200" swimtime="00:05:31.69" />
                    <SPLIT distance="250" swimtime="00:06:57.23" />
                    <SPLIT distance="300" swimtime="00:08:22.23" />
                    <SPLIT distance="350" swimtime="00:09:30.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-04-22" firstname="Tomasz" gender="M" lastname="Skoczylas" nation="POL" athleteid="4938">
              <RESULTS>
                <RESULT eventid="1105" points="438" reactiontime="+84" swimtime="00:00:35.84" resultid="4939" heatid="7966" lane="9" entrytime="00:00:34.50" />
                <RESULT eventid="1165" points="483" reactiontime="+102" swimtime="00:21:54.31" resultid="4940" heatid="8143" lane="0" entrytime="00:21:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                    <SPLIT distance="100" swimtime="00:01:17.30" />
                    <SPLIT distance="150" swimtime="00:01:59.20" />
                    <SPLIT distance="200" swimtime="00:02:42.78" />
                    <SPLIT distance="250" swimtime="00:03:25.35" />
                    <SPLIT distance="300" swimtime="00:04:08.73" />
                    <SPLIT distance="350" swimtime="00:04:51.84" />
                    <SPLIT distance="400" swimtime="00:05:35.51" />
                    <SPLIT distance="450" swimtime="00:06:19.13" />
                    <SPLIT distance="500" swimtime="00:07:03.50" />
                    <SPLIT distance="550" swimtime="00:07:47.35" />
                    <SPLIT distance="600" swimtime="00:08:31.62" />
                    <SPLIT distance="650" swimtime="00:09:15.56" />
                    <SPLIT distance="700" swimtime="00:09:59.72" />
                    <SPLIT distance="750" swimtime="00:10:43.95" />
                    <SPLIT distance="800" swimtime="00:11:28.81" />
                    <SPLIT distance="850" swimtime="00:12:13.70" />
                    <SPLIT distance="900" swimtime="00:12:58.54" />
                    <SPLIT distance="950" swimtime="00:13:43.15" />
                    <SPLIT distance="1000" swimtime="00:14:28.08" />
                    <SPLIT distance="1050" swimtime="00:15:12.89" />
                    <SPLIT distance="1100" swimtime="00:15:57.93" />
                    <SPLIT distance="1150" swimtime="00:16:42.82" />
                    <SPLIT distance="1200" swimtime="00:17:27.72" />
                    <SPLIT distance="1250" swimtime="00:18:12.56" />
                    <SPLIT distance="1300" swimtime="00:18:57.33" />
                    <SPLIT distance="1350" swimtime="00:19:42.88" />
                    <SPLIT distance="1400" swimtime="00:20:27.42" />
                    <SPLIT distance="1450" swimtime="00:21:11.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="601" reactiontime="+89" swimtime="00:01:06.16" resultid="4941" heatid="7988" lane="4" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="530" reactiontime="+90" swimtime="00:02:54.92" resultid="4942" heatid="8025" lane="8" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.53" />
                    <SPLIT distance="100" swimtime="00:01:24.81" />
                    <SPLIT distance="150" swimtime="00:02:11.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="633" reactiontime="+90" swimtime="00:00:29.29" resultid="4943" heatid="8058" lane="7" entrytime="00:00:29.50" />
                <RESULT eventid="1432" points="499" reactiontime="+97" swimtime="00:05:22.86" resultid="4944" heatid="8153" lane="7" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                    <SPLIT distance="100" swimtime="00:01:19.24" />
                    <SPLIT distance="150" swimtime="00:02:00.73" />
                    <SPLIT distance="200" swimtime="00:02:42.73" />
                    <SPLIT distance="250" swimtime="00:03:22.57" />
                    <SPLIT distance="300" swimtime="00:04:03.31" />
                    <SPLIT distance="350" swimtime="00:04:43.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="495" reactiontime="+90" swimtime="00:02:30.81" resultid="4945" heatid="8099" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                    <SPLIT distance="100" swimtime="00:01:12.65" />
                    <SPLIT distance="150" swimtime="00:01:52.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="512" reactiontime="+91" swimtime="00:00:36.55" resultid="4946" heatid="8113" lane="4" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-03-01" firstname="Jan" gender="M" lastname="Wilczek" nation="POL" athleteid="4962">
              <RESULTS>
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="4963" heatid="7968" lane="2" entrytime="00:00:31.50" />
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="4964" heatid="7986" lane="3" entrytime="00:01:08.00" />
                <RESULT eventid="1372" status="DNS" swimtime="00:00:00.00" resultid="4965" heatid="8058" lane="3" entrytime="00:00:29.40" />
                <RESULT eventid="1462" status="DNS" swimtime="00:00:00.00" resultid="4966" heatid="8084" lane="3" entrytime="00:01:16.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-28" firstname="Jerzy" gender="M" lastname="Mroziński" nation="POL" athleteid="4947">
              <RESULTS>
                <RESULT eventid="1105" points="626" reactiontime="+84" swimtime="00:00:33.35" resultid="4948" heatid="7965" lane="4" entrytime="00:00:35.00" />
                <RESULT eventid="1228" points="651" swimtime="00:00:35.81" resultid="4949" heatid="8007" lane="2" entrytime="00:00:36.00" />
                <RESULT eventid="1402" points="740" reactiontime="+87" swimtime="00:03:03.07" resultid="4950" heatid="8075" lane="9" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.68" />
                    <SPLIT distance="100" swimtime="00:01:27.08" />
                    <SPLIT distance="150" swimtime="00:02:15.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="537" reactiontime="+86" swimtime="00:02:47.46" resultid="4951" heatid="8098" lane="0" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.33" />
                    <SPLIT distance="100" swimtime="00:01:18.25" />
                    <SPLIT distance="150" swimtime="00:02:02.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="710" reactiontime="+84" swimtime="00:01:21.64" resultid="4952" heatid="8129" lane="4" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="MAL" clubid="4983" name="Unia Oświęcim Masters">
          <CONTACT name="Szpara" />
          <ATHLETES>
            <ATHLETE birthdate="1969-02-05" firstname="Krzysztof" gender="M" lastname="Szpara" nation="POL" athleteid="4984">
              <RESULTS>
                <RESULT eventid="1198" points="730" reactiontime="+74" swimtime="00:01:02.00" resultid="4985" heatid="7990" lane="3" entrytime="00:01:01.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="667" reactiontime="+74" swimtime="00:02:42.08" resultid="4986" heatid="8027" lane="0" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.36" />
                    <SPLIT distance="100" swimtime="00:01:16.46" />
                    <SPLIT distance="150" swimtime="00:01:59.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="681" reactiontime="+71" swimtime="00:01:12.62" resultid="4987" heatid="8042" lane="2" entrytime="00:01:09.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="741" reactiontime="+78" swimtime="00:00:27.80" resultid="4988" heatid="8059" lane="6" entrytime="00:00:28.98" />
                <RESULT eventid="1539" points="644" reactiontime="+72" status="EXH" swimtime="00:00:33.85" resultid="8274" heatid="8108" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="031" nation="POL" region="LOD" clubid="4989" name="UTW &quot;Masters&quot; Zgierz">
          <CONTACT city="ZGIERZ" email="roman.wiczel@gmail.com" name="WICZEL" phone="691-928-922" state="ŁÓDZK" street="ŁĘCZYCKA 24" zip="95-100" />
          <ATHLETES>
            <ATHLETE birthdate="1957-01-09" firstname="Włodzimierz" gender="M" lastname="Przytulski" nation="POL" license="503105700027" athleteid="5054">
              <RESULTS>
                <RESULT eventid="1075" points="698" reactiontime="+91" swimtime="00:02:54.72" resultid="5055" heatid="7950" lane="2" entrytime="00:02:55.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.76" />
                    <SPLIT distance="100" swimtime="00:01:21.80" />
                    <SPLIT distance="150" swimtime="00:02:15.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="674" reactiontime="+89" swimtime="00:00:32.53" resultid="5056" heatid="7967" lane="3" entrytime="00:00:32.50" entrycourse="LCM" />
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="5057" heatid="7987" lane="0" entrytime="00:01:07.50" entrycourse="LCM" />
                <RESULT eventid="1258" points="541" reactiontime="+97" swimtime="00:03:10.39" resultid="5058" heatid="8016" lane="7" entrytime="00:03:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.95" />
                    <SPLIT distance="100" swimtime="00:01:29.62" />
                    <SPLIT distance="150" swimtime="00:02:19.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" status="DNS" swimtime="00:00:00.00" resultid="5059" heatid="8040" lane="0" entrytime="00:01:20.00" entrycourse="LCM" />
                <RESULT eventid="1462" points="526" reactiontime="+88" swimtime="00:01:20.02" resultid="5060" heatid="8084" lane="7" entrytime="00:01:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="713" reactiontime="+85" swimtime="00:02:32.33" resultid="5061" heatid="8099" lane="8" entrytime="00:02:32.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                    <SPLIT distance="100" swimtime="00:01:11.13" />
                    <SPLIT distance="150" swimtime="00:01:51.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" status="DNS" swimtime="00:00:00.00" resultid="5062" heatid="8113" lane="0" entrytime="00:00:36.20" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-03-03" firstname="Urszula" gender="F" lastname="Mróz" nation="POL" license="503105600030" athleteid="5006">
              <RESULTS>
                <RESULT eventid="1058" points="603" reactiontime="+96" swimtime="00:03:12.03" resultid="5007" heatid="7942" lane="5" entrytime="00:03:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.99" />
                    <SPLIT distance="100" swimtime="00:01:27.47" />
                    <SPLIT distance="150" swimtime="00:02:26.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="609" reactiontime="+88" swimtime="00:00:35.66" resultid="5008" heatid="7958" lane="9" entrytime="00:00:37.30" entrycourse="LCM" />
                <RESULT eventid="1181" points="589" reactiontime="+92" swimtime="00:01:16.60" resultid="5009" heatid="7976" lane="1" entrytime="00:01:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="626" reactiontime="+85" swimtime="00:03:15.10" resultid="5010" heatid="8019" lane="3" entrytime="00:03:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.91" />
                    <SPLIT distance="100" swimtime="00:01:34.29" />
                    <SPLIT distance="150" swimtime="00:02:25.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="623" reactiontime="+74" swimtime="00:01:28.27" resultid="5011" heatid="8033" lane="4" entrytime="00:01:31.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="550" reactiontime="+91" swimtime="00:01:27.19" resultid="5012" heatid="8079" lane="6" entrytime="00:01:27.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="636" reactiontime="+82" swimtime="00:00:39.94" resultid="5013" heatid="8106" lane="0" entrytime="00:00:39.30" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1922-01-04" firstname="Kazimierz" gender="M" lastname="Mrówczyński" nation="POL" license="503105700021" athleteid="5075">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1198" points="537" reactiontime="+107" swimtime="00:02:22.78" resultid="5076" heatid="7981" lane="0" entrytime="00:02:53.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.31" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1228" points="505" reactiontime="+118" swimtime="00:01:16.54" resultid="5077" heatid="8000" lane="1" entrytime="00:01:18.00" entrycourse="LCM" />
                <RESULT comment="Rekord Polski Masters" eventid="1372" points="471" reactiontime="+99" swimtime="00:00:59.76" resultid="5078" heatid="8052" lane="1" entrytime="00:01:00.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-05-12" firstname="Tadeusz" gender="M" lastname="Obiedziński" nation="POL" license="503105700038" athleteid="5030">
              <RESULTS>
                <RESULT eventid="1075" points="362" reactiontime="+110" swimtime="00:03:37.48" resultid="5031" heatid="7948" lane="9" entrytime="00:03:27.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.41" />
                    <SPLIT distance="100" swimtime="00:01:48.34" />
                    <SPLIT distance="150" swimtime="00:02:45.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="456" reactiontime="+88" swimtime="00:00:40.33" resultid="5032" heatid="8004" lane="2" entrytime="00:00:40.88" entrycourse="LCM" />
                <RESULT eventid="1402" points="402" reactiontime="+97" swimtime="00:03:44.21" resultid="5033" heatid="8072" lane="5" entrytime="00:03:43.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.31" />
                    <SPLIT distance="100" swimtime="00:01:44.90" />
                    <SPLIT distance="150" swimtime="00:02:45.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="397" reactiontime="+88" swimtime="00:01:39.07" resultid="5034" heatid="8127" lane="3" entrytime="00:01:34.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-03-18" firstname="Daria" gender="F" lastname="Fajkowska" nation="POL" license="503105600018" athleteid="4999">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1058" points="863" reactiontime="+95" swimtime="00:02:39.04" resultid="5000" heatid="7944" lane="5" entrytime="00:02:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.66" />
                    <SPLIT distance="100" swimtime="00:01:11.93" />
                    <SPLIT distance="150" swimtime="00:01:58.63" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1273" points="854" reactiontime="+78" swimtime="00:02:42.29" resultid="5001" heatid="8021" lane="6" entrytime="00:02:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                    <SPLIT distance="100" swimtime="00:01:16.89" />
                    <SPLIT distance="150" swimtime="00:01:59.79" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1326" points="894" reactiontime="+76" swimtime="00:01:12.74" resultid="5002" heatid="8035" lane="5" entrytime="00:01:14.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="771" reactiontime="+91" swimtime="00:00:30.04" resultid="5003" heatid="8050" lane="9" entrytime="00:00:29.40" entrycourse="LCM" />
                <RESULT comment="Rekord Polski Masters" eventid="1524" points="904" reactiontime="+64" swimtime="00:00:33.79" resultid="5004" heatid="8107" lane="6" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT comment="Rekord Polski Masters" eventid="1584" points="783" reactiontime="+97" swimtime="00:05:51.92" resultid="5005" heatid="8159" lane="4" entrytime="00:05:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                    <SPLIT distance="100" swimtime="00:01:16.55" />
                    <SPLIT distance="150" swimtime="00:02:02.10" />
                    <SPLIT distance="200" swimtime="00:02:46.61" />
                    <SPLIT distance="250" swimtime="00:03:36.60" />
                    <SPLIT distance="300" swimtime="00:04:27.06" />
                    <SPLIT distance="350" swimtime="00:05:10.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-02-07" firstname="Krzysztof" gender="M" lastname="Wojciechowski" nation="POL" license="503105700024" athleteid="5021">
              <RESULTS>
                <RESULT eventid="1075" points="474" reactiontime="+110" swimtime="00:03:32.33" resultid="5022" heatid="7947" lane="4" entrytime="00:03:29.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.94" />
                    <SPLIT distance="100" swimtime="00:01:48.35" />
                    <SPLIT distance="150" swimtime="00:02:45.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="716" reactiontime="+104" swimtime="00:00:40.52" resultid="5023" heatid="8005" lane="0" entrytime="00:00:39.90" entrycourse="LCM" />
                <RESULT eventid="1402" points="635" reactiontime="+104" swimtime="00:03:40.42" resultid="5024" heatid="8073" lane="5" entrytime="00:03:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.25" />
                    <SPLIT distance="100" swimtime="00:01:44.53" />
                    <SPLIT distance="150" swimtime="00:02:43.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="654" reactiontime="+104" swimtime="00:01:34.87" resultid="5025" heatid="8128" lane="8" entrytime="00:01:32.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-09-12" firstname="Małgorzata" gender="F" lastname="Ścibiorek" nation="POL" license="503105600028" athleteid="4994">
              <RESULTS>
                <RESULT eventid="1090" points="797" reactiontime="+94" swimtime="00:00:32.13" resultid="4995" heatid="7960" lane="7" entrytime="00:00:32.30" entrycourse="LCM" />
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1243" points="728" reactiontime="+88" swimtime="00:02:49.96" resultid="4996" heatid="8012" lane="4" entrytime="00:02:46.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.37" />
                    <SPLIT distance="100" swimtime="00:01:16.81" />
                    <SPLIT distance="150" swimtime="00:02:01.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="804" reactiontime="+88" swimtime="00:01:11.90" resultid="4997" heatid="8080" lane="3" entrytime="00:01:11.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="674" reactiontime="+89" swimtime="00:01:27.57" resultid="4998" heatid="8123" lane="3" entrytime="00:01:24.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-22" firstname="Roman" gender="M" lastname="Wiczel" nation="POL" license="503105700034" athleteid="4990">
              <RESULTS>
                <RESULT eventid="1228" points="738" reactiontime="+75" swimtime="00:00:40.11" resultid="4991" heatid="8005" lane="8" entrytime="00:00:39.50" entrycourse="LCM" />
                <RESULT eventid="1402" points="774" reactiontime="+77" swimtime="00:03:26.37" resultid="4992" heatid="8074" lane="8" entrytime="00:03:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.00" />
                    <SPLIT distance="100" swimtime="00:01:39.55" />
                    <SPLIT distance="150" swimtime="00:02:33.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="749" reactiontime="+86" swimtime="00:01:30.68" resultid="4993" heatid="8128" lane="2" entrytime="00:01:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-04-07" firstname="Ewa" gender="F" lastname="Stępień" nation="POL" license="503105600029" athleteid="5063">
              <RESULTS>
                <RESULT eventid="1090" points="648" reactiontime="+69" swimtime="00:00:34.93" resultid="5064" heatid="7957" lane="4" entrytime="00:00:37.31" entrycourse="LCM" />
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1181" points="677" reactiontime="+70" swimtime="00:01:13.10" resultid="5065" heatid="7977" lane="2" entrytime="00:01:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="839" reactiontime="+71" swimtime="00:00:40.01" resultid="5066" heatid="7999" lane="0" entrytime="00:00:40.00" entrycourse="LCM" />
                <RESULT comment="Rekord Polski Masters" eventid="1357" points="710" reactiontime="+71" swimtime="00:00:31.84" resultid="5067" heatid="8048" lane="6" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="1387" status="DNS" swimtime="00:00:00.00" resultid="5068" heatid="8069" lane="5" entrytime="00:03:20.00" entrycourse="LCM" />
                <RESULT eventid="1554" points="789" reactiontime="+67" swimtime="00:01:30.32" resultid="5069" heatid="8122" lane="6" entrytime="00:01:30.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-06-10" firstname="Sonia" gender="F" lastname="Bochyńska" nation="POL" license="503105600046" athleteid="5035">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1090" points="813" reactiontime="+76" swimtime="00:00:30.32" resultid="5036" heatid="7960" lane="4" entrytime="00:00:29.70" entrycourse="LCM" />
                <RESULT eventid="1181" points="799" reactiontime="+76" swimtime="00:01:03.31" resultid="5037" heatid="7979" lane="5" entrytime="00:01:00.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="836" reactiontime="+75" swimtime="00:00:28.71" resultid="5038" heatid="8050" lane="5" entrytime="00:00:28.00" entrycourse="LCM" />
                <RESULT eventid="1493" status="DNS" swimtime="00:00:00.00" resultid="5039" heatid="8092" lane="4" entrytime="00:02:10.00" entrycourse="LCM" />
                <RESULT comment="Rekord Polski Masters" eventid="1524" points="901" reactiontime="+66" swimtime="00:00:32.19" resultid="5040" heatid="8107" lane="4" entrytime="00:00:30.30" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-03-11" firstname="Adrian" gender="M" lastname="Pawlak" nation="POL" license="503105700045" athleteid="5026">
              <RESULTS>
                <RESULT eventid="1075" points="455" reactiontime="+66" swimtime="00:02:43.68" resultid="5027" heatid="7952" lane="3" entrytime="00:02:35.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.92" />
                    <SPLIT distance="100" swimtime="00:01:13.92" />
                    <SPLIT distance="150" swimtime="00:02:03.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="529" reactiontime="+62" swimtime="00:00:36.22" resultid="5028" heatid="8009" lane="2" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT eventid="1372" points="696" reactiontime="+63" swimtime="00:00:26.12" resultid="5029" heatid="8065" lane="8" entrytime="00:00:26.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-03-01" firstname="Waldemar" gender="M" lastname="Jagiełło" nation="POL" license="503105700036" athleteid="5046">
              <RESULTS>
                <RESULT eventid="1075" points="723" reactiontime="+85" swimtime="00:02:30.54" resultid="5047" heatid="7953" lane="9" entrytime="00:02:27.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.57" />
                    <SPLIT distance="100" swimtime="00:01:09.70" />
                    <SPLIT distance="150" swimtime="00:01:53.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="703" reactiontime="+85" swimtime="00:00:28.69" resultid="5048" heatid="7972" lane="7" entrytime="00:00:27.30" entrycourse="LCM" />
                <RESULT eventid="1198" points="645" reactiontime="+88" swimtime="00:01:00.15" resultid="5049" heatid="7991" lane="2" entrytime="00:01:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="635" reactiontime="+94" swimtime="00:00:33.97" resultid="5050" heatid="8009" lane="6" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT comment="Rekord Polski Masters" eventid="1372" points="728" reactiontime="+80" swimtime="00:00:26.15" resultid="5051" heatid="8063" lane="2" entrytime="00:00:26.50" entrycourse="LCM" />
                <RESULT eventid="1462" points="645" reactiontime="+91" swimtime="00:01:07.38" resultid="5052" heatid="8085" lane="3" entrytime="00:01:06.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="740" reactiontime="+79" swimtime="00:00:31.17" resultid="5053" heatid="8116" lane="6" entrytime="00:00:30.70" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-12-03" firstname="Zbigniew" gender="M" lastname="Maciejczyk" nation="POL" license="503105700026" athleteid="5014">
              <RESULTS>
                <RESULT eventid="1105" points="545" reactiontime="+96" swimtime="00:00:37.36" resultid="5015" heatid="7964" lane="7" entrytime="00:00:38.00" entrycourse="LCM" />
                <RESULT eventid="1198" points="544" reactiontime="+106" swimtime="00:01:20.83" resultid="5016" heatid="7984" lane="0" entrytime="00:01:19.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="226" reactiontime="+112" swimtime="00:04:48.91" resultid="5017" heatid="8015" lane="9" entrytime="00:04:10.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.58" />
                    <SPLIT distance="100" swimtime="00:02:26.81" />
                    <SPLIT distance="150" swimtime="00:03:44.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="618" reactiontime="+95" swimtime="00:00:33.80" resultid="5018" heatid="8055" lane="9" entrytime="00:00:34.00" entrycourse="LCM" />
                <RESULT eventid="1462" points="278" reactiontime="+105" swimtime="00:01:51.94" resultid="5019" heatid="8082" lane="5" entrytime="00:01:37.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="380" reactiontime="+75" swimtime="00:00:46.25" resultid="5020" heatid="8110" lane="4" entrytime="00:00:45.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-02-16" firstname="Adrian" gender="M" lastname="Styrzyński" nation="POL" license="503105700033" athleteid="5041">
              <RESULTS>
                <RESULT eventid="1075" points="683" reactiontime="+77" swimtime="00:02:23.03" resultid="5042" heatid="7953" lane="6" entrytime="00:02:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.76" />
                    <SPLIT distance="100" swimtime="00:01:05.65" />
                    <SPLIT distance="150" swimtime="00:01:48.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="722" reactiontime="+71" swimtime="00:00:32.65" resultid="5043" heatid="8010" lane="8" entrytime="00:00:32.00" entrycourse="LCM" />
                <RESULT eventid="1462" points="787" reactiontime="+75" swimtime="00:01:01.57" resultid="5044" heatid="8086" lane="3" entrytime="00:01:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="633" reactiontime="+69" swimtime="00:01:15.28" resultid="5045" heatid="8132" lane="6" entrytime="00:01:09.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1318" reactiontime="+74" swimtime="00:04:20.37" resultid="5070" heatid="8030" lane="5" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.43" />
                    <SPLIT distance="100" swimtime="00:00:57.45" />
                    <SPLIT distance="150" swimtime="00:01:35.14" />
                    <SPLIT distance="200" swimtime="00:02:20.56" />
                    <SPLIT distance="250" swimtime="00:02:48.82" />
                    <SPLIT distance="300" swimtime="00:03:20.56" />
                    <SPLIT distance="350" swimtime="00:03:49.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5046" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="5014" number="2" reactiontime="+88" />
                    <RELAYPOSITION athleteid="5026" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="5041" number="4" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1614" swimtime="00:02:02.77" resultid="5071" heatid="8135" lane="5" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                    <SPLIT distance="100" swimtime="00:01:04.97" />
                    <SPLIT distance="150" swimtime="00:01:37.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5035" number="1" />
                    <RELAYPOSITION athleteid="5041" number="2" />
                    <RELAYPOSITION athleteid="4994" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="5026" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1614" reactiontime="+77" swimtime="00:02:26.34" resultid="5072" heatid="8134" lane="8" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.87" />
                    <SPLIT distance="100" swimtime="00:01:18.60" />
                    <SPLIT distance="150" swimtime="00:01:53.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5006" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="4990" number="2" />
                    <RELAYPOSITION athleteid="5063" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="5014" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" region="WAR" clubid="5079" name="Victory Masters Elbląg">
          <CONTACT city="Elbląg" name="Latecki Grzegorz" street="Łokietka 45" zip="82-300" />
          <ATHLETES>
            <ATHLETE birthdate="1954-02-04" firstname="Ewa" gender="F" lastname="Kerner-Mateusiak" nation="POL" athleteid="5100">
              <RESULTS>
                <RESULT eventid="1120" points="252" swimtime="00:18:38.44" resultid="5101" heatid="8138" lane="5" entrytime="00:20:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.36" />
                    <SPLIT distance="100" swimtime="00:02:07.72" />
                    <SPLIT distance="150" swimtime="00:03:19.72" />
                    <SPLIT distance="200" swimtime="00:04:31.60" />
                    <SPLIT distance="250" swimtime="00:05:42.96" />
                    <SPLIT distance="300" swimtime="00:06:53.58" />
                    <SPLIT distance="350" swimtime="00:08:04.24" />
                    <SPLIT distance="400" swimtime="00:09:15.62" />
                    <SPLIT distance="450" swimtime="00:10:26.90" />
                    <SPLIT distance="500" swimtime="00:11:38.22" />
                    <SPLIT distance="550" swimtime="00:12:49.65" />
                    <SPLIT distance="600" swimtime="00:14:00.92" />
                    <SPLIT distance="650" swimtime="00:15:11.40" />
                    <SPLIT distance="700" swimtime="00:16:22.72" />
                    <SPLIT distance="750" swimtime="00:17:32.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="184" reactiontime="+116" swimtime="00:02:03.43" resultid="5102" heatid="7973" lane="6" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="164" reactiontime="+122" swimtime="00:01:10.28" resultid="5103" heatid="7994" lane="5" entrytime="00:01:10.00" />
                <RESULT eventid="1326" points="180" reactiontime="+98" swimtime="00:02:26.44" resultid="5104" heatid="8032" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="267" reactiontime="+114" swimtime="00:09:01.55" resultid="5105" heatid="8150" lane="4" entrytime="00:09:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.73" />
                    <SPLIT distance="100" swimtime="00:02:04.68" />
                    <SPLIT distance="150" swimtime="00:03:15.52" />
                    <SPLIT distance="200" swimtime="00:04:25.83" />
                    <SPLIT distance="250" swimtime="00:05:35.87" />
                    <SPLIT distance="300" swimtime="00:06:45.79" />
                    <SPLIT distance="350" swimtime="00:07:54.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="237" reactiontime="+82" swimtime="00:01:04.85" resultid="5106" heatid="8103" lane="4" entrytime="00:01:10.00" />
                <RESULT eventid="1554" points="188" reactiontime="+126" swimtime="00:02:36.86" resultid="5107" heatid="8119" lane="0" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-03-12" firstname="Grzegorz" gender="M" lastname="Latecki" nation="POL" athleteid="5080">
              <RESULTS>
                <RESULT eventid="1105" points="769" reactiontime="+83" swimtime="00:00:30.33" resultid="5081" heatid="7969" lane="0" entrytime="00:00:31.00" />
                <RESULT eventid="1228" points="573" reactiontime="+77" swimtime="00:00:38.74" resultid="5082" heatid="8004" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1372" points="651" reactiontime="+80" swimtime="00:00:29.30" resultid="5083" heatid="8060" lane="8" entrytime="00:00:28.50" />
                <RESULT eventid="1539" points="702" reactiontime="+75" swimtime="00:00:34.34" resultid="5084" heatid="8114" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="1599" points="635" reactiontime="+83" swimtime="00:06:10.68" resultid="5085" heatid="8164" lane="4" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.41" />
                    <SPLIT distance="100" swimtime="00:01:31.74" />
                    <SPLIT distance="150" swimtime="00:02:19.56" />
                    <SPLIT distance="200" swimtime="00:03:06.62" />
                    <SPLIT distance="250" swimtime="00:03:57.49" />
                    <SPLIT distance="300" swimtime="00:04:48.65" />
                    <SPLIT distance="350" swimtime="00:05:30.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-05-05" firstname="Beata" gender="F" lastname="Karaś" nation="POL" athleteid="5092">
              <RESULTS>
                <RESULT eventid="1150" points="484" reactiontime="+107" swimtime="00:28:00.40" resultid="5093" heatid="8142" lane="7" entrytime="00:30:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.77" />
                    <SPLIT distance="100" swimtime="00:01:46.78" />
                    <SPLIT distance="150" swimtime="00:02:42.06" />
                    <SPLIT distance="200" swimtime="00:03:37.95" />
                    <SPLIT distance="250" swimtime="00:04:34.51" />
                    <SPLIT distance="300" swimtime="00:05:31.43" />
                    <SPLIT distance="350" swimtime="00:06:27.67" />
                    <SPLIT distance="400" swimtime="00:07:25.67" />
                    <SPLIT distance="450" swimtime="00:08:22.74" />
                    <SPLIT distance="500" swimtime="00:09:19.37" />
                    <SPLIT distance="550" swimtime="00:10:16.02" />
                    <SPLIT distance="600" swimtime="00:11:13.22" />
                    <SPLIT distance="650" swimtime="00:12:10.62" />
                    <SPLIT distance="700" swimtime="00:13:08.26" />
                    <SPLIT distance="750" swimtime="00:14:04.38" />
                    <SPLIT distance="800" swimtime="00:15:00.54" />
                    <SPLIT distance="850" swimtime="00:15:56.66" />
                    <SPLIT distance="900" swimtime="00:16:51.51" />
                    <SPLIT distance="950" swimtime="00:17:48.38" />
                    <SPLIT distance="1000" swimtime="00:18:45.19" />
                    <SPLIT distance="1050" swimtime="00:19:41.01" />
                    <SPLIT distance="1100" swimtime="00:20:37.28" />
                    <SPLIT distance="1150" swimtime="00:21:33.36" />
                    <SPLIT distance="1200" swimtime="00:22:30.28" />
                    <SPLIT distance="1250" swimtime="00:23:26.52" />
                    <SPLIT distance="1300" swimtime="00:24:22.87" />
                    <SPLIT distance="1350" swimtime="00:25:18.49" />
                    <SPLIT distance="1400" swimtime="00:26:13.63" />
                    <SPLIT distance="1450" swimtime="00:27:07.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="272" reactiontime="+97" swimtime="00:01:39.10" resultid="5094" heatid="7974" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1243" points="323" reactiontime="+106" swimtime="00:04:18.38" resultid="5095" heatid="8011" lane="4" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.80" />
                    <SPLIT distance="100" swimtime="00:02:01.17" />
                    <SPLIT distance="150" swimtime="00:03:08.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="289" reactiontime="+98" swimtime="00:07:19.98" resultid="5096" heatid="8149" lane="8" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.52" />
                    <SPLIT distance="100" swimtime="00:01:47.07" />
                    <SPLIT distance="150" swimtime="00:02:43.51" />
                    <SPLIT distance="200" swimtime="00:03:40.95" />
                    <SPLIT distance="250" swimtime="00:04:36.49" />
                    <SPLIT distance="300" swimtime="00:05:32.97" />
                    <SPLIT distance="350" swimtime="00:06:27.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="217" reactiontime="+109" swimtime="00:01:58.88" resultid="5097" heatid="8078" lane="7" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="279" reactiontime="+102" swimtime="00:03:31.17" resultid="5098" heatid="8089" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.88" />
                    <SPLIT distance="100" swimtime="00:01:42.90" />
                    <SPLIT distance="150" swimtime="00:02:37.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1584" points="307" reactiontime="+109" swimtime="00:08:44.38" resultid="5099" heatid="8161" lane="5" entrytime="00:08:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.03" />
                    <SPLIT distance="100" swimtime="00:01:57.49" />
                    <SPLIT distance="150" swimtime="00:03:13.79" />
                    <SPLIT distance="200" swimtime="00:04:25.24" />
                    <SPLIT distance="250" swimtime="00:05:41.33" />
                    <SPLIT distance="300" swimtime="00:06:58.62" />
                    <SPLIT distance="350" swimtime="00:07:52.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-08-31" firstname="Karolina" gender="F" lastname="Karaś" nation="POL" athleteid="5086">
              <RESULTS>
                <RESULT eventid="1120" points="247" reactiontime="+100" swimtime="00:14:47.55" resultid="5087" heatid="8137" lane="5" entrytime="00:13:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.27" />
                    <SPLIT distance="100" swimtime="00:01:48.08" />
                    <SPLIT distance="150" swimtime="00:02:45.55" />
                    <SPLIT distance="200" swimtime="00:03:43.26" />
                    <SPLIT distance="250" swimtime="00:04:40.81" />
                    <SPLIT distance="300" swimtime="00:05:38.46" />
                    <SPLIT distance="350" swimtime="00:06:35.86" />
                    <SPLIT distance="400" swimtime="00:07:32.84" />
                    <SPLIT distance="450" swimtime="00:08:27.65" />
                    <SPLIT distance="500" swimtime="00:09:22.54" />
                    <SPLIT distance="550" swimtime="00:10:16.80" />
                    <SPLIT distance="600" swimtime="00:11:12.44" />
                    <SPLIT distance="650" swimtime="00:12:07.47" />
                    <SPLIT distance="700" swimtime="00:13:02.18" />
                    <SPLIT distance="750" swimtime="00:13:56.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="230" reactiontime="+98" swimtime="00:01:35.79" resultid="5088" heatid="7974" lane="7" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="238" reactiontime="+91" swimtime="00:00:43.63" resultid="5089" heatid="8045" lane="1" entrytime="00:00:45.00" />
                <RESULT eventid="1417" points="258" reactiontime="+99" swimtime="00:07:08.66" resultid="5090" heatid="8148" lane="0" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.93" />
                    <SPLIT distance="100" swimtime="00:01:39.02" />
                    <SPLIT distance="150" swimtime="00:02:32.69" />
                    <SPLIT distance="200" swimtime="00:03:28.26" />
                    <SPLIT distance="250" swimtime="00:04:25.05" />
                    <SPLIT distance="300" swimtime="00:05:20.81" />
                    <SPLIT distance="350" swimtime="00:06:15.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="270" reactiontime="+88" swimtime="00:03:19.36" resultid="5091" heatid="8088" lane="2" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.23" />
                    <SPLIT distance="100" swimtime="00:01:37.20" />
                    <SPLIT distance="150" swimtime="00:02:28.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WMT" nation="POL" region="MAZ" clubid="2762" name="Warsaw Masters Team">
          <CONTACT city="Warszawa" email="wojciech.kaluzynski@gmail.com" name="Kałużyński Wojciech" phone="607 45 4444" />
          <ATHLETES>
            <ATHLETE birthdate="1989-07-10" firstname="Sandra" gender="F" lastname="Pietrzak" nation="POL" athleteid="2956">
              <RESULTS>
                <RESULT eventid="1120" points="738" reactiontime="+77" swimtime="00:10:16.32" resultid="2957" heatid="8136" lane="5" entrytime="00:10:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                    <SPLIT distance="100" swimtime="00:01:09.22" />
                    <SPLIT distance="150" swimtime="00:01:46.67" />
                    <SPLIT distance="200" swimtime="00:02:25.06" />
                    <SPLIT distance="250" swimtime="00:03:03.43" />
                    <SPLIT distance="300" swimtime="00:03:42.25" />
                    <SPLIT distance="350" swimtime="00:04:21.21" />
                    <SPLIT distance="400" swimtime="00:05:00.48" />
                    <SPLIT distance="450" swimtime="00:05:40.00" />
                    <SPLIT distance="500" swimtime="00:06:19.39" />
                    <SPLIT distance="550" swimtime="00:06:59.06" />
                    <SPLIT distance="600" swimtime="00:07:38.89" />
                    <SPLIT distance="650" swimtime="00:08:18.70" />
                    <SPLIT distance="700" swimtime="00:08:58.09" />
                    <SPLIT distance="750" swimtime="00:09:37.54" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1273" points="796" reactiontime="+70" swimtime="00:02:38.44" resultid="2958" heatid="8021" lane="7" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                    <SPLIT distance="100" swimtime="00:01:15.87" />
                    <SPLIT distance="150" swimtime="00:01:56.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="768" reactiontime="+73" swimtime="00:01:14.02" resultid="2959" heatid="8035" lane="7" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="740" reactiontime="+80" swimtime="00:05:01.75" resultid="2960" heatid="8147" lane="4" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.50" />
                    <SPLIT distance="100" swimtime="00:01:10.20" />
                    <SPLIT distance="150" swimtime="00:01:48.19" />
                    <SPLIT distance="200" swimtime="00:02:26.10" />
                    <SPLIT distance="250" swimtime="00:03:04.43" />
                    <SPLIT distance="300" swimtime="00:03:43.45" />
                    <SPLIT distance="350" swimtime="00:04:23.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="781" reactiontime="+77" swimtime="00:02:19.98" resultid="2961" heatid="8092" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                    <SPLIT distance="100" swimtime="00:01:06.61" />
                    <SPLIT distance="150" swimtime="00:01:42.81" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1584" points="787" reactiontime="+80" swimtime="00:05:37.73" resultid="2962" heatid="8159" lane="5" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.00" />
                    <SPLIT distance="100" swimtime="00:01:14.81" />
                    <SPLIT distance="150" swimtime="00:01:57.75" />
                    <SPLIT distance="200" swimtime="00:02:41.13" />
                    <SPLIT distance="250" swimtime="00:03:29.63" />
                    <SPLIT distance="300" swimtime="00:04:19.00" />
                    <SPLIT distance="350" swimtime="00:05:00.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-10" firstname="Michał" gender="M" lastname="Rudziński" nation="POL" athleteid="2853">
              <RESULTS>
                <RESULT eventid="1105" points="303" reactiontime="+101" swimtime="00:00:40.52" resultid="2854" heatid="7963" lane="2" entrytime="00:00:43.79" />
                <RESULT eventid="1258" points="162" reactiontime="+115" swimtime="00:04:15.31" resultid="2855" heatid="8014" lane="1" entrytime="00:04:43.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.69" />
                    <SPLIT distance="100" swimtime="00:01:58.37" />
                    <SPLIT distance="150" swimtime="00:03:06.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="397" reactiontime="+106" swimtime="00:03:29.11" resultid="2856" heatid="8073" lane="3" entrytime="00:03:30.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.22" />
                    <SPLIT distance="100" swimtime="00:01:38.76" />
                    <SPLIT distance="150" swimtime="00:02:34.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="357" reactiontime="+116" swimtime="00:01:37.08" resultid="2857" heatid="8124" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="299" reactiontime="+102" swimtime="00:07:46.98" resultid="2858" heatid="8166" lane="2" entrytime="00:07:44.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.65" />
                    <SPLIT distance="100" swimtime="00:01:50.01" />
                    <SPLIT distance="150" swimtime="00:02:59.85" />
                    <SPLIT distance="200" swimtime="00:04:08.30" />
                    <SPLIT distance="250" swimtime="00:05:02.78" />
                    <SPLIT distance="300" swimtime="00:05:59.78" />
                    <SPLIT distance="350" swimtime="00:06:55.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-05-14" firstname="Wojciech" gender="M" lastname="Kałużyński" nation="POL" athleteid="2969">
              <RESULTS>
                <RESULT eventid="1105" points="369" reactiontime="+74" swimtime="00:00:35.57" resultid="2970" heatid="7965" lane="9" entrytime="00:00:35.77" />
                <RESULT eventid="1198" points="419" reactiontime="+75" swimtime="00:01:09.43" resultid="2971" heatid="7986" lane="4" entrytime="00:01:07.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="414" reactiontime="+80" swimtime="00:00:31.55" resultid="2972" heatid="8057" lane="9" entrytime="00:00:30.53" />
                <RESULT eventid="1432" points="364" reactiontime="+84" swimtime="00:05:59.06" resultid="2973" heatid="8153" lane="0" entrytime="00:05:37.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                    <SPLIT distance="100" swimtime="00:01:20.22" />
                    <SPLIT distance="150" swimtime="00:02:04.48" />
                    <SPLIT distance="200" swimtime="00:02:50.57" />
                    <SPLIT distance="250" swimtime="00:03:37.16" />
                    <SPLIT distance="300" swimtime="00:04:24.54" />
                    <SPLIT distance="350" swimtime="00:05:12.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="349" reactiontime="+85" swimtime="00:02:44.16" resultid="2974" heatid="8099" lane="9" entrytime="00:02:33.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                    <SPLIT distance="100" swimtime="00:01:17.93" />
                    <SPLIT distance="150" swimtime="00:02:00.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="333" reactiontime="+96" swimtime="00:00:40.68" resultid="2975" heatid="8112" lane="1" entrytime="00:00:38.02" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-03" firstname="Robert" gender="M" lastname="Sutowski" nation="POL" athleteid="2910">
              <RESULTS>
                <RESULT eventid="1135" points="389" reactiontime="+106" swimtime="00:13:59.34" resultid="2912" heatid="8140" lane="0" entrytime="00:14:30.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.18" />
                    <SPLIT distance="100" swimtime="00:01:40.28" />
                    <SPLIT distance="150" swimtime="00:02:34.94" />
                    <SPLIT distance="200" swimtime="00:03:29.07" />
                    <SPLIT distance="250" swimtime="00:04:24.49" />
                    <SPLIT distance="300" swimtime="00:05:18.66" />
                    <SPLIT distance="350" swimtime="00:06:12.61" />
                    <SPLIT distance="400" swimtime="00:07:06.36" />
                    <SPLIT distance="450" swimtime="00:07:58.46" />
                    <SPLIT distance="500" swimtime="00:08:50.96" />
                    <SPLIT distance="550" swimtime="00:09:43.85" />
                    <SPLIT distance="600" swimtime="00:10:36.60" />
                    <SPLIT distance="650" swimtime="00:11:29.23" />
                    <SPLIT distance="700" swimtime="00:12:21.70" />
                    <SPLIT distance="750" swimtime="00:13:12.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="320" reactiontime="+109" swimtime="00:01:28.79" resultid="2913" heatid="7983" lane="9" entrytime="00:01:27.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="238" reactiontime="+85" swimtime="00:04:18.39" resultid="2914" heatid="8024" lane="0" entrytime="00:03:58.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.90" />
                    <SPLIT distance="100" swimtime="00:02:11.21" />
                    <SPLIT distance="150" swimtime="00:03:17.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="303" reactiontime="+115" swimtime="00:00:39.60" resultid="2915" heatid="8053" lane="9" entrytime="00:00:42.20" />
                <RESULT eventid="1432" points="377" reactiontime="+109" swimtime="00:06:48.35" resultid="2916" heatid="8155" lane="5" entrytime="00:06:39.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.95" />
                    <SPLIT distance="100" swimtime="00:01:39.02" />
                    <SPLIT distance="150" swimtime="00:02:32.71" />
                    <SPLIT distance="200" swimtime="00:03:25.63" />
                    <SPLIT distance="250" swimtime="00:04:18.51" />
                    <SPLIT distance="300" swimtime="00:05:10.59" />
                    <SPLIT distance="350" swimtime="00:06:01.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="349" reactiontime="+110" swimtime="00:03:13.33" resultid="2917" heatid="8095" lane="3" entrytime="00:03:13.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.61" />
                    <SPLIT distance="100" swimtime="00:01:35.67" />
                    <SPLIT distance="150" swimtime="00:02:26.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="193" reactiontime="+84" swimtime="00:00:56.21" resultid="2918" heatid="8110" lane="2" entrytime="00:00:47.20" />
                <RESULT eventid="1105" points="194" reactiontime="+109" swimtime="00:00:49.26" resultid="6025" heatid="7963" lane="8" entrytime="00:00:47.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-12-11" firstname="Igor" gender="M" lastname="Rębas" nation="POL" athleteid="2879">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="2880" heatid="7945" lane="1" />
                <RESULT eventid="1105" points="795" reactiontime="+71" swimtime="00:00:27.06" resultid="2881" heatid="7972" lane="2" entrytime="00:00:27.05" />
                <RESULT eventid="1198" points="685" reactiontime="+78" swimtime="00:00:58.66" resultid="2882" heatid="7993" lane="8" entrytime="00:00:57.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="715" reactiontime="+71" swimtime="00:00:25.88" resultid="2883" heatid="8064" lane="6" entrytime="00:00:26.04" />
                <RESULT eventid="1462" points="753" reactiontime="+72" swimtime="00:01:02.48" resultid="2884" heatid="8086" lane="2" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="521" reactiontime="+71" swimtime="00:00:33.27" resultid="2885" heatid="8114" lane="7" entrytime="00:00:34.00" />
                <RESULT eventid="1599" status="DNS" swimtime="00:00:00.00" resultid="2886" heatid="8162" lane="9" entrytime="00:05:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-11-11" firstname="Bolesław" gender="M" lastname="Szuter" nation="POL" athleteid="2777">
              <RESULTS>
                <RESULT eventid="1105" points="886" reactiontime="+79" swimtime="00:00:28.35" resultid="2778" heatid="7968" lane="7" entrytime="00:00:31.55" />
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1198" points="978" reactiontime="+75" swimtime="00:00:56.26" resultid="2779" heatid="7992" lane="5" entrytime="00:00:58.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.26" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1372" points="942" reactiontime="+81" swimtime="00:00:25.66" resultid="2780" heatid="8063" lane="5" entrytime="00:00:26.34" />
                <RESULT comment="Rekord Polski Masters" eventid="1509" points="849" reactiontime="+79" swimtime="00:02:06.06" resultid="2781" heatid="8102" lane="1" entrytime="00:02:10.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.68" />
                    <SPLIT distance="100" swimtime="00:01:02.11" />
                    <SPLIT distance="150" swimtime="00:01:33.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-04-17" firstname="Andrzej" gender="M" lastname="Skorykow" nation="POL" athleteid="2951">
              <RESULTS>
                <RESULT eventid="1105" points="880" reactiontime="+69" swimtime="00:00:28.41" resultid="2952" heatid="7971" lane="3" entrytime="00:00:28.00" />
                <RESULT eventid="1258" status="DNS" swimtime="00:00:00.00" resultid="2953" heatid="8017" lane="7" entrytime="00:02:30.00" />
                <RESULT comment="Rekord Polski Masters" eventid="1462" points="888" reactiontime="+72" swimtime="00:01:03.27" resultid="2954" heatid="8085" lane="4" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="725" reactiontime="+76" swimtime="00:02:12.83" resultid="2955" heatid="8101" lane="5" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="100" swimtime="00:01:05.50" />
                    <SPLIT distance="150" swimtime="00:01:40.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-06-13" firstname="Agnieszka" gender="F" lastname="Mazurkiewicz" nation="POL" athleteid="2940">
              <RESULTS>
                <RESULT eventid="1090" points="448" reactiontime="+91" swimtime="00:00:38.29" resultid="2941" heatid="7958" lane="0" entrytime="00:00:37.27" />
                <RESULT eventid="1181" points="407" reactiontime="+82" swimtime="00:01:19.52" resultid="2942" heatid="7976" lane="7" entrytime="00:01:18.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="322" reactiontime="+88" swimtime="00:01:35.47" resultid="2943" heatid="8079" lane="3" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="383" reactiontime="+85" swimtime="00:02:56.03" resultid="2944" heatid="8090" lane="1" entrytime="00:02:54.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.48" />
                    <SPLIT distance="100" swimtime="00:01:25.04" />
                    <SPLIT distance="150" swimtime="00:02:11.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-02-29" firstname="Jan" gender="M" lastname="Boboli" nation="POL" athleteid="2796">
              <RESULTS>
                <RESULT eventid="1105" points="418" reactiontime="+99" swimtime="00:00:40.82" resultid="2797" heatid="7964" lane="0" entrytime="00:00:39.00" />
                <RESULT eventid="1198" points="378" reactiontime="+90" swimtime="00:01:31.24" resultid="2798" heatid="7982" lane="2" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="412" reactiontime="+82" swimtime="00:00:38.68" resultid="2799" heatid="8054" lane="1" entrytime="00:00:37.00" />
                <RESULT eventid="1539" points="179" reactiontime="+73" swimtime="00:00:59.37" resultid="2800" heatid="8109" lane="2" entrytime="00:00:56.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-10-03" firstname="Ryszard" gender="M" lastname="Sielski" nation="POL" athleteid="2768">
              <RESULTS>
                <RESULT eventid="1075" points="158" reactiontime="+117" swimtime="00:05:46.16" resultid="2769" heatid="7945" lane="7" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:34.16" />
                    <SPLIT distance="100" swimtime="00:02:58.64" />
                    <SPLIT distance="150" swimtime="00:04:31.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="141" reactiontime="+113" swimtime="00:01:10.44" resultid="2770" heatid="7962" lane="8" entrytime="00:01:25.00" />
                <RESULT eventid="1228" points="293" reactiontime="+111" swimtime="00:00:59.52" resultid="2771" heatid="8000" lane="6" entrytime="00:01:10.00" />
                <RESULT eventid="1288" points="207" reactiontime="+77" swimtime="00:05:26.95" resultid="2772" heatid="8023" lane="9" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.45" />
                    <SPLIT distance="100" swimtime="00:02:42.67" />
                    <SPLIT distance="150" swimtime="00:04:02.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="204" reactiontime="+76" swimtime="00:02:31.87" resultid="2773" heatid="8036" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="274" reactiontime="+118" swimtime="00:05:13.98" resultid="2774" heatid="8071" lane="7" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.99" />
                    <SPLIT distance="100" swimtime="00:02:26.10" />
                    <SPLIT distance="150" swimtime="00:03:51.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="189" reactiontime="+75" swimtime="00:01:10.00" resultid="2775" heatid="8108" lane="4" entrytime="00:01:20.00" />
                <RESULT eventid="1569" points="239" reactiontime="+118" swimtime="00:02:24.78" resultid="2776" heatid="8125" lane="0" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-10-02" firstname="Andrzej" gender="M" lastname="Wiszniewski" nation="POL" athleteid="2832">
              <RESULTS>
                <RESULT eventid="1075" points="229" reactiontime="+99" swimtime="00:03:55.65" resultid="2833" heatid="7946" lane="2" entrytime="00:03:56.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.67" />
                    <SPLIT distance="100" swimtime="00:02:10.40" />
                    <SPLIT distance="150" swimtime="00:03:07.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="137" reactiontime="+103" swimtime="00:00:53.79" resultid="2834" heatid="7962" lane="3" entrytime="00:00:53.30" />
                <RESULT eventid="1258" points="221" reactiontime="+101" swimtime="00:04:10.53" resultid="2835" heatid="8014" lane="4" entrytime="00:04:15.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.93" />
                    <SPLIT distance="100" swimtime="00:02:03.60" />
                    <SPLIT distance="150" swimtime="00:03:07.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="136" reactiontime="+94" swimtime="00:04:48.63" resultid="2836" heatid="8023" lane="6" entrytime="00:04:23.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.05" />
                    <SPLIT distance="100" swimtime="00:02:25.11" />
                    <SPLIT distance="150" swimtime="00:03:42.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="139" reactiontime="+85" swimtime="00:02:07.11" resultid="2837" heatid="8036" lane="4" entrytime="00:02:10.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1402" points="379" reactiontime="+95" swimtime="00:03:41.07" resultid="2838" heatid="8072" lane="2" entrytime="00:03:54.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.76" />
                    <SPLIT distance="100" swimtime="00:01:47.52" />
                    <SPLIT distance="150" swimtime="00:02:44.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="356" reactiontime="+97" swimtime="00:01:42.24" resultid="2839" heatid="8125" lane="5" entrytime="00:01:56.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="264" reactiontime="+102" swimtime="00:08:16.25" resultid="2840" heatid="8167" lane="4" entrytime="00:08:25.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.98" />
                    <SPLIT distance="100" swimtime="00:02:11.05" />
                    <SPLIT distance="150" swimtime="00:03:26.22" />
                    <SPLIT distance="200" swimtime="00:04:41.16" />
                    <SPLIT distance="250" swimtime="00:05:38.24" />
                    <SPLIT distance="300" swimtime="00:06:34.60" />
                    <SPLIT distance="350" swimtime="00:07:26.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-05" firstname="Bartłomiej" gender="M" lastname="Pawłowski" nation="POL" athleteid="2801">
              <RESULTS>
                <RESULT eventid="1228" points="614" reactiontime="+77" swimtime="00:00:35.88" resultid="2802" heatid="8008" lane="8" entrytime="00:00:35.00" />
                <RESULT eventid="1372" points="636" reactiontime="+83" swimtime="00:00:28.57" resultid="2803" heatid="8060" lane="5" entrytime="00:00:28.38" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-08-12" firstname="Jakub" gender="M" lastname="Szulc" nation="POL" athleteid="2903">
              <RESULTS>
                <RESULT eventid="1105" points="534" reactiontime="+71" swimtime="00:00:31.44" resultid="2904" heatid="7968" lane="6" entrytime="00:00:31.00" />
                <RESULT eventid="1135" points="559" reactiontime="+83" swimtime="00:10:49.76" resultid="2905" heatid="8139" lane="9" entrytime="00:11:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                    <SPLIT distance="100" swimtime="00:01:13.02" />
                    <SPLIT distance="150" swimtime="00:01:52.59" />
                    <SPLIT distance="200" swimtime="00:02:33.07" />
                    <SPLIT distance="250" swimtime="00:03:14.12" />
                    <SPLIT distance="300" swimtime="00:03:55.25" />
                    <SPLIT distance="350" swimtime="00:04:36.37" />
                    <SPLIT distance="400" swimtime="00:05:17.62" />
                    <SPLIT distance="450" swimtime="00:05:59.25" />
                    <SPLIT distance="500" swimtime="00:06:41.52" />
                    <SPLIT distance="550" swimtime="00:07:23.65" />
                    <SPLIT distance="600" swimtime="00:08:05.51" />
                    <SPLIT distance="650" swimtime="00:08:47.44" />
                    <SPLIT distance="700" swimtime="00:09:29.59" />
                    <SPLIT distance="750" swimtime="00:10:10.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="565" reactiontime="+82" swimtime="00:01:02.86" resultid="2906" heatid="7988" lane="0" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="559" reactiontime="+77" swimtime="00:00:28.55" resultid="2907" heatid="8059" lane="0" entrytime="00:00:29.00" />
                <RESULT eventid="1509" points="554" reactiontime="+74" swimtime="00:02:20.79" resultid="2909" heatid="8100" lane="0" entrytime="00:02:24.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                    <SPLIT distance="100" swimtime="00:01:07.36" />
                    <SPLIT distance="150" swimtime="00:01:43.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="575" reactiontime="+84" swimtime="00:05:08.33" resultid="8292" heatid="8156" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                    <SPLIT distance="100" swimtime="00:01:11.31" />
                    <SPLIT distance="150" swimtime="00:01:49.97" />
                    <SPLIT distance="200" swimtime="00:02:29.83" />
                    <SPLIT distance="250" swimtime="00:03:10.53" />
                    <SPLIT distance="300" swimtime="00:03:50.84" />
                    <SPLIT distance="350" swimtime="00:04:31.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-02-23" firstname="Joanna" gender="F" lastname="Gołębiowska" nation="POL" athleteid="2868">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters" eventid="1181" points="870" reactiontime="+71" swimtime="00:01:01.75" resultid="2869" heatid="7979" lane="3" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.72" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1357" points="885" reactiontime="+75" swimtime="00:00:28.27" resultid="2870" heatid="8050" lane="7" entrytime="00:00:28.80" />
                <RESULT comment="Rekord Polski Masters" eventid="1447" points="923" reactiontime="+71" swimtime="00:01:07.27" resultid="2871" heatid="8080" lane="4" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-06-13" firstname="Marcin" gender="M" lastname="Giejsztowt" nation="POL" athleteid="2863">
              <RESULTS>
                <RESULT eventid="1105" points="492" reactiontime="+82" swimtime="00:00:32.32" resultid="2864" heatid="7966" lane="1" entrytime="00:00:34.45" />
                <RESULT eventid="1198" points="475" reactiontime="+77" swimtime="00:01:06.59" resultid="2865" heatid="7986" lane="9" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="533" reactiontime="+83" swimtime="00:05:16.22" resultid="2866" heatid="8153" lane="1" entrytime="00:05:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.25" />
                    <SPLIT distance="100" swimtime="00:01:14.56" />
                    <SPLIT distance="150" swimtime="00:01:54.01" />
                    <SPLIT distance="200" swimtime="00:02:34.84" />
                    <SPLIT distance="250" swimtime="00:03:15.93" />
                    <SPLIT distance="300" swimtime="00:03:55.79" />
                    <SPLIT distance="350" swimtime="00:04:36.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="496" reactiontime="+80" swimtime="00:02:26.05" resultid="2867" heatid="8099" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                    <SPLIT distance="100" swimtime="00:01:10.64" />
                    <SPLIT distance="150" swimtime="00:01:48.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-30" firstname="Monika" gender="F" lastname="Jarecka-Skorykow" nation="POL" athleteid="2945">
              <RESULTS>
                <RESULT eventid="1090" points="611" reactiontime="+71" swimtime="00:00:35.09" resultid="2946" heatid="7957" lane="5" entrytime="00:00:37.50" />
                <RESULT eventid="1213" points="620" reactiontime="+79" swimtime="00:00:40.99" resultid="2947" heatid="7997" lane="7" entrytime="00:00:43.50" />
                <RESULT eventid="1357" points="625" reactiontime="+74" swimtime="00:00:32.21" resultid="2948" heatid="8047" lane="4" entrytime="00:00:33.50" />
                <RESULT eventid="1387" points="568" reactiontime="+82" swimtime="00:03:25.11" resultid="2949" heatid="8068" lane="4" entrytime="00:03:30.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.96" />
                    <SPLIT distance="100" swimtime="00:01:36.90" />
                    <SPLIT distance="150" swimtime="00:02:30.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="606" reactiontime="+77" swimtime="00:01:30.74" resultid="2950" heatid="8121" lane="6" entrytime="00:01:35.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-04-28" firstname="Paweł" gender="M" lastname="Rogosz" nation="POL" athleteid="2816">
              <RESULTS>
                <RESULT eventid="1075" points="617" reactiontime="+87" swimtime="00:02:38.70" resultid="2817" heatid="7951" lane="5" entrytime="00:02:42.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                    <SPLIT distance="100" swimtime="00:01:17.20" />
                    <SPLIT distance="150" swimtime="00:02:02.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="533" reactiontime="+100" swimtime="00:21:08.11" resultid="2818" heatid="8143" lane="8" entrytime="00:21:35.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.96" />
                    <SPLIT distance="100" swimtime="00:01:20.15" />
                    <SPLIT distance="150" swimtime="00:02:03.10" />
                    <SPLIT distance="200" swimtime="00:02:46.54" />
                    <SPLIT distance="250" swimtime="00:03:29.14" />
                    <SPLIT distance="300" swimtime="00:04:12.10" />
                    <SPLIT distance="350" swimtime="00:04:54.97" />
                    <SPLIT distance="400" swimtime="00:05:37.73" />
                    <SPLIT distance="450" swimtime="00:06:20.61" />
                    <SPLIT distance="500" swimtime="00:07:03.31" />
                    <SPLIT distance="550" swimtime="00:07:45.61" />
                    <SPLIT distance="600" swimtime="00:08:27.86" />
                    <SPLIT distance="650" swimtime="00:09:10.48" />
                    <SPLIT distance="700" swimtime="00:09:52.33" />
                    <SPLIT distance="750" swimtime="00:10:35.14" />
                    <SPLIT distance="800" swimtime="00:11:17.87" />
                    <SPLIT distance="850" swimtime="00:12:00.45" />
                    <SPLIT distance="900" swimtime="00:12:43.16" />
                    <SPLIT distance="950" swimtime="00:13:25.53" />
                    <SPLIT distance="1000" swimtime="00:14:08.07" />
                    <SPLIT distance="1050" swimtime="00:14:51.27" />
                    <SPLIT distance="1100" swimtime="00:15:33.49" />
                    <SPLIT distance="1150" swimtime="00:16:17.38" />
                    <SPLIT distance="1200" swimtime="00:16:59.65" />
                    <SPLIT distance="1250" swimtime="00:17:43.16" />
                    <SPLIT distance="1300" swimtime="00:18:25.56" />
                    <SPLIT distance="1350" swimtime="00:19:08.39" />
                    <SPLIT distance="1400" swimtime="00:19:50.26" />
                    <SPLIT distance="1450" swimtime="00:20:31.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="467" reactiontime="+92" swimtime="00:01:06.99" resultid="2819" heatid="7989" lane="0" entrytime="00:01:04.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="511" reactiontime="+97" swimtime="00:02:48.29" resultid="2820" heatid="8016" lane="5" entrytime="00:02:49.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.07" />
                    <SPLIT distance="100" swimtime="00:01:20.45" />
                    <SPLIT distance="150" swimtime="00:02:03.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Mirosław" gender="M" lastname="Warchoł" nation="POL" athleteid="2963">
              <RESULTS>
                <RESULT eventid="1075" points="954" reactiontime="+86" swimtime="00:02:44.89" resultid="2964" heatid="7950" lane="3" entrytime="00:02:51.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                    <SPLIT distance="100" swimtime="00:01:15.42" />
                    <SPLIT distance="150" swimtime="00:02:08.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="1094" reactiontime="+86" swimtime="00:02:44.24" resultid="2965" heatid="8026" lane="0" entrytime="00:02:52.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                    <SPLIT distance="100" swimtime="00:01:19.62" />
                    <SPLIT distance="150" swimtime="00:02:01.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="910" reactiontime="+75" swimtime="00:01:16.99" resultid="2966" heatid="8041" lane="9" entrytime="00:01:16.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="824" reactiontime="+68" swimtime="00:00:29.15" resultid="2967" heatid="8058" lane="9" entrytime="00:00:29.99" />
                <RESULT eventid="1509" points="966" reactiontime="+71" swimtime="00:02:23.34" resultid="2968" heatid="8100" lane="9" entrytime="00:02:24.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.52" />
                    <SPLIT distance="100" swimtime="00:01:09.85" />
                    <SPLIT distance="150" swimtime="00:01:46.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-06-07" firstname="Olga" gender="F" lastname="Krysiak" nation="POL" athleteid="2846">
              <RESULTS>
                <RESULT eventid="1090" points="531" reactiontime="+76" swimtime="00:00:34.42" resultid="2847" heatid="7959" lane="5" entrytime="00:00:34.30" />
                <RESULT eventid="1181" points="690" reactiontime="+74" swimtime="00:01:06.39" resultid="2848" heatid="7979" lane="1" entrytime="00:01:03.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="2849" heatid="8018" lane="1" />
                <RESULT eventid="1357" points="702" reactiontime="+71" swimtime="00:00:29.94" resultid="2850" heatid="8050" lane="8" entrytime="00:00:29.00" />
                <RESULT eventid="1417" points="557" reactiontime="+84" swimtime="00:05:26.31" resultid="2851" heatid="8147" lane="8" entrytime="00:05:30.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.90" />
                    <SPLIT distance="100" swimtime="00:01:16.52" />
                    <SPLIT distance="150" swimtime="00:01:58.64" />
                    <SPLIT distance="200" swimtime="00:02:41.26" />
                    <SPLIT distance="250" swimtime="00:03:23.45" />
                    <SPLIT distance="300" swimtime="00:04:06.13" />
                    <SPLIT distance="350" swimtime="00:04:47.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="598" reactiontime="+75" swimtime="00:02:32.09" resultid="2852" heatid="8092" lane="0" entrytime="00:02:25.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                    <SPLIT distance="100" swimtime="00:01:11.88" />
                    <SPLIT distance="150" swimtime="00:01:52.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-11-05" firstname="Mirosława" gender="F" lastname="Przyłuska" nation="POL" athleteid="2827">
              <RESULTS>
                <RESULT eventid="1213" points="262" reactiontime="+97" swimtime="00:01:00.07" resultid="2828" heatid="7995" lane="2" entrytime="00:00:56.00" />
                <RESULT eventid="1387" points="314" reactiontime="+98" swimtime="00:04:48.31" resultid="2829" heatid="8067" lane="7" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.72" />
                    <SPLIT distance="100" swimtime="00:02:21.28" />
                    <SPLIT distance="150" swimtime="00:03:38.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="195" reactiontime="+89" swimtime="00:04:34.05" resultid="2830" heatid="8087" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.27" />
                    <SPLIT distance="100" swimtime="00:02:11.54" />
                    <SPLIT distance="150" swimtime="00:03:23.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="300" reactiontime="+105" swimtime="00:02:14.23" resultid="2831" heatid="8119" lane="3" entrytime="00:01:56.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-05" firstname="Rafał" gender="M" lastname="Skośkiewicz" nation="POL" athleteid="2809">
              <RESULTS>
                <RESULT eventid="1075" points="833" reactiontime="+80" swimtime="00:02:34.99" resultid="2810" heatid="7947" lane="5" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                    <SPLIT distance="100" swimtime="00:01:11.61" />
                    <SPLIT distance="150" swimtime="00:01:59.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="692" reactiontime="+86" swimtime="00:00:30.78" resultid="2811" heatid="7968" lane="0" entrytime="00:00:32.00" />
                <RESULT eventid="1288" points="748" reactiontime="+77" swimtime="00:02:35.99" resultid="2812" heatid="8027" lane="6" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.87" />
                    <SPLIT distance="100" swimtime="00:01:14.83" />
                    <SPLIT distance="150" swimtime="00:01:54.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="710" reactiontime="+77" swimtime="00:01:11.60" resultid="2813" heatid="8042" lane="4" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="631" reactiontime="+82" swimtime="00:02:19.15" resultid="2814" heatid="8099" lane="4" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                    <SPLIT distance="100" swimtime="00:01:08.34" />
                    <SPLIT distance="150" swimtime="00:01:44.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="663" reactiontime="+79" swimtime="00:00:33.52" resultid="2815" heatid="8116" lane="9" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-10-19" firstname="Emilia" gender="F" lastname="Sączyńska" nation="POL" athleteid="2924">
              <RESULTS>
                <RESULT eventid="1273" points="593" reactiontime="+77" swimtime="00:02:54.79" resultid="2925" heatid="8021" lane="8" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.76" />
                    <SPLIT distance="100" swimtime="00:01:24.15" />
                    <SPLIT distance="150" swimtime="00:02:10.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="592" reactiontime="+76" swimtime="00:01:20.69" resultid="2926" heatid="8034" lane="4" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="434" reactiontime="+93" swimtime="00:01:24.70" resultid="2927" heatid="8080" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="533" reactiontime="+76" swimtime="00:00:38.35" resultid="2928" heatid="8107" lane="9" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-05-10" firstname="Katarzyna" gender="F" lastname="Czarnecka" nation="POL" athleteid="2919">
              <RESULTS>
                <RESULT eventid="1213" points="456" swimtime="00:00:42.41" resultid="2920" heatid="7998" lane="7" entrytime="00:00:41.27" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="2921" heatid="8018" lane="7" />
                <RESULT eventid="1387" points="478" reactiontime="+81" swimtime="00:03:25.15" resultid="2922" heatid="8066" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.89" />
                    <SPLIT distance="100" swimtime="00:01:40.67" />
                    <SPLIT distance="150" swimtime="00:02:33.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="482" reactiontime="+71" swimtime="00:01:33.21" resultid="2923" heatid="8118" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-24" firstname="Jan" gender="M" lastname="Pfitzner" nation="POL" athleteid="2821">
              <RESULTS>
                <RESULT eventid="1198" points="667" reactiontime="+73" swimtime="00:00:59.16" resultid="2822" heatid="7992" lane="0" entrytime="00:00:58.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="645" reactiontime="+78" swimtime="00:00:26.79" resultid="2823" heatid="8063" lane="7" entrytime="00:00:26.83" />
                <RESULT eventid="1462" points="515" reactiontime="+70" swimtime="00:01:10.91" resultid="2824" heatid="8085" lane="2" entrytime="00:01:08.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="611" reactiontime="+72" swimtime="00:02:15.67" resultid="2825" heatid="8102" lane="9" entrytime="00:02:12.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                    <SPLIT distance="100" swimtime="00:01:08.02" />
                    <SPLIT distance="150" swimtime="00:01:42.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="606" reactiontime="+83" swimtime="00:00:31.63" resultid="2826" heatid="8116" lane="1" entrytime="00:00:31.64" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-11-10" firstname="Anna" gender="F" lastname="Turczyn" nation="POL" athleteid="2935">
              <RESULTS>
                <RESULT eventid="1181" points="200" reactiontime="+97" swimtime="00:01:40.46" resultid="2936" heatid="7975" lane="7" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="264" swimtime="00:00:50.89" resultid="2937" heatid="7996" lane="7" entrytime="00:00:48.00" />
                <RESULT eventid="1357" points="239" reactiontime="+93" swimtime="00:00:43.56" resultid="2938" heatid="8046" lane="0" entrytime="00:00:38.00" />
                <RESULT comment="O4 - Start wykonany przed sygnałem (przedwczesny start)" eventid="1524" reactiontime="+58" status="DSQ" swimtime="00:00:51.34" resultid="2939" heatid="8105" lane="8" entrytime="00:00:46.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-06-16" firstname="Paweł" gender="M" lastname="Witkowski" nation="POL" athleteid="2841">
              <RESULTS>
                <RESULT eventid="1228" points="701" reactiontime="+82" swimtime="00:00:32.85" resultid="2842" heatid="8010" lane="0" entrytime="00:00:32.45" />
                <RESULT eventid="1372" points="524" reactiontime="+89" swimtime="00:00:28.83" resultid="2843" heatid="8055" lane="3" entrytime="00:00:32.50" />
                <RESULT eventid="1402" points="621" reactiontime="+93" swimtime="00:02:51.55" resultid="2844" heatid="8076" lane="1" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.78" />
                    <SPLIT distance="100" swimtime="00:01:24.10" />
                    <SPLIT distance="150" swimtime="00:02:08.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="634" reactiontime="+87" swimtime="00:01:15.81" resultid="2845" heatid="8131" lane="6" entrytime="00:01:15.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-02-15" firstname="Manuela" gender="F" lastname="Nawrocka" nation="POL" athleteid="2782">
              <RESULTS>
                <RESULT eventid="1058" points="689" reactiontime="+86" swimtime="00:02:44.57" resultid="2783" heatid="7944" lane="3" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                    <SPLIT distance="100" swimtime="00:01:17.27" />
                    <SPLIT distance="150" swimtime="00:02:05.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="564" swimtime="00:00:39.50" resultid="2784" heatid="7998" lane="4" entrytime="00:00:40.50" />
                <RESULT eventid="1387" points="588" reactiontime="+86" swimtime="00:03:05.92" resultid="2785" heatid="8070" lane="2" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.79" />
                    <SPLIT distance="100" swimtime="00:01:27.84" />
                    <SPLIT distance="150" swimtime="00:02:16.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1447" points="472" reactiontime="+85" swimtime="00:01:22.40" resultid="2786" heatid="8079" lane="4" entrytime="00:01:22.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="602" reactiontime="+84" swimtime="00:01:25.68" resultid="2787" heatid="8123" lane="0" entrytime="00:01:28.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-30" firstname="Monika" gender="F" lastname="Jarecka - Skorykow" nation="POL" athleteid="6001" />
            <ATHLETE birthdate="1949-07-26" firstname="Anna" gender="F" lastname="Szemberg" nation="POL" athleteid="2887">
              <RESULTS>
                <RESULT eventid="1120" points="381" reactiontime="+78" swimtime="00:17:05.74" resultid="2888" heatid="8137" lane="4" entrytime="00:16:55.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.32" />
                    <SPLIT distance="100" swimtime="00:01:57.15" />
                    <SPLIT distance="150" swimtime="00:03:02.97" />
                    <SPLIT distance="200" swimtime="00:04:09.30" />
                    <SPLIT distance="250" swimtime="00:05:15.24" />
                    <SPLIT distance="300" swimtime="00:06:21.32" />
                    <SPLIT distance="350" swimtime="00:07:25.83" />
                    <SPLIT distance="400" swimtime="00:08:29.99" />
                    <SPLIT distance="450" swimtime="00:09:33.31" />
                    <SPLIT distance="500" swimtime="00:10:37.72" />
                    <SPLIT distance="550" swimtime="00:11:41.70" />
                    <SPLIT distance="600" swimtime="00:12:46.50" />
                    <SPLIT distance="650" swimtime="00:13:51.18" />
                    <SPLIT distance="700" swimtime="00:14:56.22" />
                    <SPLIT distance="750" swimtime="00:16:00.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="216" reactiontime="+78" swimtime="00:01:59.82" resultid="2889" heatid="7973" lane="4" entrytime="00:01:55.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="220" swimtime="00:01:08.76" resultid="2890" heatid="7995" lane="9" entrytime="00:01:06.89" />
                <RESULT eventid="1357" points="284" reactiontime="+80" swimtime="00:00:49.43" resultid="2891" heatid="8044" lane="4" entrytime="00:00:50.02" />
                <RESULT eventid="1417" points="336" swimtime="00:08:38.37" resultid="2892" heatid="8149" lane="9" entrytime="00:08:16.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.04" />
                    <SPLIT distance="100" swimtime="00:01:59.89" />
                    <SPLIT distance="150" swimtime="00:03:07.30" />
                    <SPLIT distance="200" swimtime="00:04:15.49" />
                    <SPLIT distance="250" swimtime="00:05:22.67" />
                    <SPLIT distance="300" swimtime="00:06:29.19" />
                    <SPLIT distance="350" swimtime="00:07:34.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="265" swimtime="00:04:12.31" resultid="2893" heatid="8087" lane="3" entrytime="00:04:04.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.34" />
                    <SPLIT distance="100" swimtime="00:02:01.39" />
                    <SPLIT distance="150" swimtime="00:03:07.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-06-17" firstname="Leszek" gender="M" lastname="Madej" nation="POL" athleteid="2763">
              <RESULTS>
                <RESULT eventid="1198" points="1086" reactiontime="+79" swimtime="00:00:59.11" resultid="2764" heatid="7991" lane="3" entrytime="00:00:59.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="697" swimtime="00:00:35.02" resultid="2765" heatid="8007" lane="1" entrytime="00:00:36.52" />
                <RESULT eventid="1509" points="1120" reactiontime="+77" swimtime="00:02:11.08" resultid="2766" heatid="8101" lane="3" entrytime="00:02:13.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                    <SPLIT distance="100" swimtime="00:01:02.98" />
                    <SPLIT distance="150" swimtime="00:01:35.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="810" reactiontime="+78" swimtime="00:01:18.15" resultid="2767" heatid="8130" lane="2" entrytime="00:01:20.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Anna" gender="M" lastname="Kotusińska" nation="POL" athleteid="6003" />
            <ATHLETE birthdate="1983-06-10" firstname="Tomasz" gender="M" lastname="Porada" nation="POL" athleteid="2788">
              <RESULTS>
                <RESULT eventid="1075" points="643" reactiontime="+76" swimtime="00:02:32.44" resultid="2789" heatid="7952" lane="2" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                    <SPLIT distance="100" swimtime="00:01:14.35" />
                    <SPLIT distance="150" swimtime="00:01:56.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="494" swimtime="00:10:17.90" resultid="2790" heatid="8141" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.63" />
                    <SPLIT distance="100" swimtime="00:01:09.20" />
                    <SPLIT distance="150" swimtime="00:01:47.19" />
                    <SPLIT distance="200" swimtime="00:02:25.28" />
                    <SPLIT distance="250" swimtime="00:03:03.95" />
                    <SPLIT distance="300" swimtime="00:03:42.94" />
                    <SPLIT distance="350" swimtime="00:04:22.25" />
                    <SPLIT distance="400" swimtime="00:05:01.64" />
                    <SPLIT distance="450" swimtime="00:05:41.41" />
                    <SPLIT distance="500" swimtime="00:06:20.91" />
                    <SPLIT distance="550" swimtime="00:07:01.09" />
                    <SPLIT distance="600" swimtime="00:07:40.19" />
                    <SPLIT distance="650" swimtime="00:08:19.60" />
                    <SPLIT distance="700" swimtime="00:08:59.33" />
                    <SPLIT distance="750" swimtime="00:09:39.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="615" reactiontime="+74" swimtime="00:00:34.31" resultid="2791" heatid="8008" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1402" points="728" reactiontime="+78" swimtime="00:02:42.76" resultid="2792" heatid="8077" lane="9" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.00" />
                    <SPLIT distance="100" swimtime="00:01:18.26" />
                    <SPLIT distance="150" swimtime="00:02:00.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="613" reactiontime="+81" swimtime="00:04:52.53" resultid="2793" heatid="8156" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                    <SPLIT distance="100" swimtime="00:01:07.55" />
                    <SPLIT distance="150" swimtime="00:01:44.28" />
                    <SPLIT distance="200" swimtime="00:02:21.41" />
                    <SPLIT distance="250" swimtime="00:02:58.93" />
                    <SPLIT distance="300" swimtime="00:03:36.87" />
                    <SPLIT distance="350" swimtime="00:04:15.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="671" reactiontime="+72" swimtime="00:01:14.41" resultid="2794" heatid="8131" lane="2" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="569" reactiontime="+80" swimtime="00:05:30.43" resultid="2795" heatid="8167" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                    <SPLIT distance="100" swimtime="00:01:14.69" />
                    <SPLIT distance="150" swimtime="00:02:02.27" />
                    <SPLIT distance="200" swimtime="00:02:48.19" />
                    <SPLIT distance="250" swimtime="00:03:31.59" />
                    <SPLIT distance="300" swimtime="00:04:15.91" />
                    <SPLIT distance="350" swimtime="00:04:54.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-10-20" firstname="Norbert" gender="M" lastname="Stablewski" nation="POL" athleteid="2876">
              <RESULTS>
                <RESULT eventid="1372" points="522" reactiontime="+89" swimtime="00:00:30.52" resultid="2877" heatid="8058" lane="1" entrytime="00:00:29.50" />
                <RESULT eventid="1509" points="406" reactiontime="+89" swimtime="00:02:39.93" resultid="2878" heatid="8097" lane="2" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.15" />
                    <SPLIT distance="100" swimtime="00:01:19.46" />
                    <SPLIT distance="150" swimtime="00:02:01.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-13" firstname="Stanisław" gender="M" lastname="Kozak" nation="POL" athleteid="2872">
              <RESULTS>
                <RESULT eventid="1228" points="759" reactiontime="+76" swimtime="00:00:32.11" resultid="2873" heatid="8009" lane="8" entrytime="00:00:33.50" />
                <RESULT eventid="1402" points="622" reactiontime="+91" swimtime="00:02:51.39" resultid="2874" heatid="8076" lane="2" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.90" />
                    <SPLIT distance="100" swimtime="00:01:24.91" />
                    <SPLIT distance="150" swimtime="00:02:09.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="663" reactiontime="+78" swimtime="00:01:14.16" resultid="2875" heatid="8131" lane="3" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-08-02" firstname="Tomasz" gender="M" lastname="Jąkalski" nation="POL" athleteid="2894">
              <RESULTS>
                <RESULT eventid="1228" status="DNS" swimtime="00:00:00.00" resultid="2895" heatid="8000" lane="0" />
                <RESULT eventid="1288" points="464" reactiontime="+63" swimtime="00:02:39.82" resultid="2896" heatid="8024" lane="9" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                    <SPLIT distance="100" swimtime="00:01:14.86" />
                    <SPLIT distance="150" swimtime="00:01:57.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="625" reactiontime="+62" swimtime="00:01:09.29" resultid="2897" heatid="8043" lane="9" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="595" reactiontime="+82" swimtime="00:01:07.59" resultid="2898" heatid="8085" lane="6" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="655" reactiontime="+64" swimtime="00:00:30.83" resultid="2899" heatid="8116" lane="3" entrytime="00:00:30.49" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Anna" gender="F" lastname="Kotusińska" nation="POL" athleteid="2900">
              <RESULTS>
                <RESULT eventid="1181" points="353" reactiontime="+89" swimtime="00:01:23.12" resultid="2901" heatid="7976" lane="6" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="477" reactiontime="+84" swimtime="00:00:34.61" resultid="2902" heatid="8047" lane="0" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-10-04" firstname="Maciej" gender="M" lastname="Szymański" nation="POL" athleteid="6432">
              <RESULTS>
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="6433" heatid="7993" lane="3" entrytime="00:00:55.50" />
                <RESULT eventid="1372" status="DNS" swimtime="00:00:00.00" resultid="6434" heatid="8065" lane="7" entrytime="00:00:24.82" />
                <RESULT eventid="1462" status="DNS" swimtime="00:00:00.00" resultid="6435" heatid="8086" lane="0" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-02-15" firstname="Manuela" gender="M" lastname="Nawrocka" nation="POL" athleteid="6002" />
            <ATHLETE birthdate="1988-05-24" firstname="Marlena" gender="F" lastname="Dobrasiewicz" nation="POL" athleteid="2929">
              <RESULTS>
                <RESULT eventid="1181" points="723" reactiontime="+81" swimtime="00:01:05.45" resultid="2930" heatid="7979" lane="8" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="596" reactiontime="+80" swimtime="00:00:38.79" resultid="2931" heatid="7999" lane="8" entrytime="00:00:39.50" />
                <RESULT eventid="1387" points="653" reactiontime="+89" swimtime="00:02:59.53" resultid="2932" heatid="8070" lane="3" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.32" />
                    <SPLIT distance="100" swimtime="00:01:25.81" />
                    <SPLIT distance="150" swimtime="00:02:12.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="680" reactiontime="+90" swimtime="00:02:26.60" resultid="2933" heatid="8092" lane="8" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                    <SPLIT distance="100" swimtime="00:01:10.95" />
                    <SPLIT distance="150" swimtime="00:01:49.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="611" reactiontime="+88" swimtime="00:01:25.26" resultid="2934" heatid="8123" lane="7" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-08-01" firstname="Edyta" gender="F" lastname="Olszewska" nation="POL" athleteid="2859">
              <RESULTS>
                <RESULT eventid="1213" points="694" swimtime="00:00:42.63" resultid="2860" heatid="7998" lane="2" entrytime="00:00:41.06" />
                <RESULT eventid="1387" points="747" reactiontime="+81" swimtime="00:03:21.91" resultid="2861" heatid="8070" lane="7" entrytime="00:03:14.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.78" />
                    <SPLIT distance="100" swimtime="00:01:40.49" />
                    <SPLIT distance="150" swimtime="00:02:31.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="673" reactiontime="+75" swimtime="00:01:35.22" resultid="2862" heatid="8122" lane="2" entrytime="00:01:30.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-05-18" firstname="Barbara" gender="F" lastname="Łowkis" nation="POL" athleteid="2804">
              <RESULTS>
                <RESULT eventid="1181" points="381" reactiontime="+122" swimtime="00:01:39.27" resultid="2805" heatid="7974" lane="8" entrytime="00:01:43.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="558" reactiontime="+84" swimtime="00:01:49.58" resultid="2806" heatid="8033" lane="8" entrytime="00:01:53.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="571" reactiontime="+110" swimtime="00:00:39.19" resultid="2807" heatid="8045" lane="7" entrytime="00:00:43.59" />
                <RESULT eventid="1524" points="661" reactiontime="+101" swimtime="00:00:46.66" resultid="2808" heatid="8104" lane="3" entrytime="00:00:50.70" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="M" number="3">
              <RESULTS>
                <RESULT comment="O4 - Start wykonany przed sygnałem (przedwczesny start)" eventid="1318" reactiontime="+73" status="DSQ" swimtime="00:03:56.91" resultid="2978" heatid="8031" lane="5" entrytime="00:03:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.83" />
                    <SPLIT distance="100" swimtime="00:00:58.14" />
                    <SPLIT distance="150" swimtime="00:01:26.65" />
                    <SPLIT distance="200" swimtime="00:01:59.36" />
                    <SPLIT distance="250" swimtime="00:02:27.41" />
                    <SPLIT distance="300" swimtime="00:02:59.46" />
                    <SPLIT distance="350" swimtime="00:03:25.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2821" number="1" reactiontime="+73" status="DSQ" />
                    <RELAYPOSITION athleteid="2788" number="2" reactiontime="+42" status="DSQ" />
                    <RELAYPOSITION athleteid="2894" number="3" reactiontime="+34" status="DSQ" />
                    <RELAYPOSITION athleteid="2879" number="4" reactiontime="-8" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" number="4">
              <RESULTS>
                <RESULT comment="Rekord Polski" eventid="1318" reactiontime="+72" swimtime="00:03:57.53" resultid="2979" heatid="8031" lane="3" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.51" />
                    <SPLIT distance="100" swimtime="00:00:59.05" />
                    <SPLIT distance="150" swimtime="00:01:26.29" />
                    <SPLIT distance="200" swimtime="00:01:54.87" />
                    <SPLIT distance="250" swimtime="00:02:22.89" />
                    <SPLIT distance="300" swimtime="00:02:53.55" />
                    <SPLIT distance="350" swimtime="00:03:24.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2951" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="2777" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="2763" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="2963" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="1318" reactiontime="+86" swimtime="00:04:23.50" resultid="2980" heatid="8031" lane="9" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.06" />
                    <SPLIT distance="100" swimtime="00:01:05.39" />
                    <SPLIT distance="150" swimtime="00:01:36.84" />
                    <SPLIT distance="200" swimtime="00:02:11.38" />
                    <SPLIT distance="250" swimtime="00:02:43.78" />
                    <SPLIT distance="300" swimtime="00:03:20.19" />
                    <SPLIT distance="350" swimtime="00:03:50.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2872" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="2816" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="2876" number="3" reactiontime="+72" />
                    <RELAYPOSITION athleteid="2903" number="4" reactiontime="+50" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1303" reactiontime="+89" swimtime="00:05:11.71" resultid="2976" heatid="8029" lane="0" entrytime="00:05:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.09" />
                    <SPLIT distance="100" swimtime="00:01:19.93" />
                    <SPLIT distance="150" swimtime="00:01:57.68" />
                    <SPLIT distance="200" swimtime="00:02:40.04" />
                    <SPLIT distance="250" swimtime="00:03:15.64" />
                    <SPLIT distance="300" swimtime="00:03:56.45" />
                    <SPLIT distance="350" swimtime="00:04:31.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2900" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="2940" number="2" reactiontime="+65" />
                    <RELAYPOSITION athleteid="2919" number="3" reactiontime="+65" />
                    <RELAYPOSITION athleteid="2924" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1303" reactiontime="+86" swimtime="00:04:22.70" resultid="2977" heatid="8029" lane="3" entrytime="00:04:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.80" />
                    <SPLIT distance="100" swimtime="00:01:05.78" />
                    <SPLIT distance="150" swimtime="00:01:36.66" />
                    <SPLIT distance="200" swimtime="00:02:12.18" />
                    <SPLIT distance="250" swimtime="00:02:42.93" />
                    <SPLIT distance="300" swimtime="00:03:16.50" />
                    <SPLIT distance="350" swimtime="00:03:47.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2929" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="2782" number="2" reactiontime="+70" />
                    <RELAYPOSITION athleteid="2956" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="2868" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="6">
              <RESULTS>
                <RESULT eventid="1614" reactiontime="+76" swimtime="00:02:12.62" resultid="6004" heatid="8135" lane="2" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                    <SPLIT distance="100" swimtime="00:01:12.63" />
                    <SPLIT distance="150" swimtime="00:01:45.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2809" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="6001" number="2" />
                    <RELAYPOSITION athleteid="2929" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="2763" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="X" number="7">
              <RESULTS>
                <RESULT eventid="1614" reactiontime="+69" swimtime="00:02:08.92" resultid="6005" heatid="8135" lane="4" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                    <SPLIT distance="100" swimtime="00:01:11.57" />
                    <SPLIT distance="150" swimtime="00:01:39.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2894" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="2919" number="2" />
                    <RELAYPOSITION athleteid="2879" number="3" reactiontime="+29" />
                    <RELAYPOSITION athleteid="6002" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" number="8">
              <RESULTS>
                <RESULT eventid="1614" reactiontime="+74" swimtime="00:02:18.74" resultid="6006" heatid="8134" lane="6" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                    <SPLIT distance="100" swimtime="00:01:11.31" />
                    <SPLIT distance="150" swimtime="00:01:43.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2924" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="2841" number="2" />
                    <RELAYPOSITION athleteid="2863" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="2940" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="X" number="9">
              <RESULTS>
                <RESULT eventid="1614" reactiontime="+77" swimtime="00:02:09.42" resultid="6007" heatid="8135" lane="7" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                    <SPLIT distance="100" swimtime="00:01:03.43" />
                    <SPLIT distance="150" swimtime="00:01:35.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2821" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="2872" number="2" />
                    <RELAYPOSITION athleteid="2956" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="6003" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5108" name="Weteran Zabrze">
          <CONTACT city="ZABRZE" email="weteranzabrze@op.pl" name="BO9SOWSKI  WŁODZIMIERZ" street="ŚW.JANA  4A/4" zip="41803" />
          <ATHLETES>
            <ATHLETE birthdate="1943-03-12" firstname="Krystyna" gender="F" lastname="Fecica" nation="POL" license="502611100002" athleteid="5133">
              <RESULTS>
                <RESULT comment="Rekord Polski Masters, Rekord Polski" eventid="1150" points="767" reactiontime="+109" swimtime="00:31:30.18" resultid="5134" heatid="8142" lane="8" entrytime="00:31:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.03" />
                    <SPLIT distance="100" swimtime="00:01:57.67" />
                    <SPLIT distance="150" swimtime="00:03:00.48" />
                    <SPLIT distance="200" swimtime="00:04:03.82" />
                    <SPLIT distance="250" swimtime="00:05:06.78" />
                    <SPLIT distance="300" swimtime="00:06:10.02" />
                    <SPLIT distance="350" swimtime="00:07:14.66" />
                    <SPLIT distance="400" swimtime="00:08:17.23" />
                    <SPLIT distance="450" swimtime="00:09:20.63" />
                    <SPLIT distance="500" swimtime="00:10:23.96" />
                    <SPLIT distance="550" swimtime="00:11:27.17" />
                    <SPLIT distance="600" swimtime="00:12:29.38" />
                    <SPLIT distance="650" swimtime="00:13:32.39" />
                    <SPLIT distance="700" swimtime="00:14:34.64" />
                    <SPLIT distance="750" swimtime="00:15:36.79" />
                    <SPLIT distance="800" swimtime="00:16:39.21" />
                    <SPLIT distance="850" swimtime="00:17:42.59" />
                    <SPLIT distance="900" swimtime="00:18:44.99" />
                    <SPLIT distance="950" swimtime="00:19:48.17" />
                    <SPLIT distance="1000" swimtime="00:20:51.41" />
                    <SPLIT distance="1050" swimtime="00:24:03.64" />
                    <SPLIT distance="1100" swimtime="00:22:59.69" />
                    <SPLIT distance="1200" swimtime="00:25:08.22" />
                    <SPLIT distance="1250" swimtime="00:28:22.03" />
                    <SPLIT distance="1300" swimtime="00:27:17.41" />
                    <SPLIT distance="1350" swimtime="00:30:29.87" />
                    <SPLIT distance="1400" swimtime="00:29:25.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="549" swimtime="00:00:52.25" resultid="5135" heatid="7996" lane="9" entrytime="00:00:50.00" />
                <RESULT eventid="1387" points="649" reactiontime="+106" swimtime="00:04:09.89" resultid="5136" heatid="8067" lane="3" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.16" />
                    <SPLIT distance="100" swimtime="00:02:01.60" />
                    <SPLIT distance="150" swimtime="00:03:06.90" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1554" points="773" swimtime="00:01:50.35" resultid="5137" heatid="8120" lane="9" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-11-02" firstname="Beata" gender="F" lastname="Sulewska" nation="POL" license="502611100009" athleteid="5138">
              <RESULTS>
                <RESULT eventid="1120" points="763" reactiontime="+81" swimtime="00:10:43.29" resultid="5139" heatid="8136" lane="3" entrytime="00:10:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                    <SPLIT distance="100" swimtime="00:01:14.03" />
                    <SPLIT distance="150" swimtime="00:01:53.49" />
                    <SPLIT distance="200" swimtime="00:02:33.35" />
                    <SPLIT distance="250" swimtime="00:03:13.38" />
                    <SPLIT distance="300" swimtime="00:03:53.97" />
                    <SPLIT distance="350" swimtime="00:04:34.32" />
                    <SPLIT distance="400" swimtime="00:05:15.79" />
                    <SPLIT distance="450" swimtime="00:05:56.83" />
                    <SPLIT distance="500" swimtime="00:06:38.29" />
                    <SPLIT distance="550" swimtime="00:07:19.31" />
                    <SPLIT distance="600" swimtime="00:08:00.84" />
                    <SPLIT distance="650" swimtime="00:08:41.78" />
                    <SPLIT distance="700" swimtime="00:09:23.39" />
                    <SPLIT distance="750" swimtime="00:10:03.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="655" reactiontime="+75" swimtime="00:01:10.08" resultid="5140" heatid="7978" lane="5" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1387" points="753" reactiontime="+81" swimtime="00:03:06.73" resultid="5141" heatid="8066" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.54" />
                    <SPLIT distance="100" swimtime="00:01:28.64" />
                    <SPLIT distance="150" swimtime="00:02:17.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1417" points="719" reactiontime="+85" swimtime="00:05:15.50" resultid="5142" heatid="8150" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.10" />
                    <SPLIT distance="100" swimtime="00:01:15.56" />
                    <SPLIT distance="150" swimtime="00:01:55.59" />
                    <SPLIT distance="200" swimtime="00:02:35.68" />
                    <SPLIT distance="250" swimtime="00:03:16.15" />
                    <SPLIT distance="300" swimtime="00:03:56.73" />
                    <SPLIT distance="350" swimtime="00:04:36.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="676" reactiontime="+81" swimtime="00:01:27.48" resultid="5143" heatid="8123" lane="6" entrytime="00:01:26.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-28" firstname="Wiesław" gender="M" lastname="Kornicki" nation="POL" license="502611200007" athleteid="5114">
              <RESULTS>
                <RESULT eventid="1105" points="611" reactiontime="+84" swimtime="00:00:35.97" resultid="5115" heatid="7964" lane="5" entrytime="00:00:36.00" />
                <RESULT eventid="1198" points="620" reactiontime="+89" swimtime="00:01:17.38" resultid="5116" heatid="7985" lane="1" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="733" reactiontime="+78" swimtime="00:00:31.93" resultid="5117" heatid="8055" lane="4" entrytime="00:00:32.00" />
                <RESULT eventid="1539" points="389" reactiontime="+73" swimtime="00:00:45.86" resultid="5118" heatid="8110" lane="3" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-11-29" firstname="Daniel" gender="M" lastname="Fecica" nation="POL" license="502611200002" athleteid="5124">
              <RESULTS>
                <RESULT eventid="1228" points="560" reactiontime="+75" swimtime="00:00:47.99" resultid="5125" heatid="8002" lane="8" entrytime="00:00:46.00" />
                <RESULT comment="Rekord Polski Masters" eventid="1402" points="818" reactiontime="+92" swimtime="00:03:38.14" resultid="5126" heatid="8073" lane="0" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.35" />
                    <SPLIT distance="100" swimtime="00:01:46.93" />
                    <SPLIT distance="150" swimtime="00:02:43.11" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski Masters" eventid="1569" points="708" reactiontime="+94" swimtime="00:01:40.85" resultid="5127" heatid="8126" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-10-05" firstname="Barbara" gender="F" lastname="Brendler" nation="POL" license="502611100005" athleteid="5145">
              <RESULTS>
                <RESULT eventid="1181" points="390" reactiontime="+100" swimtime="00:01:38.52" resultid="5146" heatid="7974" lane="3" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="281" reactiontime="+83" swimtime="00:04:58.96" resultid="5147" heatid="8019" lane="9" entrytime="00:04:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.98" />
                    <SPLIT distance="100" swimtime="00:02:28.08" />
                    <SPLIT distance="150" swimtime="00:03:44.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="497" reactiontime="+94" swimtime="00:00:41.03" resultid="5148" heatid="8045" lane="5" entrytime="00:00:40.00" />
                <RESULT eventid="1493" points="329" reactiontime="+92" swimtime="00:03:54.86" resultid="5149" heatid="8088" lane="9" entrytime="00:03:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.95" />
                    <SPLIT distance="100" swimtime="00:01:47.49" />
                    <SPLIT distance="150" swimtime="00:02:51.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-05-22" firstname="Włodzimierz" gender="M" lastname="Bosowski" nation="POL" license="502611200005" athleteid="5109">
              <RESULTS>
                <RESULT eventid="1105" points="226" reactiontime="+92" swimtime="00:00:50.08" resultid="5110" heatid="7963" lane="3" entrytime="00:00:42.00" />
                <RESULT eventid="1342" points="177" reactiontime="+110" swimtime="00:02:11.31" resultid="5111" heatid="8037" lane="3" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="312" reactiontime="+89" swimtime="00:00:42.42" resultid="5112" heatid="8053" lane="3" entrytime="00:00:38.00" />
                <RESULT eventid="1539" points="236" reactiontime="+96" swimtime="00:00:54.18" resultid="5113" heatid="8110" lane="8" entrytime="00:00:48.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SLOWRO" nation="POL" region="DOL" clubid="5156" name="WKS Śląsk Wrocław">
          <CONTACT email="murtacha68@gmail.com" name="Frank Marta" phone="604 231 250" />
          <ATHLETES>
            <ATHLETE birthdate="1970-03-11" firstname="Anna" gender="F" lastname="Głowiak" nation="POL" athleteid="5175">
              <RESULTS>
                <RESULT eventid="1181" points="526" reactiontime="+87" swimtime="00:01:17.67" resultid="5176" heatid="7977" lane="0" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="542" reactiontime="+91" swimtime="00:00:44.86" resultid="5177" heatid="7997" lane="0" entrytime="00:00:46.00" />
                <RESULT eventid="1357" points="612" reactiontime="+88" swimtime="00:00:33.38" resultid="5178" heatid="8047" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="1493" points="485" reactiontime="+88" swimtime="00:02:52.96" resultid="5179" heatid="8090" lane="2" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.78" />
                    <SPLIT distance="100" swimtime="00:01:19.69" />
                    <SPLIT distance="150" swimtime="00:02:05.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="520" reactiontime="+92" swimtime="00:01:39.63" resultid="5180" heatid="8120" lane="0" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-05-13" firstname="Maciej" gender="M" lastname="Dąbrowski" nation="POL" athleteid="5162">
              <RESULTS>
                <RESULT eventid="1075" points="590" reactiontime="+126" swimtime="00:02:53.81" resultid="5163" heatid="7949" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                    <SPLIT distance="100" swimtime="00:01:19.54" />
                    <SPLIT distance="150" swimtime="00:02:11.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="341" reactiontime="+111" swimtime="00:24:36.28" resultid="5164" heatid="8144" lane="8" entrytime="00:24:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.73" />
                    <SPLIT distance="100" swimtime="00:01:20.13" />
                    <SPLIT distance="150" swimtime="00:02:06.34" />
                    <SPLIT distance="200" swimtime="00:02:53.97" />
                    <SPLIT distance="250" swimtime="00:03:42.64" />
                    <SPLIT distance="300" swimtime="00:04:31.62" />
                    <SPLIT distance="350" swimtime="00:05:20.94" />
                    <SPLIT distance="400" swimtime="00:06:11.10" />
                    <SPLIT distance="450" swimtime="00:07:00.89" />
                    <SPLIT distance="500" swimtime="00:07:50.61" />
                    <SPLIT distance="550" swimtime="00:08:40.52" />
                    <SPLIT distance="600" swimtime="00:09:30.69" />
                    <SPLIT distance="650" swimtime="00:10:20.27" />
                    <SPLIT distance="700" swimtime="00:11:10.48" />
                    <SPLIT distance="750" swimtime="00:12:00.75" />
                    <SPLIT distance="800" swimtime="00:12:50.35" />
                    <SPLIT distance="850" swimtime="00:13:39.57" />
                    <SPLIT distance="900" swimtime="00:14:29.52" />
                    <SPLIT distance="950" swimtime="00:16:59.91" />
                    <SPLIT distance="1000" swimtime="00:16:09.87" />
                    <SPLIT distance="1050" swimtime="00:18:39.95" />
                    <SPLIT distance="1100" swimtime="00:17:49.53" />
                    <SPLIT distance="1200" swimtime="00:19:32.01" />
                    <SPLIT distance="1250" swimtime="00:20:24.12" />
                    <SPLIT distance="1300" swimtime="00:21:14.22" />
                    <SPLIT distance="1350" swimtime="00:22:05.50" />
                    <SPLIT distance="1400" swimtime="00:22:55.53" />
                    <SPLIT distance="1450" swimtime="00:23:46.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="5165" heatid="8025" lane="4" entrytime="00:02:55.00" />
                <RESULT eventid="1342" points="550" reactiontime="+76" swimtime="00:01:17.95" resultid="5166" heatid="8040" lane="6" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="397" reactiontime="+106" swimtime="00:01:22.69" resultid="5167" heatid="8084" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="552" reactiontime="+78" swimtime="00:00:35.63" resultid="5168" heatid="8113" lane="8" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-05-03" firstname="Marta" gender="F" lastname="Frank" nation="POL" athleteid="5169">
              <RESULTS>
                <RESULT eventid="1090" points="689" reactiontime="+70" swimtime="00:00:34.30" resultid="5170" heatid="7959" lane="2" entrytime="00:00:35.00" />
                <RESULT eventid="1273" points="724" reactiontime="+78" swimtime="00:02:57.22" resultid="5171" heatid="8020" lane="6" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.38" />
                    <SPLIT distance="100" swimtime="00:01:27.79" />
                    <SPLIT distance="150" swimtime="00:02:13.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="742" reactiontime="+74" swimtime="00:01:20.68" resultid="5172" heatid="8035" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="458" reactiontime="+86" swimtime="00:00:36.77" resultid="5173" heatid="8048" lane="0" entrytime="00:00:33.00" />
                <RESULT eventid="1524" points="787" reactiontime="+72" swimtime="00:00:35.93" resultid="5174" heatid="8106" lane="4" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-05-21" firstname="Marek" gender="M" lastname="Rother" nation="POL" athleteid="5157">
              <RESULTS>
                <RESULT eventid="1105" points="788" reactiontime="+83" swimtime="00:00:29.48" resultid="5158" heatid="7969" lane="7" entrytime="00:00:30.50" />
                <RESULT eventid="1288" points="952" reactiontime="+71" swimtime="00:02:23.96" resultid="5159" heatid="8028" lane="2" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                    <SPLIT distance="100" swimtime="00:01:10.14" />
                    <SPLIT distance="150" swimtime="00:01:47.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="926" reactiontime="+74" swimtime="00:01:05.54" resultid="5160" heatid="8043" lane="0" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="877" reactiontime="+66" swimtime="00:00:30.54" resultid="5161" heatid="8116" lane="5" entrytime="00:00:30.40" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1614" reactiontime="+65" swimtime="00:02:18.25" resultid="5181" heatid="8134" lane="1" entrytime="00:02:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.01" />
                    <SPLIT distance="100" swimtime="00:01:12.70" />
                    <SPLIT distance="150" swimtime="00:01:47.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5157" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="5175" number="2" />
                    <RELAYPOSITION athleteid="5169" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="5162" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="4689" name="Wodnik Siemianowice">
          <CONTACT email="bartolomeo863@wp.pl" name="Szymik" street="osiedle andaluzja 13/4/11" />
          <ATHLETES>
            <ATHLETE birthdate="1960-02-18" firstname="Piotr" gender="M" lastname="Szymik" nation="POL" athleteid="4690">
              <RESULTS>
                <RESULT eventid="1105" points="449" swimtime="00:00:37.24" resultid="4691" heatid="7964" lane="6" entrytime="00:00:36.50" />
                <RESULT eventid="1165" points="666" swimtime="00:22:35.50" resultid="4692" heatid="8144" lane="5" entrytime="00:22:15.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.61" />
                    <SPLIT distance="100" swimtime="00:01:22.81" />
                    <SPLIT distance="150" swimtime="00:02:08.20" />
                    <SPLIT distance="200" swimtime="00:02:54.13" />
                    <SPLIT distance="250" swimtime="00:03:39.96" />
                    <SPLIT distance="300" swimtime="00:04:25.70" />
                    <SPLIT distance="350" swimtime="00:05:11.13" />
                    <SPLIT distance="400" swimtime="00:05:56.30" />
                    <SPLIT distance="450" swimtime="00:06:42.50" />
                    <SPLIT distance="500" swimtime="00:07:28.04" />
                    <SPLIT distance="550" swimtime="00:08:12.98" />
                    <SPLIT distance="600" swimtime="00:08:58.72" />
                    <SPLIT distance="650" swimtime="00:09:44.34" />
                    <SPLIT distance="700" swimtime="00:10:29.75" />
                    <SPLIT distance="750" swimtime="00:11:14.71" />
                    <SPLIT distance="800" swimtime="00:11:59.24" />
                    <SPLIT distance="850" swimtime="00:12:45.50" />
                    <SPLIT distance="900" swimtime="00:13:30.46" />
                    <SPLIT distance="950" swimtime="00:14:15.84" />
                    <SPLIT distance="1000" swimtime="00:15:01.46" />
                    <SPLIT distance="1050" swimtime="00:15:47.85" />
                    <SPLIT distance="1100" swimtime="00:16:32.02" />
                    <SPLIT distance="1150" swimtime="00:17:17.75" />
                    <SPLIT distance="1200" swimtime="00:18:03.86" />
                    <SPLIT distance="1250" swimtime="00:18:50.19" />
                    <SPLIT distance="1300" swimtime="00:19:35.06" />
                    <SPLIT distance="1350" swimtime="00:20:20.92" />
                    <SPLIT distance="1400" swimtime="00:21:06.41" />
                    <SPLIT distance="1450" swimtime="00:21:51.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="456" reactiontime="+51" swimtime="00:03:21.50" resultid="4693" heatid="8015" lane="3" entrytime="00:03:20.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.60" />
                    <SPLIT distance="100" swimtime="00:01:38.33" />
                    <SPLIT distance="150" swimtime="00:02:29.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="569" reactiontime="+56" swimtime="00:05:56.02" resultid="4694" heatid="8153" lane="8" entrytime="00:05:37.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.41" />
                    <SPLIT distance="100" swimtime="00:01:22.87" />
                    <SPLIT distance="150" swimtime="00:02:09.07" />
                    <SPLIT distance="200" swimtime="00:02:55.08" />
                    <SPLIT distance="250" swimtime="00:03:41.57" />
                    <SPLIT distance="300" swimtime="00:04:27.12" />
                    <SPLIT distance="350" swimtime="00:05:13.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="385" reactiontime="+54" swimtime="00:01:28.82" resultid="4695" heatid="8083" lane="5" entrytime="00:01:25.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="561" reactiontime="+80" swimtime="00:06:43.20" resultid="4696" heatid="8164" lane="0" entrytime="00:06:39.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.98" />
                    <SPLIT distance="100" swimtime="00:01:39.36" />
                    <SPLIT distance="150" swimtime="00:02:30.89" />
                    <SPLIT distance="200" swimtime="00:03:22.74" />
                    <SPLIT distance="250" swimtime="00:04:19.16" />
                    <SPLIT distance="300" swimtime="00:05:16.82" />
                    <SPLIT distance="350" swimtime="00:06:00.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="POL" clubid="5230" name="WOPR Tczew">
          <CONTACT email="aleksandra.hebel@wp.pl" name="Aleksandra Hebel" />
          <ATHLETES>
            <ATHLETE birthdate="1987-06-22" firstname="Aleksandra" gender="F" lastname="Hebel" nation="POL" athleteid="5236">
              <RESULTS>
                <RESULT eventid="1181" points="465" reactiontime="+93" swimtime="00:01:15.83" resultid="5237" heatid="7977" lane="8" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="385" reactiontime="+99" swimtime="00:03:21.90" resultid="5238" heatid="8019" lane="6" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.06" />
                    <SPLIT distance="100" swimtime="00:01:37.89" />
                    <SPLIT distance="150" swimtime="00:02:30.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="400" reactiontime="+88" swimtime="00:01:32.00" resultid="5239" heatid="8034" lane="0" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="556" reactiontime="+89" swimtime="00:00:32.89" resultid="5240" heatid="8047" lane="7" entrytime="00:00:34.00" />
                <RESULT eventid="1493" points="399" reactiontime="+85" swimtime="00:02:55.11" resultid="5241" heatid="8089" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.27" />
                    <SPLIT distance="100" swimtime="00:01:22.28" />
                    <SPLIT distance="150" swimtime="00:02:09.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="373" reactiontime="+100" swimtime="00:00:43.19" resultid="5242" heatid="8105" lane="1" entrytime="00:00:44.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-09-12" firstname="Maciej" gender="M" lastname="Reschke" nation="POL" athleteid="5251">
              <RESULTS>
                <RESULT eventid="1105" points="486" reactiontime="+93" swimtime="00:00:31.87" resultid="5252" heatid="7965" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1198" points="599" reactiontime="+92" swimtime="00:01:01.32" resultid="5253" heatid="7988" lane="9" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="532" swimtime="00:00:36.16" resultid="5254" heatid="8007" lane="3" entrytime="00:00:36.00" />
                <RESULT eventid="1372" points="563" reactiontime="+78" swimtime="00:00:28.03" resultid="5255" heatid="8061" lane="4" entrytime="00:00:28.00" />
                <RESULT eventid="1432" points="528" reactiontime="+82" swimtime="00:05:10.33" resultid="5256" heatid="8151" lane="9" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                    <SPLIT distance="100" swimtime="00:01:09.29" />
                    <SPLIT distance="150" swimtime="00:01:47.85" />
                    <SPLIT distance="200" swimtime="00:02:27.20" />
                    <SPLIT distance="250" swimtime="00:03:07.77" />
                    <SPLIT distance="300" swimtime="00:03:49.30" />
                    <SPLIT distance="350" swimtime="00:04:30.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-02-18" firstname="Marek" gender="M" lastname="Stuczyński" nation="POL" athleteid="5257">
              <RESULTS>
                <RESULT eventid="1105" points="681" reactiontime="+77" swimtime="00:00:28.43" resultid="5258" heatid="7971" lane="8" entrytime="00:00:28.70" />
                <RESULT eventid="1228" points="811" reactiontime="+78" swimtime="00:00:31.29" resultid="5259" heatid="8010" lane="6" entrytime="00:00:31.50" />
                <RESULT eventid="1402" points="668" reactiontime="+80" swimtime="00:02:47.48" resultid="5260" heatid="8077" lane="8" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                    <SPLIT distance="100" swimtime="00:01:17.19" />
                    <SPLIT distance="150" swimtime="00:02:01.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="706" reactiontime="+76" swimtime="00:01:13.14" resultid="5261" heatid="8132" lane="1" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-10-28" firstname="Andrzej" gender="M" lastname="Gołembiewski" nation="POL" athleteid="5243">
              <RESULTS>
                <RESULT eventid="1135" points="522" reactiontime="+87" swimtime="00:10:47.03" resultid="5244" heatid="8139" lane="7" entrytime="00:11:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                    <SPLIT distance="100" swimtime="00:01:11.29" />
                    <SPLIT distance="150" swimtime="00:01:51.30" />
                    <SPLIT distance="200" swimtime="00:02:32.48" />
                    <SPLIT distance="250" swimtime="00:03:13.61" />
                    <SPLIT distance="300" swimtime="00:03:55.18" />
                    <SPLIT distance="350" swimtime="00:04:37.07" />
                    <SPLIT distance="400" swimtime="00:05:18.98" />
                    <SPLIT distance="450" swimtime="00:06:01.04" />
                    <SPLIT distance="500" swimtime="00:06:43.34" />
                    <SPLIT distance="550" swimtime="00:07:25.48" />
                    <SPLIT distance="600" swimtime="00:08:06.85" />
                    <SPLIT distance="650" swimtime="00:08:48.59" />
                    <SPLIT distance="700" swimtime="00:09:29.67" />
                    <SPLIT distance="750" swimtime="00:10:10.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="590" reactiontime="+82" swimtime="00:01:01.63" resultid="5245" heatid="7989" lane="2" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="660" reactiontime="+85" swimtime="00:00:33.65" resultid="5246" heatid="8008" lane="3" entrytime="00:00:34.00" />
                <RESULT eventid="1402" points="589" reactiontime="+83" swimtime="00:02:54.52" resultid="5247" heatid="8076" lane="6" entrytime="00:02:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.58" />
                    <SPLIT distance="100" swimtime="00:01:23.98" />
                    <SPLIT distance="150" swimtime="00:02:09.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="581" reactiontime="+85" swimtime="00:05:00.52" resultid="5248" heatid="8152" lane="4" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                    <SPLIT distance="100" swimtime="00:01:10.30" />
                    <SPLIT distance="150" swimtime="00:01:48.16" />
                    <SPLIT distance="200" swimtime="00:02:27.35" />
                    <SPLIT distance="250" swimtime="00:03:06.72" />
                    <SPLIT distance="300" swimtime="00:03:46.20" />
                    <SPLIT distance="350" swimtime="00:04:25.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="574" reactiontime="+86" swimtime="00:02:18.54" resultid="5249" heatid="8100" lane="1" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.27" />
                    <SPLIT distance="100" swimtime="00:01:06.21" />
                    <SPLIT distance="150" swimtime="00:01:42.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="556" reactiontime="+96" swimtime="00:01:18.62" resultid="5250" heatid="8132" lane="9" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WOPRWL" nation="POL" region="LBS" clubid="5185" name="WOPR Województwa Lubuskiego">
          <CONTACT city="Zielona Góra" email="kifertnat@gmail.com" name="Kifert" phone="606793089" state="LUBUS" street="Lisowskiego 1" zip="65-072" />
          <ATHLETES>
            <ATHLETE birthdate="1984-07-06" firstname="Małgorzata" gender="F" lastname="Fijałek-Żuk" nation="POL" athleteid="5204">
              <RESULTS>
                <RESULT eventid="1058" points="580" reactiontime="+81" swimtime="00:02:55.77" resultid="5205" heatid="7944" lane="4" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="100" swimtime="00:01:18.97" />
                    <SPLIT distance="150" swimtime="00:02:11.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1387" points="545" reactiontime="+75" swimtime="00:03:16.30" resultid="5206" heatid="8070" lane="9" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.05" />
                    <SPLIT distance="100" swimtime="00:01:32.66" />
                    <SPLIT distance="150" swimtime="00:02:24.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-02-20" firstname="Kalina" gender="F" lastname="Chęcińska" nation="POL" athleteid="5195">
              <RESULTS>
                <RESULT eventid="1090" points="449" reactiontime="+89" swimtime="00:00:38.78" resultid="5196" heatid="7957" lane="7" entrytime="00:00:38.80" />
                <RESULT eventid="1181" points="515" reactiontime="+86" swimtime="00:01:14.48" resultid="5197" heatid="7976" lane="4" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="560" reactiontime="+83" swimtime="00:00:33.30" resultid="5198" heatid="8047" lane="3" entrytime="00:00:34.00" />
                <RESULT eventid="1447" points="348" reactiontime="+87" swimtime="00:01:34.67" resultid="5199" heatid="8078" lane="5" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-07-16" firstname="Mariusz" gender="M" lastname="Kachel" nation="POL" athleteid="5218">
              <RESULTS>
                <RESULT eventid="1105" points="680" reactiontime="+82" swimtime="00:00:29.44" resultid="5219" heatid="7970" lane="2" entrytime="00:00:29.00" />
                <RESULT eventid="1228" points="608" reactiontime="+81" swimtime="00:00:36.00" resultid="5220" heatid="8008" lane="9" entrytime="00:00:35.00" />
                <RESULT eventid="1569" points="589" reactiontime="+87" swimtime="00:01:21.97" resultid="5221" heatid="8130" lane="4" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-03-23" firstname="Lilianna" gender="F" lastname="Wilk" nation="POL" athleteid="5207">
              <RESULTS>
                <RESULT eventid="1090" points="663" reactiontime="+79" swimtime="00:00:32.45" resultid="5208" heatid="7960" lane="1" entrytime="00:00:33.00" />
                <RESULT eventid="1181" points="598" reactiontime="+73" swimtime="00:01:09.72" resultid="5209" heatid="7978" lane="3" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="594" reactiontime="+75" swimtime="00:02:54.69" resultid="5210" heatid="8021" lane="0" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                    <SPLIT distance="100" swimtime="00:01:23.84" />
                    <SPLIT distance="150" swimtime="00:02:09.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="619" reactiontime="+82" swimtime="00:00:31.74" resultid="5211" heatid="8049" lane="1" entrytime="00:00:31.50" />
                <RESULT eventid="1447" points="609" reactiontime="+69" swimtime="00:01:15.67" resultid="5212" heatid="8080" lane="8" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="524" reactiontime="+78" swimtime="00:02:39.91" resultid="5213" heatid="8091" lane="7" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                    <SPLIT distance="100" swimtime="00:01:16.40" />
                    <SPLIT distance="150" swimtime="00:01:58.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-06-10" firstname="Łukasz" gender="M" lastname="Osik" nation="POL" athleteid="5214">
              <RESULTS>
                <RESULT eventid="1105" points="491" reactiontime="+91" swimtime="00:00:32.33" resultid="5215" heatid="7970" lane="3" entrytime="00:00:29.00" />
                <RESULT eventid="1198" points="557" reactiontime="+92" swimtime="00:01:03.16" resultid="5216" heatid="7990" lane="0" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="554" reactiontime="+89" swimtime="00:00:28.64" resultid="5217" heatid="8061" lane="9" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-07-02" firstname="Natalia" gender="F" lastname="Kifert" nation="POL" athleteid="5191">
              <RESULTS>
                <RESULT eventid="1273" points="432" reactiontime="+79" swimtime="00:03:09.70" resultid="5192" heatid="8020" lane="7" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.49" />
                    <SPLIT distance="100" swimtime="00:01:34.70" />
                    <SPLIT distance="150" swimtime="00:02:23.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="545" reactiontime="+73" swimtime="00:01:24.65" resultid="5193" heatid="8034" lane="3" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1524" points="568" reactiontime="+67" swimtime="00:00:38.51" resultid="5194" heatid="8106" lane="2" entrytime="00:00:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-02-20" firstname="Mateusz" gender="M" lastname="Chęciński" nation="POL" athleteid="5200">
              <RESULTS>
                <RESULT eventid="1288" points="793" reactiontime="+75" swimtime="00:02:24.22" resultid="5201" heatid="8028" lane="6" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                    <SPLIT distance="100" swimtime="00:01:08.82" />
                    <SPLIT distance="150" swimtime="00:01:45.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="769" reactiontime="+76" swimtime="00:01:07.71" resultid="5202" heatid="8043" lane="2" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="766" reactiontime="+74" swimtime="00:00:30.81" resultid="5203" heatid="8116" lane="4" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-04-11" firstname="Radomir" gender="M" lastname="Kifert" nation="POL" athleteid="5186">
              <RESULTS>
                <RESULT eventid="1105" points="680" reactiontime="+87" swimtime="00:00:29.44" resultid="5187" heatid="7968" lane="9" entrytime="00:00:32.00" />
                <RESULT eventid="1228" points="596" swimtime="00:00:36.24" resultid="5188" heatid="8007" lane="6" entrytime="00:00:36.00" />
                <RESULT eventid="1342" points="682" reactiontime="+74" swimtime="00:01:11.51" resultid="5189" heatid="8042" lane="6" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1539" points="688" reactiontime="+67" swimtime="00:00:32.27" resultid="5190" heatid="8115" lane="5" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-04-23" firstname="Wojciech" gender="M" lastname="Pabiński" nation="POL" athleteid="5222">
              <RESULTS>
                <RESULT eventid="1105" points="376" reactiontime="+84" swimtime="00:00:34.64" resultid="5223" heatid="7970" lane="5" entrytime="00:00:29.00" />
                <RESULT eventid="1228" points="408" reactiontime="+79" swimtime="00:00:39.33" resultid="5224" heatid="8006" lane="2" entrytime="00:00:37.00" />
                <RESULT eventid="1372" points="527" reactiontime="+67" swimtime="00:00:28.78" resultid="5225" heatid="8063" lane="8" entrytime="00:00:27.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1318" reactiontime="+84" swimtime="00:04:16.79" resultid="5227" heatid="8030" lane="4" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                    <SPLIT distance="100" swimtime="00:01:04.46" />
                    <SPLIT distance="150" swimtime="00:01:36.30" />
                    <SPLIT distance="200" swimtime="00:02:09.36" />
                    <SPLIT distance="250" swimtime="00:02:38.54" />
                    <SPLIT distance="300" swimtime="00:03:12.01" />
                    <SPLIT distance="350" swimtime="00:03:42.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5214" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="5218" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="5186" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="5200" number="4" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1303" reactiontime="+80" swimtime="00:05:00.47" resultid="5228" heatid="8029" lane="2" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                    <SPLIT distance="100" swimtime="00:01:13.99" />
                    <SPLIT distance="150" swimtime="00:01:48.26" />
                    <SPLIT distance="200" swimtime="00:02:28.68" />
                    <SPLIT distance="250" swimtime="00:03:06.90" />
                    <SPLIT distance="300" swimtime="00:03:48.23" />
                    <SPLIT distance="350" swimtime="00:04:21.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5204" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="5195" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="5191" number="3" reactiontime="+70" />
                    <RELAYPOSITION athleteid="5207" number="4" reactiontime="+67" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1614" reactiontime="+78" swimtime="00:02:11.54" resultid="5229" heatid="8135" lane="1" entrytime="00:02:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.51" />
                    <SPLIT distance="100" swimtime="00:01:06.23" />
                    <SPLIT distance="150" swimtime="00:01:38.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5186" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="5204" number="2" />
                    <RELAYPOSITION athleteid="5207" number="3" reactiontime="+69" />
                    <RELAYPOSITION athleteid="5200" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1614" reactiontime="+67" swimtime="00:02:19.11" resultid="5226" heatid="8134" lane="5" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.07" />
                    <SPLIT distance="100" swimtime="00:01:14.29" />
                    <SPLIT distance="150" swimtime="00:01:46.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5191" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="5218" number="2" />
                    <RELAYPOSITION athleteid="5214" number="3" reactiontime="+61" />
                    <RELAYPOSITION athleteid="5195" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WAGRO" nation="POL" region="WIE" clubid="3473" name="Wągrowiec">
          <CONTACT city="WĄGROWIEC" email="obywatel-ag@xl.wp.pl" name="GUZIAŁ ANDRZEJ" phone="508030407" state="WIELK" street="OSIEDLE NIEPODLEGŁOŚCI 9/4" zip="62-100" />
          <ATHLETES>
            <ATHLETE birthdate="1954-09-30" firstname="Andrzej" gender="M" lastname="Guział" nation="POL" athleteid="3483">
              <RESULTS>
                <RESULT eventid="1198" points="462" reactiontime="+85" swimtime="00:01:18.91" resultid="3484" heatid="7984" lane="8" entrytime="00:01:18.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="445" reactiontime="+93" swimtime="00:00:44.99" resultid="3485" heatid="8003" lane="8" entrytime="00:00:42.36" />
                <RESULT eventid="1372" points="526" reactiontime="+104" swimtime="00:00:33.84" resultid="3486" heatid="8054" lane="4" entrytime="00:00:34.41" />
                <RESULT eventid="1569" points="496" reactiontime="+98" swimtime="00:01:40.20" resultid="3487" heatid="8127" lane="7" entrytime="00:01:36.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ZKS DRZONK" nation="POL" region="LBS" clubid="5345" name="ZKS Drzonków">
          <CONTACT city="ZIELONA GÓRA /ŁĘŻYCA" email="llfpiotr@gmail.com" name="BARTA PIOTR" phone="602347348" state="LUBUS" street="ODRZAŃSKA 21" zip="66-016" />
          <ATHLETES>
            <ATHLETE birthdate="1971-03-18" firstname="Piotr" gender="M" lastname="Barta" nation="POL" athleteid="5346">
              <RESULTS>
                <RESULT eventid="1228" points="736" reactiontime="+87" swimtime="00:00:33.78" resultid="5347" heatid="8008" lane="2" entrytime="00:00:34.21" entrycourse="LCM" />
                <RESULT comment="Rekord Polski Masters" eventid="1402" points="834" reactiontime="+85" swimtime="00:02:40.21" resultid="5348" heatid="8077" lane="1" entrytime="00:02:42.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.49" />
                    <SPLIT distance="100" swimtime="00:01:15.77" />
                    <SPLIT distance="150" swimtime="00:01:57.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="830" reactiontime="+84" swimtime="00:01:13.13" resultid="5350" heatid="8132" lane="0" entrytime="00:01:13.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="647" reactiontime="+91" swimtime="00:05:27.19" resultid="5351" heatid="8162" lane="1" entrytime="00:05:39.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                    <SPLIT distance="100" swimtime="00:01:12.54" />
                    <SPLIT distance="150" swimtime="00:02:00.46" />
                    <SPLIT distance="200" swimtime="00:02:46.30" />
                    <SPLIT distance="250" swimtime="00:03:30.22" />
                    <SPLIT distance="300" swimtime="00:04:15.45" />
                    <SPLIT distance="350" swimtime="00:04:52.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="714" reactiontime="+86" swimtime="00:04:44.55" resultid="8291" heatid="8156" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.96" />
                    <SPLIT distance="100" swimtime="00:01:09.93" />
                    <SPLIT distance="150" swimtime="00:01:45.88" />
                    <SPLIT distance="200" swimtime="00:02:22.08" />
                    <SPLIT distance="250" swimtime="00:02:58.01" />
                    <SPLIT distance="300" swimtime="00:03:33.70" />
                    <SPLIT distance="350" swimtime="00:04:09.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" nation="RUS" clubid="5352" name="Zvezdy Rossii">
          <CONTACT email="a.tervinsky@gov39.ru" name="Tervinsky" />
          <ATHLETES>
            <ATHLETE birthdate="1963-01-01" firstname="Sergei" gender="M" lastname="Dirindyaev" nation="RUS" athleteid="5433">
              <RESULTS>
                <RESULT eventid="1135" points="377" reactiontime="+100" swimtime="00:12:59.99" resultid="5434" heatid="8140" lane="4" entrytime="00:11:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.61" />
                    <SPLIT distance="100" swimtime="00:01:27.52" />
                    <SPLIT distance="150" swimtime="00:02:15.56" />
                    <SPLIT distance="200" swimtime="00:03:05.11" />
                    <SPLIT distance="250" swimtime="00:03:54.83" />
                    <SPLIT distance="300" swimtime="00:04:45.24" />
                    <SPLIT distance="350" swimtime="00:05:35.34" />
                    <SPLIT distance="400" swimtime="00:06:25.37" />
                    <SPLIT distance="450" swimtime="00:07:14.65" />
                    <SPLIT distance="500" swimtime="00:08:04.91" />
                    <SPLIT distance="550" swimtime="00:08:54.42" />
                    <SPLIT distance="600" swimtime="00:09:44.28" />
                    <SPLIT distance="650" swimtime="00:10:33.18" />
                    <SPLIT distance="700" swimtime="00:11:23.03" />
                    <SPLIT distance="750" swimtime="00:12:12.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="5435" heatid="7987" lane="3" entrytime="00:01:06.00" />
                <RESULT eventid="1372" status="DNS" swimtime="00:00:00.00" resultid="5436" heatid="8057" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1509" status="DNS" swimtime="00:00:00.00" resultid="5438" heatid="8098" lane="2" entrytime="00:02:38.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Irina" gender="F" lastname="Shangina" nation="RUS" athleteid="5358">
              <RESULTS>
                <RESULT eventid="1058" points="804" reactiontime="+83" swimtime="00:03:11.50" resultid="5359" heatid="7943" lane="8" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                    <SPLIT distance="100" swimtime="00:01:31.36" />
                    <SPLIT distance="150" swimtime="00:02:24.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="738" swimtime="00:00:42.57" resultid="5360" heatid="7998" lane="9" entrytime="00:00:42.00" />
                <RESULT eventid="1387" points="993" reactiontime="+89" swimtime="00:03:16.51" resultid="5361" heatid="8070" lane="0" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.25" />
                    <SPLIT distance="100" swimtime="00:01:34.88" />
                    <SPLIT distance="150" swimtime="00:02:26.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="977" reactiontime="+86" swimtime="00:01:30.55" resultid="5362" heatid="8122" lane="0" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Elena" gender="F" lastname="Kolyadina" nation="RUS" athleteid="5363">
              <RESULTS>
                <RESULT eventid="1090" points="538" reactiontime="+88" swimtime="00:00:43.09" resultid="5364" heatid="7956" lane="2" entrytime="00:00:45.00" />
                <RESULT eventid="1181" points="692" reactiontime="+81" swimtime="00:01:19.44" resultid="5365" heatid="7976" lane="9" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="705" reactiontime="+90" swimtime="00:00:43.22" resultid="5366" heatid="7997" lane="2" entrytime="00:00:43.00" />
                <RESULT eventid="1357" points="775" reactiontime="+80" swimtime="00:00:34.34" resultid="5367" heatid="8046" lane="4" entrytime="00:00:35.50" />
                <RESULT eventid="1387" points="761" reactiontime="+88" swimtime="00:03:34.75" resultid="5368" heatid="8069" lane="0" entrytime="00:03:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.74" />
                    <SPLIT distance="100" swimtime="00:01:42.66" />
                    <SPLIT distance="150" swimtime="00:02:38.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="762" reactiontime="+87" swimtime="00:01:38.35" resultid="5369" heatid="8121" lane="2" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-01-01" firstname="Svetlana" gender="F" lastname="Kozlova" nation="RUS" athleteid="5387">
              <RESULTS>
                <RESULT eventid="1058" points="781" reactiontime="+86" swimtime="00:02:56.20" resultid="5388" heatid="7943" lane="3" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.32" />
                    <SPLIT distance="100" swimtime="00:01:25.25" />
                    <SPLIT distance="150" swimtime="00:02:14.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="701" swimtime="00:00:42.48" resultid="5389" heatid="7998" lane="1" entrytime="00:00:41.50" />
                <RESULT eventid="1387" points="819" reactiontime="+92" swimtime="00:03:15.80" resultid="5390" heatid="8070" lane="6" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.67" />
                    <SPLIT distance="100" swimtime="00:01:36.64" />
                    <SPLIT distance="150" swimtime="00:02:26.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="792" reactiontime="+83" swimtime="00:01:30.21" resultid="5391" heatid="8123" lane="8" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1584" points="763" reactiontime="+90" swimtime="00:06:27.22" resultid="5392" heatid="8159" lane="9" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.36" />
                    <SPLIT distance="100" swimtime="00:01:30.34" />
                    <SPLIT distance="150" swimtime="00:02:21.75" />
                    <SPLIT distance="200" swimtime="00:03:11.93" />
                    <SPLIT distance="250" swimtime="00:04:03.96" />
                    <SPLIT distance="300" swimtime="00:04:55.39" />
                    <SPLIT distance="350" swimtime="00:05:42.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Aleksandr" gender="M" lastname="Smirnov" nation="RUS" athleteid="5452">
              <RESULTS>
                <RESULT eventid="1165" points="662" reactiontime="+86" swimtime="00:19:43.23" resultid="5453" heatid="8143" lane="2" entrytime="00:20:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.76" />
                    <SPLIT distance="100" swimtime="00:01:13.38" />
                    <SPLIT distance="150" swimtime="00:01:52.87" />
                    <SPLIT distance="200" swimtime="00:02:32.72" />
                    <SPLIT distance="250" swimtime="00:03:12.02" />
                    <SPLIT distance="300" swimtime="00:03:52.18" />
                    <SPLIT distance="350" swimtime="00:04:31.95" />
                    <SPLIT distance="400" swimtime="00:05:11.94" />
                    <SPLIT distance="450" swimtime="00:05:51.47" />
                    <SPLIT distance="500" swimtime="00:06:31.36" />
                    <SPLIT distance="550" swimtime="00:07:11.07" />
                    <SPLIT distance="600" swimtime="00:07:50.99" />
                    <SPLIT distance="650" swimtime="00:08:30.50" />
                    <SPLIT distance="700" swimtime="00:09:10.41" />
                    <SPLIT distance="750" swimtime="00:09:50.10" />
                    <SPLIT distance="800" swimtime="00:10:30.31" />
                    <SPLIT distance="850" swimtime="00:11:10.26" />
                    <SPLIT distance="900" swimtime="00:11:50.19" />
                    <SPLIT distance="950" swimtime="00:12:29.47" />
                    <SPLIT distance="1000" swimtime="00:13:09.48" />
                    <SPLIT distance="1050" swimtime="00:13:48.94" />
                    <SPLIT distance="1100" swimtime="00:14:29.28" />
                    <SPLIT distance="1150" swimtime="00:15:08.89" />
                    <SPLIT distance="1200" swimtime="00:15:49.08" />
                    <SPLIT distance="1250" swimtime="00:16:28.62" />
                    <SPLIT distance="1300" swimtime="00:17:08.79" />
                    <SPLIT distance="1350" swimtime="00:17:48.28" />
                    <SPLIT distance="1400" swimtime="00:18:28.12" />
                    <SPLIT distance="1450" swimtime="00:19:07.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="635" reactiontime="+79" swimtime="00:02:18.87" resultid="5455" heatid="8101" lane="8" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                    <SPLIT distance="100" swimtime="00:01:07.39" />
                    <SPLIT distance="150" swimtime="00:01:43.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1432" points="653" swimtime="00:04:55.20" resultid="8326" heatid="8325" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                    <SPLIT distance="100" swimtime="00:01:10.44" />
                    <SPLIT distance="150" swimtime="00:01:48.35" />
                    <SPLIT distance="200" swimtime="00:02:26.91" />
                    <SPLIT distance="250" swimtime="00:03:05.06" />
                    <SPLIT distance="300" swimtime="00:03:42.99" />
                    <SPLIT distance="350" swimtime="00:04:20.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-01" firstname="Olga" gender="F" lastname="Veryukina" nation="RUS" athleteid="5398">
              <RESULTS>
                <RESULT eventid="1090" points="661" reactiontime="+89" swimtime="00:00:34.19" resultid="5399" heatid="7960" lane="0" entrytime="00:00:34.00" />
                <RESULT eventid="1120" points="663" reactiontime="+89" swimtime="00:11:14.10" resultid="5400" heatid="8136" lane="2" entrytime="00:11:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.42" />
                    <SPLIT distance="100" swimtime="00:01:18.03" />
                    <SPLIT distance="150" swimtime="00:01:59.74" />
                    <SPLIT distance="200" swimtime="00:02:42.15" />
                    <SPLIT distance="250" swimtime="00:03:24.49" />
                    <SPLIT distance="300" swimtime="00:04:07.40" />
                    <SPLIT distance="350" swimtime="00:04:50.46" />
                    <SPLIT distance="400" swimtime="00:05:33.41" />
                    <SPLIT distance="450" swimtime="00:06:16.37" />
                    <SPLIT distance="500" swimtime="00:06:59.65" />
                    <SPLIT distance="550" swimtime="00:07:42.62" />
                    <SPLIT distance="600" swimtime="00:08:25.60" />
                    <SPLIT distance="650" swimtime="00:09:08.31" />
                    <SPLIT distance="700" swimtime="00:09:50.88" />
                    <SPLIT distance="750" swimtime="00:10:32.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="652" reactiontime="+84" swimtime="00:01:10.18" resultid="5401" heatid="7978" lane="1" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="621" reactiontime="+82" swimtime="00:00:32.29" resultid="5402" heatid="8049" lane="9" entrytime="00:00:32.00" />
                <RESULT eventid="1417" points="651" reactiontime="+93" swimtime="00:05:26.16" resultid="5403" heatid="8147" lane="7" entrytime="00:05:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="100" swimtime="00:01:17.73" />
                    <SPLIT distance="150" swimtime="00:01:59.34" />
                    <SPLIT distance="200" swimtime="00:02:41.66" />
                    <SPLIT distance="250" swimtime="00:03:23.65" />
                    <SPLIT distance="300" swimtime="00:04:05.66" />
                    <SPLIT distance="350" swimtime="00:04:46.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="660" reactiontime="+88" swimtime="00:02:33.09" resultid="5404" heatid="8091" lane="4" entrytime="00:02:33.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                    <SPLIT distance="100" swimtime="00:01:12.85" />
                    <SPLIT distance="150" swimtime="00:01:52.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Viktor" gender="M" lastname="Lyubavin" nation="RUS" athleteid="5439">
              <RESULTS>
                <RESULT eventid="1135" points="483" reactiontime="+85" swimtime="00:11:15.49" resultid="5440" heatid="8139" lane="1" entrytime="00:11:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.13" />
                    <SPLIT distance="100" swimtime="00:01:15.17" />
                    <SPLIT distance="150" swimtime="00:01:56.97" />
                    <SPLIT distance="200" swimtime="00:02:39.92" />
                    <SPLIT distance="250" swimtime="00:03:22.88" />
                    <SPLIT distance="300" swimtime="00:04:04.92" />
                    <SPLIT distance="350" swimtime="00:04:47.33" />
                    <SPLIT distance="400" swimtime="00:05:30.65" />
                    <SPLIT distance="450" swimtime="00:06:14.56" />
                    <SPLIT distance="500" swimtime="00:06:57.98" />
                    <SPLIT distance="550" swimtime="00:07:41.47" />
                    <SPLIT distance="600" swimtime="00:08:25.44" />
                    <SPLIT distance="650" swimtime="00:09:08.39" />
                    <SPLIT distance="700" swimtime="00:09:51.78" />
                    <SPLIT distance="750" swimtime="00:10:34.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="641" reactiontime="+83" swimtime="00:01:04.76" resultid="5441" heatid="7990" lane="8" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="489" swimtime="00:00:37.95" resultid="5442" heatid="8007" lane="7" entrytime="00:00:36.50" />
                <RESULT eventid="1372" points="666" reactiontime="+79" swimtime="00:00:28.81" resultid="5443" heatid="8060" lane="1" entrytime="00:00:28.50" />
                <RESULT eventid="1402" points="541" reactiontime="+86" swimtime="00:03:08.57" resultid="5444" heatid="8075" lane="2" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.81" />
                    <SPLIT distance="100" swimtime="00:01:31.33" />
                    <SPLIT distance="150" swimtime="00:02:20.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="537" reactiontime="+81" swimtime="00:02:26.82" resultid="5445" heatid="8100" lane="6" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                    <SPLIT distance="100" swimtime="00:01:10.75" />
                    <SPLIT distance="150" swimtime="00:01:49.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1569" points="546" reactiontime="+83" swimtime="00:01:24.30" resultid="5446" heatid="8130" lane="1" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-01" firstname="Vladimir" gender="M" lastname="Chekutov" nation="RUS" athleteid="5447">
              <RESULTS>
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="5448" heatid="7989" lane="7" entrytime="00:01:04.00" />
                <RESULT eventid="1342" status="DNS" swimtime="00:00:00.00" resultid="5449" heatid="8041" lane="3" entrytime="00:01:14.00" />
                <RESULT eventid="1372" status="DNS" swimtime="00:00:00.00" resultid="5450" heatid="8060" lane="7" entrytime="00:00:28.50" />
                <RESULT eventid="1539" status="DNS" swimtime="00:00:00.00" resultid="5451" heatid="8114" lane="5" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Sergei" gender="M" lastname="Mikhaylov" nation="RUS" athleteid="5422">
              <RESULTS>
                <RESULT eventid="1165" points="461" reactiontime="+99" swimtime="00:25:31.50" resultid="5423" heatid="8145" lane="3" entrytime="00:27:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.21" />
                    <SPLIT distance="100" swimtime="00:01:34.78" />
                    <SPLIT distance="150" swimtime="00:02:24.84" />
                    <SPLIT distance="200" swimtime="00:03:15.23" />
                    <SPLIT distance="250" swimtime="00:04:05.89" />
                    <SPLIT distance="300" swimtime="00:04:57.17" />
                    <SPLIT distance="350" swimtime="00:05:48.03" />
                    <SPLIT distance="400" swimtime="00:06:39.42" />
                    <SPLIT distance="450" swimtime="00:07:30.32" />
                    <SPLIT distance="500" swimtime="00:08:21.56" />
                    <SPLIT distance="550" swimtime="00:09:13.08" />
                    <SPLIT distance="600" swimtime="00:10:04.11" />
                    <SPLIT distance="650" swimtime="00:10:55.63" />
                    <SPLIT distance="700" swimtime="00:11:47.48" />
                    <SPLIT distance="750" swimtime="00:12:38.96" />
                    <SPLIT distance="800" swimtime="00:13:29.66" />
                    <SPLIT distance="850" swimtime="00:14:20.74" />
                    <SPLIT distance="900" swimtime="00:15:12.19" />
                    <SPLIT distance="950" swimtime="00:16:03.57" />
                    <SPLIT distance="1000" swimtime="00:16:56.01" />
                    <SPLIT distance="1050" swimtime="00:17:47.87" />
                    <SPLIT distance="1100" swimtime="00:18:39.78" />
                    <SPLIT distance="1150" swimtime="00:19:30.84" />
                    <SPLIT distance="1200" swimtime="00:20:23.01" />
                    <SPLIT distance="1250" swimtime="00:21:15.02" />
                    <SPLIT distance="1300" swimtime="00:22:06.68" />
                    <SPLIT distance="1350" swimtime="00:22:58.16" />
                    <SPLIT distance="1400" swimtime="00:23:50.90" />
                    <SPLIT distance="1450" swimtime="00:24:41.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="317" reactiontime="+94" swimtime="00:01:29.10" resultid="5424" heatid="7982" lane="5" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1372" points="305" reactiontime="+94" swimtime="00:00:39.52" resultid="5425" heatid="8053" lane="1" entrytime="00:00:39.50" />
                <RESULT eventid="1432" points="445" reactiontime="+96" swimtime="00:06:26.44" resultid="5426" heatid="8155" lane="3" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.58" />
                    <SPLIT distance="100" swimtime="00:01:30.34" />
                    <SPLIT distance="150" swimtime="00:02:20.12" />
                    <SPLIT distance="200" swimtime="00:03:09.72" />
                    <SPLIT distance="250" swimtime="00:03:59.66" />
                    <SPLIT distance="300" swimtime="00:04:48.90" />
                    <SPLIT distance="350" swimtime="00:05:38.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1509" points="382" reactiontime="+92" swimtime="00:03:07.58" resultid="5427" heatid="8095" lane="7" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.61" />
                    <SPLIT distance="100" swimtime="00:01:29.34" />
                    <SPLIT distance="150" swimtime="00:02:18.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-20" firstname="Sergey" gender="M" lastname="Petrov" nation="RUS" athleteid="2212">
              <RESULTS>
                <RESULT eventid="1105" points="703" reactiontime="+71" swimtime="00:00:29.12" resultid="2213" heatid="7971" lane="9" entrytime="00:00:29.00" entrycourse="LCM" />
                <RESULT eventid="1228" points="785" reactiontime="+71" swimtime="00:00:33.07" resultid="2214" heatid="8009" lane="3" entrytime="00:00:33.00" entrycourse="LCM" />
                <RESULT eventid="1372" points="700" reactiontime="+73" swimtime="00:00:27.68" resultid="2215" heatid="8061" lane="1" entrytime="00:00:28.00" entrycourse="LCM" />
                <RESULT eventid="1569" points="722" reactiontime="+72" swimtime="00:01:16.58" resultid="2216" heatid="8131" lane="5" entrytime="00:01:15.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1938-01-01" firstname="Luiza" gender="F" lastname="Shcherbich" nation="RUS" athleteid="5353">
              <RESULTS>
                <RESULT eventid="1181" points="208" reactiontime="+137" swimtime="00:02:34.68" resultid="5354" heatid="7973" lane="2" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="274" reactiontime="+127" swimtime="00:01:13.21" resultid="5355" heatid="7994" lane="4" entrytime="00:01:09.00" />
                <RESULT eventid="1357" points="235" reactiontime="+129" swimtime="00:01:04.48" resultid="5356" heatid="8044" lane="5" entrytime="00:00:59.00" />
                <RESULT eventid="1554" points="285" reactiontime="+125" swimtime="00:02:53.61" resultid="5357" heatid="8119" lane="9" entrytime="00:02:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-01-01" firstname="Irina" gender="F" lastname="Titova" nation="RUS" athleteid="5377">
              <RESULTS>
                <RESULT eventid="1181" points="570" reactiontime="+97" swimtime="00:01:17.42" resultid="5378" heatid="7976" lane="2" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="526" reactiontime="+95" swimtime="00:00:35.18" resultid="5379" heatid="8046" lane="5" entrytime="00:00:35.50" />
                <RESULT eventid="1493" points="545" reactiontime="+99" swimtime="00:02:48.96" resultid="5380" heatid="8090" lane="6" entrytime="00:02:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                    <SPLIT distance="100" swimtime="00:01:21.35" />
                    <SPLIT distance="150" swimtime="00:02:05.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Natalia" gender="F" lastname="Aleshchenko" nation="RUS" athleteid="5370">
              <RESULTS>
                <RESULT eventid="1058" points="786" reactiontime="+92" swimtime="00:03:08.17" resultid="5371" heatid="7943" lane="1" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.95" />
                    <SPLIT distance="100" swimtime="00:01:29.46" />
                    <SPLIT distance="150" swimtime="00:02:23.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="832" reactiontime="+94" swimtime="00:00:36.82" resultid="5372" heatid="7957" lane="3" entrytime="00:00:38.00" />
                <RESULT eventid="1181" points="728" reactiontime="+81" swimtime="00:01:16.85" resultid="5373" heatid="7976" lane="5" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="732" reactiontime="+82" swimtime="00:00:34.26" resultid="5374" heatid="8047" lane="1" entrytime="00:00:34.50" />
                <RESULT eventid="1447" points="789" reactiontime="+91" swimtime="00:01:25.78" resultid="5375" heatid="8079" lane="7" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1493" points="753" reactiontime="+87" swimtime="00:02:52.34" resultid="5376" heatid="8090" lane="5" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.40" />
                    <SPLIT distance="100" swimtime="00:01:23.27" />
                    <SPLIT distance="150" swimtime="00:02:09.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-01" firstname="Elena" gender="F" lastname="Dautova" nation="RUS" athleteid="5393">
              <RESULTS>
                <RESULT eventid="1273" points="466" reactiontime="+69" swimtime="00:03:18.53" resultid="5394" heatid="8019" lane="5" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.12" />
                    <SPLIT distance="100" swimtime="00:01:35.72" />
                    <SPLIT distance="150" swimtime="00:02:27.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="538" reactiontime="+77" swimtime="00:01:26.16" resultid="5395" heatid="8034" lane="1" entrytime="00:01:25.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="639" reactiontime="+87" swimtime="00:00:31.98" resultid="5396" heatid="8048" lane="1" entrytime="00:00:32.50" />
                <RESULT eventid="1524" points="610" reactiontime="+65" swimtime="00:00:38.53" resultid="5397" heatid="8106" lane="7" entrytime="00:00:39.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-01" firstname="Elena" gender="F" lastname="Mekhteleva" nation="RUS" athleteid="5405">
              <RESULTS>
                <RESULT eventid="1090" status="DNS" swimtime="00:00:00.00" resultid="5406" heatid="7959" lane="1" entrytime="00:00:35.00" />
                <RESULT eventid="1213" points="767" reactiontime="+97" swimtime="00:00:36.75" resultid="5407" heatid="7999" lane="3" entrytime="00:00:37.00" />
                <RESULT eventid="1387" points="689" reactiontime="+91" swimtime="00:03:09.27" resultid="5408" heatid="8070" lane="5" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.28" />
                    <SPLIT distance="100" swimtime="00:01:29.75" />
                    <SPLIT distance="150" swimtime="00:02:19.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1554" points="783" reactiontime="+89" swimtime="00:01:21.75" resultid="5409" heatid="8123" lane="5" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-01" firstname="Grigorii" gender="M" lastname="Lopin" nation="RUS" athleteid="5428">
              <RESULTS>
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="5429" heatid="7949" lane="8" entrytime="00:03:10.00" />
                <RESULT eventid="1228" points="514" reactiontime="+90" swimtime="00:00:40.16" resultid="5430" heatid="8005" lane="1" entrytime="00:00:39.50" />
                <RESULT eventid="1402" points="468" reactiontime="+89" swimtime="00:03:26.10" resultid="5431" heatid="8074" lane="0" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.57" />
                    <SPLIT distance="100" swimtime="00:01:44.19" />
                    <SPLIT distance="150" swimtime="00:02:36.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1599" points="488" reactiontime="+92" swimtime="00:06:44.73" resultid="5432" heatid="8165" lane="5" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.95" />
                    <SPLIT distance="100" swimtime="00:01:39.09" />
                    <SPLIT distance="150" swimtime="00:02:34.40" />
                    <SPLIT distance="200" swimtime="00:03:28.62" />
                    <SPLIT distance="250" swimtime="00:04:22.08" />
                    <SPLIT distance="300" swimtime="00:05:17.00" />
                    <SPLIT distance="350" swimtime="00:06:03.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-01-01" firstname="Regina" gender="F" lastname="Sych" nation="RUS" athleteid="5410">
              <RESULTS>
                <RESULT eventid="1090" points="880" reactiontime="+90" swimtime="00:00:29.53" resultid="5411" heatid="7960" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="1181" points="943" reactiontime="+81" swimtime="00:00:59.89" resultid="5412" heatid="7979" lane="7" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="972" reactiontime="+79" swimtime="00:00:27.30" resultid="5413" heatid="8050" lane="3" entrytime="00:00:28.50" />
                <RESULT eventid="1493" status="DNS" swimtime="00:00:00.00" resultid="5414" heatid="8092" lane="6" entrytime="00:02:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-01-01" firstname="Aleksandr" gender="M" lastname="Tervinskii" nation="RUS" athleteid="5415">
              <RESULTS>
                <RESULT eventid="1105" points="267" reactiontime="+90" swimtime="00:00:44.28" resultid="5416" heatid="7963" lane="6" entrytime="00:00:42.50" />
                <RESULT eventid="1228" points="424" reactiontime="+91" swimtime="00:00:41.32" resultid="5417" heatid="8003" lane="0" entrytime="00:00:42.50" />
                <RESULT eventid="1342" status="DNS" swimtime="00:00:00.00" resultid="5418" heatid="8038" lane="8" entrytime="00:01:40.50" />
                <RESULT eventid="1372" points="491" reactiontime="+88" swimtime="00:00:33.72" resultid="5419" heatid="8054" lane="5" entrytime="00:00:34.50" />
                <RESULT eventid="1539" status="DNS" swimtime="00:00:00.00" resultid="5420" heatid="8111" lane="1" entrytime="00:00:43.00" />
                <RESULT eventid="1569" points="392" reactiontime="+90" swimtime="00:01:39.48" resultid="5421" heatid="8126" lane="5" entrytime="00:01:40.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1318" reactiontime="+75" swimtime="00:04:22.42" resultid="5463" heatid="8030" lane="2" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                    <SPLIT distance="100" swimtime="00:01:04.02" />
                    <SPLIT distance="150" swimtime="00:01:33.13" />
                    <SPLIT distance="200" swimtime="00:02:06.57" />
                    <SPLIT distance="250" swimtime="00:02:37.39" />
                    <SPLIT distance="300" swimtime="00:03:10.37" />
                    <SPLIT distance="350" swimtime="00:03:43.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5452" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="5447" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="5439" number="3" reactiontime="+17" />
                    <RELAYPOSITION athleteid="5415" number="4" reactiontime="+76" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT comment="S4 - Przedwczesna zmiana sztafetowa" eventid="1303" reactiontime="+93" status="DSQ" swimtime="00:05:24.84" resultid="5461" heatid="8029" lane="1" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.79" />
                    <SPLIT distance="100" swimtime="00:01:24.00" />
                    <SPLIT distance="150" swimtime="00:01:56.91" />
                    <SPLIT distance="200" swimtime="00:02:38.71" />
                    <SPLIT distance="250" swimtime="00:03:17.12" />
                    <SPLIT distance="300" swimtime="00:04:05.02" />
                    <SPLIT distance="350" swimtime="00:04:42.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5370" number="1" reactiontime="+93" status="DSQ" />
                    <RELAYPOSITION athleteid="5410" number="2" reactiontime="-40" status="DSQ" />
                    <RELAYPOSITION athleteid="5358" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="5377" number="4" reactiontime="+70" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1303" reactiontime="+82" swimtime="00:04:47.33" resultid="5462" heatid="8029" lane="8" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                    <SPLIT distance="100" swimtime="00:01:11.60" />
                    <SPLIT distance="150" swimtime="00:01:44.78" />
                    <SPLIT distance="200" swimtime="00:02:21.79" />
                    <SPLIT distance="250" swimtime="00:02:56.45" />
                    <SPLIT distance="300" swimtime="00:03:33.62" />
                    <SPLIT distance="350" swimtime="00:04:08.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5393" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="5405" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="5398" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="5387" number="4" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="1614" reactiontime="+76" swimtime="00:03:27.84" resultid="5464" heatid="8133" lane="2" entrytime="00:03:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.64" />
                    <SPLIT distance="100" swimtime="00:01:41.57" />
                    <SPLIT distance="150" swimtime="00:02:22.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5415" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="5363" number="2" />
                    <RELAYPOSITION athleteid="5428" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="5353" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="X" number="5">
              <RESULTS>
                <RESULT eventid="1614" reactiontime="+78" swimtime="00:02:24.53" resultid="5465" heatid="8134" lane="0" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.81" />
                    <SPLIT distance="100" swimtime="00:01:18.39" />
                    <SPLIT distance="150" swimtime="00:01:52.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5452" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="5358" number="2" />
                    <RELAYPOSITION athleteid="5398" number="3" reactiontime="+64" />
                    <RELAYPOSITION athleteid="5433" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="6">
              <RESULTS>
                <RESULT eventid="1614" reactiontime="+73" swimtime="00:02:11.79" resultid="5466" heatid="8135" lane="9" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                    <SPLIT distance="100" swimtime="00:01:14.64" />
                    <SPLIT distance="150" swimtime="00:01:44.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5447" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="5405" number="2" />
                    <RELAYPOSITION athleteid="5410" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="5439" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>

<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Wielkopolski Okregowy Zwiazek Plywacki" version="Build 17589">
    <CONTACT name="GeoLogix AG" street="Muristrasse 60" city="Bern" zip="3006" country="CH" phone="+41 31 356 80 56" fax="+41 31 356 80 81" email="info@splash-software.ch" internet="http://www.splash-software.ch" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Poznań" name="Zimowe Otwarte Mistrzostwa Polski w Pływaniu w Kategorii Masters Poznań 2011" course="SCM" nation="POL" timing="AUTOMATIC">
      <AGEDATE value="2011-01-01" type="YEAR" />
      <POOL lanemax="8" />
      <POINTTABLE pointtableid="1013" name="DSV Performance Table" version="2009" />
      <SESSIONS>
        <SESSION date="2011-11-18" daytime="16:30" number="1">
          <EVENTS>
            <EVENT eventid="1058" daytime="16:30" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1060" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3657" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1061" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4629" />
                    <RANKING order="2" place="2" resultid="3223" />
                    <RANKING order="3" place="3" resultid="1964" />
                    <RANKING order="4" place="4" resultid="4262" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1062" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4829" />
                    <RANKING order="2" place="2" resultid="2759" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1063" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3984" />
                    <RANKING order="2" place="-1" resultid="1853" />
                    <RANKING order="3" place="-1" resultid="5193" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1064" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="1065" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2470" />
                    <RANKING order="2" place="2" resultid="5037" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4514" />
                    <RANKING order="2" place="2" resultid="1916" />
                    <RANKING order="3" place="3" resultid="1931" />
                    <RANKING order="4" place="4" resultid="1951" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3736" />
                    <RANKING order="2" place="2" resultid="2391" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1068" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2673" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1070" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4841" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4865" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1072" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1073" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1074" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1059" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6713" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6714" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6715" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1075" daytime="17:25" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1076" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4914" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1077" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4855" />
                    <RANKING order="2" place="2" resultid="4597" />
                    <RANKING order="3" place="3" resultid="2424" />
                    <RANKING order="4" place="4" resultid="4495" />
                    <RANKING order="5" place="-1" resultid="2767" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1078" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3019" />
                    <RANKING order="2" place="2" resultid="4377" />
                    <RANKING order="3" place="3" resultid="5058" />
                    <RANKING order="4" place="4" resultid="3487" />
                    <RANKING order="5" place="-1" resultid="5073" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1079" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3347" />
                    <RANKING order="2" place="2" resultid="3328" />
                    <RANKING order="3" place="3" resultid="4554" />
                    <RANKING order="4" place="4" resultid="3479" />
                    <RANKING order="5" place="5" resultid="4667" />
                    <RANKING order="6" place="6" resultid="2049" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1080" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2616" />
                    <RANKING order="2" place="2" resultid="4040" />
                    <RANKING order="3" place="3" resultid="3291" />
                    <RANKING order="4" place="4" resultid="3502" />
                    <RANKING order="5" place="5" resultid="3111" />
                    <RANKING order="6" place="6" resultid="4033" />
                    <RANKING order="7" place="7" resultid="4013" />
                    <RANKING order="8" place="8" resultid="2577" />
                    <RANKING order="9" place="9" resultid="4720" />
                    <RANKING order="10" place="10" resultid="4139" />
                    <RANKING order="11" place="-1" resultid="2293" />
                    <RANKING order="12" place="-1" resultid="2233" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1081" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3700" />
                    <RANKING order="2" place="2" resultid="3308" />
                    <RANKING order="3" place="3" resultid="5029" />
                    <RANKING order="4" place="-1" resultid="2594" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1082" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5245" />
                    <RANKING order="2" place="2" resultid="3465" />
                    <RANKING order="3" place="3" resultid="5356" />
                    <RANKING order="4" place="4" resultid="2599" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1083" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4065" />
                    <RANKING order="2" place="2" resultid="2351" />
                    <RANKING order="3" place="3" resultid="5378" />
                    <RANKING order="4" place="4" resultid="3364" />
                    <RANKING order="5" place="5" resultid="3342" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1084" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4004" />
                    <RANKING order="2" place="2" resultid="2359" />
                    <RANKING order="3" place="3" resultid="5249" />
                    <RANKING order="4" place="4" resultid="3449" />
                    <RANKING order="5" place="5" resultid="4698" />
                    <RANKING order="6" place="6" resultid="4427" />
                    <RANKING order="7" place="7" resultid="6712" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1085" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2644" />
                    <RANKING order="2" place="-1" resultid="3989" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1086" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2529" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1087" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4107" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1088" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="2321" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1089" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4197" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1090" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1091" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6716" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6717" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6718" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6719" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6720" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6721" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6722" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1092" daytime="19:10" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1093" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2053" />
                    <RANKING order="2" place="2" resultid="2522" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2956" />
                    <RANKING order="2" place="2" resultid="2916" />
                    <RANKING order="3" place="3" resultid="3804" />
                    <RANKING order="4" place="4" resultid="2921" />
                    <RANKING order="5" place="5" resultid="2723" />
                    <RANKING order="6" place="6" resultid="2961" />
                    <RANKING order="7" place="7" resultid="2119" />
                    <RANKING order="8" place="8" resultid="4388" />
                    <RANKING order="9" place="9" resultid="4395" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1095" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2753" />
                    <RANKING order="2" place="2" resultid="3665" />
                    <RANKING order="3" place="3" resultid="3970" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1096" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2835" />
                    <RANKING order="2" place="2" resultid="2623" />
                    <RANKING order="3" place="3" resultid="5187" />
                    <RANKING order="4" place="4" resultid="5371" />
                    <RANKING order="5" place="5" resultid="2780" />
                    <RANKING order="6" place="6" resultid="1945" />
                    <RANKING order="7" place="-1" resultid="2132" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1097" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4588" />
                    <RANKING order="2" place="2" resultid="2343" />
                    <RANKING order="3" place="3" resultid="3569" />
                    <RANKING order="4" place="4" resultid="3495" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2106" />
                    <RANKING order="2" place="2" resultid="2156" />
                    <RANKING order="3" place="3" resultid="2611" />
                    <RANKING order="4" place="4" resultid="3077" />
                    <RANKING order="5" place="5" resultid="5180" />
                    <RANKING order="6" place="6" resultid="2731" />
                    <RANKING order="7" place="7" resultid="4170" />
                    <RANKING order="8" place="8" resultid="4163" />
                    <RANKING order="9" place="9" resultid="4276" />
                    <RANKING order="10" place="10" resultid="3170" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1099" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5173" />
                    <RANKING order="2" place="2" resultid="2148" />
                    <RANKING order="3" place="3" resultid="1972" />
                    <RANKING order="4" place="4" resultid="2124" />
                    <RANKING order="5" place="5" resultid="3578" />
                    <RANKING order="6" place="-1" resultid="4676" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1100" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4177" />
                    <RANKING order="2" place="2" resultid="2014" />
                    <RANKING order="3" place="3" resultid="4099" />
                    <RANKING order="4" place="4" resultid="3964" />
                    <RANKING order="5" place="5" resultid="5161" />
                    <RANKING order="6" place="6" resultid="1991" />
                    <RANKING order="7" place="7" resultid="4636" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1101" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2853" />
                    <RANKING order="2" place="2" resultid="5155" />
                    <RANKING order="3" place="3" resultid="2655" />
                    <RANKING order="4" place="4" resultid="2114" />
                    <RANKING order="5" place="5" resultid="3162" />
                    <RANKING order="6" place="-1" resultid="2817" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2874" />
                    <RANKING order="2" place="2" resultid="1985" />
                    <RANKING order="3" place="3" resultid="4955" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1103" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1104" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1105" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1106" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1107" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1108" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6723" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6724" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6725" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6726" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6727" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6728" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6729" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1109" daytime="19:26" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1110" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3838" />
                    <RANKING order="2" place="2" resultid="3777" />
                    <RANKING order="3" place="3" resultid="1893" />
                    <RANKING order="4" place="4" resultid="3773" />
                    <RANKING order="5" place="5" resultid="3785" />
                    <RANKING order="6" place="6" resultid="2066" />
                    <RANKING order="7" place="7" resultid="3814" />
                    <RANKING order="8" place="8" resultid="2074" />
                    <RANKING order="9" place="9" resultid="1861" />
                    <RANKING order="10" place="10" resultid="5095" />
                    <RANKING order="11" place="11" resultid="4908" />
                    <RANKING order="12" place="12" resultid="2090" />
                    <RANKING order="13" place="-1" resultid="2082" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1111" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4412" />
                    <RANKING order="2" place="2" resultid="2903" />
                    <RANKING order="3" place="3" resultid="3872" />
                    <RANKING order="4" place="4" resultid="2932" />
                    <RANKING order="5" place="5" resultid="2950" />
                    <RANKING order="6" place="6" resultid="5050" />
                    <RANKING order="7" place="7" resultid="4211" />
                    <RANKING order="8" place="8" resultid="2739" />
                    <RANKING order="9" place="9" resultid="2910" />
                    <RANKING order="10" place="10" resultid="2667" />
                    <RANKING order="11" place="11" resultid="2939" />
                    <RANKING order="12" place="12" resultid="3867" />
                    <RANKING order="13" place="13" resultid="3205" />
                    <RANKING order="14" place="14" resultid="4128" />
                    <RANKING order="15" place="15" resultid="4756" />
                    <RANKING order="16" place="-1" resultid="2945" />
                    <RANKING order="17" place="-1" resultid="5124" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1112" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3301" />
                    <RANKING order="2" place="2" resultid="5143" />
                    <RANKING order="3" place="3" resultid="3846" />
                    <RANKING order="4" place="4" resultid="3649" />
                    <RANKING order="5" place="5" resultid="4562" />
                    <RANKING order="6" place="6" resultid="4346" />
                    <RANKING order="7" place="7" resultid="5103" />
                    <RANKING order="8" place="8" resultid="4330" />
                    <RANKING order="9" place="9" resultid="3672" />
                    <RANKING order="10" place="10" resultid="4318" />
                    <RANKING order="11" place="11" resultid="5065" />
                    <RANKING order="12" place="12" resultid="2745" />
                    <RANKING order="13" place="13" resultid="4340" />
                    <RANKING order="14" place="14" resultid="3441" />
                    <RANKING order="15" place="15" resultid="3641" />
                    <RANKING order="16" place="16" resultid="4325" />
                    <RANKING order="17" place="17" resultid="4361" />
                    <RANKING order="18" place="18" resultid="2537" />
                    <RANKING order="19" place="19" resultid="4071" />
                    <RANKING order="20" place="-1" resultid="4794" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1113" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3425" />
                    <RANKING order="2" place="2" resultid="3510" />
                    <RANKING order="3" place="3" resultid="3417" />
                    <RANKING order="4" place="4" resultid="3070" />
                    <RANKING order="5" place="5" resultid="4370" />
                    <RANKING order="6" place="6" resultid="2222" />
                    <RANKING order="7" place="7" resultid="3371" />
                    <RANKING order="8" place="8" resultid="2238" />
                    <RANKING order="9" place="9" resultid="3433" />
                    <RANKING order="10" place="10" resultid="3849" />
                    <RANKING order="11" place="-1" resultid="2679" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1114" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2511" />
                    <RANKING order="2" place="2" resultid="5363" />
                    <RANKING order="3" place="3" resultid="4547" />
                    <RANKING order="4" place="4" resultid="5333" />
                    <RANKING order="5" place="5" resultid="3457" />
                    <RANKING order="6" place="6" resultid="2187" />
                    <RANKING order="7" place="7" resultid="3859" />
                    <RANKING order="8" place="8" resultid="5261" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1115" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2561" />
                    <RANKING order="2" place="2" resultid="3591" />
                    <RANKING order="3" place="3" resultid="3085" />
                    <RANKING order="4" place="4" resultid="3261" />
                    <RANKING order="5" place="5" resultid="5045" />
                    <RANKING order="6" place="6" resultid="2193" />
                    <RANKING order="7" place="7" resultid="1888" />
                    <RANKING order="8" place="8" resultid="4658" />
                    <RANKING order="9" place="9" resultid="4712" />
                    <RANKING order="10" place="10" resultid="2214" />
                    <RANKING order="11" place="11" resultid="4218" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1116" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2706" />
                    <RANKING order="2" place="2" resultid="2556" />
                    <RANKING order="3" place="3" resultid="3035" />
                    <RANKING order="4" place="4" resultid="2477" />
                    <RANKING order="5" place="5" resultid="4823" />
                    <RANKING order="6" place="6" resultid="4203" />
                    <RANKING order="7" place="7" resultid="3910" />
                    <RANKING order="8" place="8" resultid="4529" />
                    <RANKING order="9" place="9" resultid="4225" />
                    <RANKING order="10" place="10" resultid="3894" />
                    <RANKING order="11" place="11" resultid="4244" />
                    <RANKING order="12" place="12" resultid="3393" />
                    <RANKING order="13" place="13" resultid="3730" />
                    <RANKING order="14" place="-1" resultid="3473" />
                    <RANKING order="15" place="-1" resultid="2483" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1117" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3059" />
                    <RANKING order="2" place="2" resultid="4616" />
                    <RANKING order="3" place="3" resultid="4936" />
                    <RANKING order="4" place="4" resultid="2336" />
                    <RANKING order="5" place="5" resultid="4684" />
                    <RANKING order="6" place="6" resultid="3629" />
                    <RANKING order="7" place="7" resultid="3385" />
                    <RANKING order="8" place="8" resultid="4185" />
                    <RANKING order="9" place="9" resultid="4881" />
                    <RANKING order="10" place="10" resultid="3624" />
                    <RANKING order="11" place="11" resultid="3004" />
                    <RANKING order="12" place="12" resultid="4526" />
                    <RANKING order="13" place="13" resultid="3679" />
                    <RANKING order="14" place="14" resultid="3752" />
                    <RANKING order="15" place="15" resultid="2775" />
                    <RANKING order="16" place="-1" resultid="4897" />
                    <RANKING order="17" place="-1" resultid="4520" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1118" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4291" />
                    <RANKING order="2" place="2" resultid="2888" />
                    <RANKING order="3" place="3" resultid="5226" />
                    <RANKING order="4" place="4" resultid="2713" />
                    <RANKING order="5" place="5" resultid="4503" />
                    <RANKING order="6" place="6" resultid="2375" />
                    <RANKING order="7" place="7" resultid="3830" />
                    <RANKING order="8" place="8" resultid="3376" />
                    <RANKING order="9" place="9" resultid="2582" />
                    <RANKING order="10" place="10" resultid="3141" />
                    <RANKING order="11" place="-1" resultid="3950" />
                    <RANKING order="12" place="-1" resultid="3611" />
                    <RANKING order="13" place="-1" resultid="2859" />
                    <RANKING order="14" place="-1" resultid="5427" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1119" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4056" />
                    <RANKING order="2" place="2" resultid="5220" />
                    <RANKING order="3" place="3" resultid="5348" />
                    <RANKING order="4" place="4" resultid="5208" />
                    <RANKING order="5" place="-1" resultid="2866" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1120" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1923" />
                    <RANKING order="2" place="2" resultid="2497" />
                    <RANKING order="3" place="3" resultid="4690" />
                    <RANKING order="4" place="4" resultid="2367" />
                    <RANKING order="5" place="-1" resultid="4115" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1121" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1122" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4609" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1123" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1124" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1125" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6730" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6731" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6732" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6733" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6734" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6735" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6736" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6737" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6738" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6739" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6740" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="6741" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="6742" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="6743" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="6744" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="6745" number="16" order="16" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1126" daytime="19:57" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1127" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2416" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1128" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3117" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1129" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2569" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1130" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2164" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1131" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3822" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1132" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3319" />
                    <RANKING order="2" place="2" resultid="3274" />
                    <RANKING order="3" place="3" resultid="3723" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1133" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3012" />
                    <RANKING order="2" place="2" resultid="5168" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1134" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4270" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1135" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3211" />
                    <RANKING order="2" place="-1" resultid="4948" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1136" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2846" />
                    <RANKING order="2" place="-1" resultid="4623" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1137" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1138" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1139" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1140" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1141" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1142" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6746" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6747" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1143" daytime="21:05" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1144" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1903" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1145" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2328" />
                    <RANKING order="2" place="-1" resultid="3556" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1146" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4310" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1147" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2201" />
                    <RANKING order="2" place="2" resultid="3237" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1148" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3518" />
                    <RANKING order="2" place="2" resultid="3027" />
                    <RANKING order="3" place="3" resultid="2699" />
                    <RANKING order="4" place="-1" resultid="2210" />
                    <RANKING order="5" place="-1" resultid="4049" />
                    <RANKING order="6" place="-1" resultid="3228" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1149" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4847" />
                    <RANKING order="2" place="2" resultid="4541" />
                    <RANKING order="3" place="3" resultid="5026" />
                    <RANKING order="4" place="4" resultid="2517" />
                    <RANKING order="5" place="5" resultid="4136" />
                    <RANKING order="6" place="6" resultid="3337" />
                    <RANKING order="7" place="-1" resultid="3934" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1150" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3708" />
                    <RANKING order="2" place="2" resultid="4026" />
                    <RANKING order="3" place="3" resultid="3563" />
                    <RANKING order="4" place="4" resultid="3095" />
                    <RANKING order="5" place="5" resultid="2997" />
                    <RANKING order="6" place="6" resultid="4944" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1151" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2006" />
                    <RANKING order="2" place="2" resultid="2808" />
                    <RANKING order="3" place="3" resultid="2824" />
                    <RANKING order="4" place="4" resultid="3401" />
                    <RANKING order="5" place="5" resultid="4777" />
                    <RANKING order="6" place="6" resultid="2399" />
                    <RANKING order="7" place="7" resultid="4769" />
                    <RANKING order="8" place="-1" resultid="3149" />
                    <RANKING order="9" place="-1" resultid="3760" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1152" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2463" />
                    <RANKING order="2" place="2" resultid="3717" />
                    <RANKING order="3" place="3" resultid="2407" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1153" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1154" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3998" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1155" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="4154" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1156" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1157" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1158" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1159" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6748" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6749" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6750" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6751" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6752" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1160" daytime="23:22" gender="F" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1161" agemax="96" agemin="80" />
                <AGEGROUP agegroupid="1162" agemax="119" agemin="100">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2972" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1163" agemax="159" agemin="120">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2790" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1164" agemax="199" agemin="160">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2257" />
                    <RANKING order="2" place="-1" resultid="5289" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1165" agemax="239" agemin="200">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2244" />
                    <RANKING order="2" place="2" resultid="5294" />
                    <RANKING order="3" place="3" resultid="4981" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1166" agemax="279" agemin="240">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3186" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1167" agemax="319" agemin="280" />
                <AGEGROUP agegroupid="1168" agemax="359" agemin="320" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6813" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1177" daytime="23:27" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1178" agemax="96" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3793" />
                    <RANKING order="2" place="2" resultid="2095" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1179" agemax="119" agemin="100">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2973" />
                    <RANKING order="2" place="2" resultid="3877" />
                    <RANKING order="3" place="-1" resultid="1905" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1180" agemax="159" agemin="120">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6658" />
                    <RANKING order="2" place="2" resultid="1906" />
                    <RANKING order="3" place="3" resultid="3525" />
                    <RANKING order="4" place="4" resultid="2791" />
                    <RANKING order="5" place="5" resultid="3684" />
                    <RANKING order="6" place="6" resultid="4403" />
                    <RANKING order="7" place="7" resultid="4401" />
                    <RANKING order="8" place="8" resultid="4402" />
                    <RANKING order="9" place="9" resultid="6659" />
                    <RANKING order="10" place="-1" resultid="2247" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1181" agemax="199" agemin="160">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2246" />
                    <RANKING order="2" place="2" resultid="3526" />
                    <RANKING order="3" place="3" resultid="6668" />
                    <RANKING order="4" place="-1" resultid="3313" />
                    <RANKING order="5" place="-1" resultid="3043" />
                    <RANKING order="6" place="-1" resultid="4251" />
                    <RANKING order="7" place="-1" resultid="4567" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1182" agemax="239" agemin="200">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4569" />
                    <RANKING order="2" place="2" resultid="3527" />
                    <RANKING order="3" place="3" resultid="4982" />
                    <RANKING order="4" place="4" resultid="2248" />
                    <RANKING order="5" place="-1" resultid="5293" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1183" agemax="279" agemin="240">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2380" />
                    <RANKING order="2" place="2" resultid="5291" />
                    <RANKING order="3" place="-1" resultid="3188" />
                    <RANKING order="4" place="-1" resultid="4743" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1184" agemax="319" agemin="280" />
                <AGEGROUP agegroupid="1185" agemax="359" agemin="320" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6807" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6808" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6809" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6810" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2011-11-19" daytime="09:30" number="2">
          <EVENTS>
            <EVENT eventid="1187" daytime="09:30" gender="F" number="9" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1189" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3332" />
                    <RANKING order="2" place="2" resultid="2054" />
                    <RANKING order="3" place="3" resultid="3978" />
                    <RANKING order="4" place="4" resultid="3269" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1190" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1876" />
                    <RANKING order="2" place="2" resultid="2922" />
                    <RANKING order="3" place="3" resultid="4630" />
                    <RANKING order="4" place="4" resultid="3118" />
                    <RANKING order="5" place="5" resultid="2660" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1191" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3053" />
                    <RANKING order="2" place="2" resultid="4808" />
                    <RANKING order="3" place="3" resultid="3255" />
                    <RANKING order="4" place="4" resultid="4384" />
                    <RANKING order="5" place="5" resultid="2639" />
                    <RANKING order="6" place="6" resultid="4830" />
                    <RANKING order="7" place="7" resultid="3251" />
                    <RANKING order="8" place="-1" resultid="2760" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1192" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2836" />
                    <RANKING order="2" place="2" resultid="5372" />
                    <RANKING order="3" place="3" resultid="2686" />
                    <RANKING order="4" place="4" resultid="2781" />
                    <RANKING order="5" place="5" resultid="5183" />
                    <RANKING order="6" place="6" resultid="2133" />
                    <RANKING order="7" place="7" resultid="5283" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1193" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4589" />
                    <RANKING order="2" place="-1" resultid="4728" />
                    <RANKING order="3" place="-1" resultid="4650" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1194" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2107" />
                    <RANKING order="2" place="2" resultid="2157" />
                    <RANKING order="3" place="3" resultid="3078" />
                    <RANKING order="4" place="4" resultid="4171" />
                    <RANKING order="5" place="-1" resultid="3171" />
                    <RANKING order="6" place="-1" resultid="4931" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1195" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3013" />
                    <RANKING order="2" place="2" resultid="2149" />
                    <RANKING order="3" place="3" resultid="4677" />
                    <RANKING order="4" place="4" resultid="1973" />
                    <RANKING order="5" place="5" resultid="3409" />
                    <RANKING order="6" place="6" resultid="3065" />
                    <RANKING order="7" place="7" resultid="5169" />
                    <RANKING order="8" place="8" resultid="2490" />
                    <RANKING order="9" place="9" resultid="1939" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1196" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4178" />
                    <RANKING order="2" place="2" resultid="4100" />
                    <RANKING order="3" place="3" resultid="4271" />
                    <RANKING order="4" place="4" resultid="2392" />
                    <RANKING order="5" place="-1" resultid="2015" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1197" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3956" />
                    <RANKING order="2" place="2" resultid="5156" />
                    <RANKING order="3" place="3" resultid="2818" />
                    <RANKING order="4" place="4" resultid="2656" />
                    <RANKING order="5" place="5" resultid="2674" />
                    <RANKING order="6" place="6" resultid="3212" />
                    <RANKING order="7" place="7" resultid="3163" />
                    <RANKING order="8" place="-1" resultid="4949" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1198" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2875" />
                    <RANKING order="2" place="2" resultid="2026" />
                    <RANKING order="3" place="3" resultid="2450" />
                    <RANKING order="4" place="4" resultid="4956" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1199" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4092" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1200" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1201" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3103" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1202" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3157" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1203" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1204" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6821" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6822" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6823" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6824" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6825" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6826" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6827" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6828" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1205" daytime="09:47" gender="M" number="10" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1206" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3839" />
                    <RANKING order="2" place="2" resultid="2439" />
                    <RANKING order="3" place="3" resultid="3778" />
                    <RANKING order="4" place="4" resultid="4233" />
                    <RANKING order="5" place="5" resultid="1862" />
                    <RANKING order="6" place="6" resultid="5096" />
                    <RANKING order="7" place="7" resultid="2075" />
                    <RANKING order="8" place="8" resultid="3810" />
                    <RANKING order="9" place="9" resultid="2067" />
                    <RANKING order="10" place="10" resultid="1868" />
                    <RANKING order="11" place="11" resultid="3905" />
                    <RANKING order="12" place="-1" resultid="5018" />
                    <RANKING order="13" place="-1" resultid="2083" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1207" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3769" />
                    <RANKING order="2" place="2" resultid="4856" />
                    <RANKING order="3" place="3" resultid="2933" />
                    <RANKING order="4" place="4" resultid="1882" />
                    <RANKING order="5" place="5" resultid="4598" />
                    <RANKING order="6" place="6" resultid="2927" />
                    <RANKING order="7" place="7" resultid="5135" />
                    <RANKING order="8" place="8" resultid="3868" />
                    <RANKING order="9" place="9" resultid="3206" />
                    <RANKING order="10" place="10" resultid="4129" />
                    <RANKING order="11" place="11" resultid="4757" />
                    <RANKING order="12" place="12" resultid="4491" />
                    <RANKING order="13" place="-1" resultid="2735" />
                    <RANKING order="14" place="-1" resultid="5111" />
                    <RANKING order="15" place="-1" resultid="4046" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1208" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2589" />
                    <RANKING order="2" place="2" resultid="3637" />
                    <RANKING order="3" place="3" resultid="3650" />
                    <RANKING order="4" place="4" resultid="3020" />
                    <RANKING order="5" place="5" resultid="5144" />
                    <RANKING order="6" place="6" resultid="4563" />
                    <RANKING order="7" place="7" resultid="4331" />
                    <RANKING order="8" place="8" resultid="2746" />
                    <RANKING order="9" place="9" resultid="4352" />
                    <RANKING order="10" place="10" resultid="3642" />
                    <RANKING order="11" place="11" resultid="3442" />
                    <RANKING order="12" place="12" resultid="2719" />
                    <RANKING order="13" place="13" resultid="4357" />
                    <RANKING order="14" place="14" resultid="2538" />
                    <RANKING order="15" place="15" resultid="4336" />
                    <RANKING order="16" place="16" resultid="3745" />
                    <RANKING order="17" place="17" resultid="4319" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1209" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3426" />
                    <RANKING order="2" place="2" resultid="3418" />
                    <RANKING order="3" place="3" resultid="3348" />
                    <RANKING order="4" place="4" resultid="3901" />
                    <RANKING order="5" place="5" resultid="2680" />
                    <RANKING order="6" place="6" resultid="3480" />
                    <RANKING order="7" place="7" resultid="4420" />
                    <RANKING order="8" place="8" resultid="4555" />
                    <RANKING order="9" place="9" resultid="3238" />
                    <RANKING order="10" place="10" resultid="1958" />
                    <RANKING order="11" place="11" resultid="5341" />
                    <RANKING order="12" place="12" resultid="3726" />
                    <RANKING order="13" place="-1" resultid="4371" />
                    <RANKING order="14" place="-1" resultid="4668" />
                    <RANKING order="15" place="-1" resultid="5085" />
                    <RANKING order="16" place="-1" resultid="3372" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1210" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2512" />
                    <RANKING order="2" place="2" resultid="5364" />
                    <RANKING order="3" place="3" resultid="2181" />
                    <RANKING order="4" place="4" resultid="3356" />
                    <RANKING order="5" place="5" resultid="3519" />
                    <RANKING order="6" place="6" resultid="4548" />
                    <RANKING order="7" place="7" resultid="2306" />
                    <RANKING order="8" place="8" resultid="4484" />
                    <RANKING order="9" place="9" resultid="3292" />
                    <RANKING order="10" place="10" resultid="3028" />
                    <RANKING order="11" place="11" resultid="4034" />
                    <RANKING order="12" place="12" resultid="4299" />
                    <RANKING order="13" place="13" resultid="3458" />
                    <RANKING order="14" place="14" resultid="2188" />
                    <RANKING order="15" place="15" resultid="2700" />
                    <RANKING order="16" place="16" resultid="3503" />
                    <RANKING order="17" place="17" resultid="2185" />
                    <RANKING order="18" place="18" resultid="3112" />
                    <RANKING order="19" place="19" resultid="2578" />
                    <RANKING order="20" place="20" resultid="3860" />
                    <RANKING order="21" place="21" resultid="3229" />
                    <RANKING order="22" place="-1" resultid="4022" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1211" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3592" />
                    <RANKING order="2" place="2" resultid="4542" />
                    <RANKING order="3" place="3" resultid="5046" />
                    <RANKING order="4" place="4" resultid="3262" />
                    <RANKING order="5" place="5" resultid="3086" />
                    <RANKING order="6" place="6" resultid="4848" />
                    <RANKING order="7" place="7" resultid="5254" />
                    <RANKING order="8" place="8" resultid="4713" />
                    <RANKING order="9" place="9" resultid="2518" />
                    <RANKING order="10" place="10" resultid="5030" />
                    <RANKING order="11" place="11" resultid="2207" />
                    <RANKING order="12" place="12" resultid="2629" />
                    <RANKING order="13" place="-1" resultid="3935" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1212" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2557" />
                    <RANKING order="2" place="2" resultid="4204" />
                    <RANKING order="3" place="3" resultid="4027" />
                    <RANKING order="4" place="4" resultid="3895" />
                    <RANKING order="5" place="5" resultid="2998" />
                    <RANKING order="6" place="6" resultid="5357" />
                    <RANKING order="7" place="7" resultid="2600" />
                    <RANKING order="8" place="8" resultid="4245" />
                    <RANKING order="9" place="-1" resultid="5397" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1213" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4898" />
                    <RANKING order="2" place="2" resultid="3585" />
                    <RANKING order="3" place="3" resultid="2825" />
                    <RANKING order="4" place="4" resultid="4937" />
                    <RANKING order="5" place="5" resultid="2337" />
                    <RANKING order="6" place="6" resultid="5379" />
                    <RANKING order="7" place="7" resultid="4818" />
                    <RANKING order="8" place="8" resultid="4066" />
                    <RANKING order="9" place="9" resultid="3630" />
                    <RANKING order="10" place="10" resultid="4882" />
                    <RANKING order="11" place="11" resultid="2007" />
                    <RANKING order="12" place="12" resultid="2400" />
                    <RANKING order="13" place="13" resultid="4778" />
                    <RANKING order="14" place="14" resultid="3343" />
                    <RANKING order="15" place="15" resultid="3402" />
                    <RANKING order="16" place="16" resultid="3005" />
                    <RANKING order="17" place="17" resultid="4770" />
                    <RANKING order="18" place="-1" resultid="4925" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1214" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4292" />
                    <RANKING order="2" place="2" resultid="4005" />
                    <RANKING order="3" place="3" resultid="5250" />
                    <RANKING order="4" place="4" resultid="2889" />
                    <RANKING order="5" place="5" resultid="4504" />
                    <RANKING order="6" place="6" resultid="2583" />
                    <RANKING order="7" place="7" resultid="3831" />
                    <RANKING order="8" place="8" resultid="4699" />
                    <RANKING order="9" place="9" resultid="3142" />
                    <RANKING order="10" place="-1" resultid="5428" />
                    <RANKING order="11" place="-1" resultid="2429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1215" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4057" />
                    <RANKING order="2" place="2" resultid="2867" />
                    <RANKING order="3" place="3" resultid="2645" />
                    <RANKING order="4" place="4" resultid="2454" />
                    <RANKING order="5" place="5" resultid="5209" />
                    <RANKING order="6" place="-1" resultid="5215" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1216" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2368" />
                    <RANKING order="2" place="2" resultid="3604" />
                    <RANKING order="3" place="3" resultid="4116" />
                    <RANKING order="4" place="4" resultid="4123" />
                    <RANKING order="5" place="5" resultid="3126" />
                    <RANKING order="6" place="-1" resultid="4706" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1217" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4155" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1218" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4610" />
                    <RANKING order="2" place="2" resultid="3943" />
                    <RANKING order="3" place="3" resultid="2446" />
                    <RANKING order="4" place="4" resultid="2322" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1219" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4198" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1220" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1221" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6829" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6830" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6831" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6832" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6833" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6834" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6835" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6836" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6837" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6838" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6839" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="6840" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="6841" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="6842" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="6843" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="6844" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="6845" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="6846" number="18" order="18" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1222" daytime="10:19" gender="F" number="11" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1223" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2523" />
                    <RANKING order="2" place="2" resultid="2055" />
                    <RANKING order="3" place="3" resultid="5012" />
                    <RANKING order="4" place="-1" resultid="5444" />
                    <RANKING order="5" place="-1" resultid="5446" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1224" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3888" />
                    <RANKING order="2" place="2" resultid="2120" />
                    <RANKING order="3" place="3" resultid="2661" />
                    <RANKING order="4" place="4" resultid="4263" />
                    <RANKING order="5" place="5" resultid="4389" />
                    <RANKING order="6" place="6" resultid="4396" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1225" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2754" />
                    <RANKING order="2" place="2" resultid="3666" />
                    <RANKING order="3" place="3" resultid="2570" />
                    <RANKING order="4" place="4" resultid="3971" />
                    <RANKING order="5" place="-1" resultid="5390" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1226" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2624" />
                    <RANKING order="2" place="2" resultid="1946" />
                    <RANKING order="3" place="3" resultid="2782" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1227" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4590" />
                    <RANKING order="2" place="2" resultid="3570" />
                    <RANKING order="3" place="3" resultid="3496" />
                    <RANKING order="4" place="4" resultid="4729" />
                    <RANKING order="5" place="-1" resultid="2141" />
                    <RANKING order="6" place="-1" resultid="4651" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1228" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2108" />
                    <RANKING order="2" place="2" resultid="2612" />
                    <RANKING order="3" place="3" resultid="5181" />
                    <RANKING order="4" place="4" resultid="4164" />
                    <RANKING order="5" place="5" resultid="4277" />
                    <RANKING order="6" place="6" resultid="3172" />
                    <RANKING order="7" place="7" resultid="4932" />
                    <RANKING order="8" place="-1" resultid="4511" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1229" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2150" />
                    <RANKING order="2" place="2" resultid="1974" />
                    <RANKING order="3" place="3" resultid="5174" />
                    <RANKING order="4" place="4" resultid="3579" />
                    <RANKING order="5" place="5" resultid="2138" />
                    <RANKING order="6" place="6" resultid="5170" />
                    <RANKING order="7" place="7" resultid="2458" />
                    <RANKING order="8" place="8" resultid="1940" />
                    <RANKING order="9" place="-1" resultid="3297" />
                    <RANKING order="10" place="-1" resultid="1999" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1230" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3965" />
                    <RANKING order="2" place="2" resultid="2016" />
                    <RANKING order="3" place="-1" resultid="1992" />
                    <RANKING order="4" place="-1" resultid="3178" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1231" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2880" />
                    <RANKING order="2" place="2" resultid="2115" />
                    <RANKING order="3" place="3" resultid="2486" />
                    <RANKING order="4" place="4" resultid="5151" />
                    <RANKING order="5" place="5" resultid="3164" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1232" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2862" />
                    <RANKING order="2" place="2" resultid="1986" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1233" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4086" />
                    <RANKING order="2" place="2" resultid="4093" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1234" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3324" />
                    <RANKING order="2" place="2" resultid="4861" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1235" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1236" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2022" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1237" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1238" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6847" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6848" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6849" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6850" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6851" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6852" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6853" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1239" daytime="10:30" gender="M" number="12" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1240" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3840" />
                    <RANKING order="2" place="2" resultid="2966" />
                    <RANKING order="3" place="3" resultid="3815" />
                    <RANKING order="4" place="4" resultid="2068" />
                    <RANKING order="5" place="5" resultid="1863" />
                    <RANKING order="6" place="6" resultid="2076" />
                    <RANKING order="7" place="7" resultid="2084" />
                    <RANKING order="8" place="-1" resultid="3786" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1241" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2904" />
                    <RANKING order="2" place="2" resultid="2668" />
                    <RANKING order="3" place="3" resultid="2740" />
                    <RANKING order="4" place="4" resultid="5051" />
                    <RANKING order="5" place="5" resultid="2911" />
                    <RANKING order="6" place="6" resultid="2693" />
                    <RANKING order="7" place="7" resultid="4496" />
                    <RANKING order="8" place="8" resultid="2434" />
                    <RANKING order="9" place="-1" resultid="2736" />
                    <RANKING order="10" place="-1" resultid="5125" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1242" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2652" />
                    <RANKING order="2" place="2" resultid="4347" />
                    <RANKING order="3" place="3" resultid="4642" />
                    <RANKING order="4" place="4" resultid="5104" />
                    <RANKING order="5" place="5" resultid="3302" />
                    <RANKING order="6" place="6" resultid="4764" />
                    <RANKING order="7" place="7" resultid="3651" />
                    <RANKING order="8" place="8" resultid="2747" />
                    <RANKING order="9" place="9" resultid="4326" />
                    <RANKING order="10" place="10" resultid="4358" />
                    <RANKING order="11" place="11" resultid="4362" />
                    <RANKING order="12" place="-1" resultid="4795" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1243" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3511" />
                    <RANKING order="2" place="1" resultid="3427" />
                    <RANKING order="3" place="3" resultid="3071" />
                    <RANKING order="4" place="4" resultid="3373" />
                    <RANKING order="5" place="5" resultid="2223" />
                    <RANKING order="6" place="6" resultid="3850" />
                    <RANKING order="7" place="7" resultid="3434" />
                    <RANKING order="8" place="8" resultid="2239" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1244" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2294" />
                    <RANKING order="2" place="2" resultid="5385" />
                    <RANKING order="3" place="3" resultid="2634" />
                    <RANKING order="4" place="3" resultid="5334" />
                    <RANKING order="5" place="5" resultid="3357" />
                    <RANKING order="6" place="6" resultid="4626" />
                    <RANKING order="7" place="7" resultid="3741" />
                    <RANKING order="8" place="8" resultid="3861" />
                    <RANKING order="9" place="9" resultid="5262" />
                    <RANKING order="10" place="10" resultid="5081" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1245" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3593" />
                    <RANKING order="2" place="2" resultid="5255" />
                    <RANKING order="3" place="3" resultid="3263" />
                    <RANKING order="4" place="4" resultid="3701" />
                    <RANKING order="5" place="5" resultid="2562" />
                    <RANKING order="6" place="6" resultid="4536" />
                    <RANKING order="7" place="7" resultid="4488" />
                    <RANKING order="8" place="8" resultid="2194" />
                    <RANKING order="9" place="9" resultid="4659" />
                    <RANKING order="10" place="10" resultid="4239" />
                    <RANKING order="11" place="11" resultid="5273" />
                    <RANKING order="12" place="12" resultid="1889" />
                    <RANKING order="13" place="13" resultid="3338" />
                    <RANKING order="14" place="14" resultid="2215" />
                    <RANKING order="15" place="15" resultid="2630" />
                    <RANKING order="16" place="-1" resultid="2549" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1246" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2478" />
                    <RANKING order="2" place="2" resultid="5392" />
                    <RANKING order="3" place="3" resultid="4824" />
                    <RANKING order="4" place="4" resultid="3474" />
                    <RANKING order="5" place="5" resultid="3911" />
                    <RANKING order="6" place="6" resultid="3096" />
                    <RANKING order="7" place="7" resultid="4530" />
                    <RANKING order="8" place="8" resultid="4226" />
                    <RANKING order="9" place="9" resultid="5329" />
                    <RANKING order="10" place="10" resultid="4246" />
                    <RANKING order="11" place="11" resultid="3394" />
                    <RANKING order="12" place="-1" resultid="4889" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1247" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3060" />
                    <RANKING order="2" place="2" resultid="4186" />
                    <RANKING order="3" place="3" resultid="3386" />
                    <RANKING order="4" place="4" resultid="4685" />
                    <RANKING order="5" place="5" resultid="4938" />
                    <RANKING order="6" place="6" resultid="3625" />
                    <RANKING order="7" place="7" resultid="3631" />
                    <RANKING order="8" place="8" resultid="2401" />
                    <RANKING order="9" place="9" resultid="3753" />
                    <RANKING order="10" place="9" resultid="4527" />
                    <RANKING order="11" place="11" resultid="3680" />
                    <RANKING order="12" place="12" resultid="3150" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1248" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4193" />
                    <RANKING order="2" place="2" resultid="4293" />
                    <RANKING order="3" place="3" resultid="3951" />
                    <RANKING order="4" place="4" resultid="3832" />
                    <RANKING order="5" place="5" resultid="2584" />
                    <RANKING order="6" place="6" resultid="2229" />
                    <RANKING order="7" place="-1" resultid="2408" />
                    <RANKING order="8" place="-1" resultid="5117" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1249" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2868" />
                    <RANKING order="2" place="2" resultid="5349" />
                    <RANKING order="3" place="3" resultid="2348" />
                    <RANKING order="4" place="4" resultid="3281" />
                    <RANKING order="5" place="5" resultid="3618" />
                    <RANKING order="6" place="6" resultid="5216" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1250" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2842" />
                    <RANKING order="2" place="2" resultid="1924" />
                    <RANKING order="3" place="3" resultid="3131" />
                    <RANKING order="4" place="4" resultid="5200" />
                    <RANKING order="5" place="5" resultid="4507" />
                    <RANKING order="6" place="6" resultid="4117" />
                    <RANKING order="7" place="-1" resultid="4124" />
                    <RANKING order="8" place="-1" resultid="4707" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1251" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3946" />
                    <RANKING order="2" place="2" resultid="5191" />
                    <RANKING order="3" place="3" resultid="1980" />
                    <RANKING order="4" place="-1" resultid="5196" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1252" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1253" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1254" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1255" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6854" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6855" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6856" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6857" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6858" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6859" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6860" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6861" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6862" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6863" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6864" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="6865" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="6866" number="13" order="13" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1256" daytime="10:47" gender="F" number="13" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1257" agemax="24" agemin="20" />
                <AGEGROUP agegroupid="1258" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1965" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1259" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3972" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1260" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="1261" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="1262" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2990" />
                    <RANKING order="2" place="2" resultid="2732" />
                    <RANKING order="3" place="3" resultid="3275" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1263" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4515" />
                    <RANKING order="2" place="2" resultid="2125" />
                    <RANKING order="3" place="3" resultid="2000" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1264" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1265" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="1266" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2847" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1267" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1268" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1269" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1270" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1271" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1272" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6867" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6868" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1273" daytime="10:57" gender="M" number="14" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1274" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4915" />
                    <RANKING order="2" place="2" resultid="1869" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1275" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4413" />
                    <RANKING order="2" place="2" resultid="3873" />
                    <RANKING order="3" place="3" resultid="5130" />
                    <RANKING order="4" place="4" resultid="4599" />
                    <RANKING order="5" place="5" resultid="4212" />
                    <RANKING order="6" place="6" resultid="2768" />
                    <RANKING order="7" place="7" resultid="2694" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1276" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4378" />
                    <RANKING order="2" place="2" resultid="3443" />
                    <RANKING order="3" place="3" resultid="4311" />
                    <RANKING order="4" place="4" resultid="5074" />
                    <RANKING order="5" place="5" resultid="4072" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1277" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2202" />
                    <RANKING order="2" place="2" resultid="3435" />
                    <RANKING order="3" place="3" resultid="5342" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1278" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2295" />
                    <RANKING order="2" place="2" resultid="2172" />
                    <RANKING order="3" place="3" resultid="5335" />
                    <RANKING order="4" place="4" resultid="3459" />
                    <RANKING order="5" place="5" resultid="4140" />
                    <RANKING order="6" place="6" resultid="4721" />
                    <RANKING order="7" place="-1" resultid="3218" />
                    <RANKING order="8" place="-1" resultid="3504" />
                    <RANKING order="9" place="-1" resultid="4014" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1279" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3285" />
                    <RANKING order="2" place="2" resultid="3309" />
                    <RANKING order="3" place="3" resultid="5031" />
                    <RANKING order="4" place="4" resultid="4219" />
                    <RANKING order="5" place="-1" resultid="2550" />
                    <RANKING order="6" place="-1" resultid="3936" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1280" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3912" />
                    <RANKING order="2" place="2" resultid="3466" />
                    <RANKING order="3" place="-1" resultid="3709" />
                    <RANKING order="4" place="-1" resultid="4205" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1281" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2352" />
                    <RANKING order="2" place="2" resultid="2809" />
                    <RANKING order="3" place="3" resultid="3365" />
                    <RANKING order="4" place="4" resultid="2338" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1282" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2714" />
                    <RANKING order="2" place="2" resultid="5227" />
                    <RANKING order="3" place="3" resultid="4428" />
                    <RANKING order="4" place="4" resultid="2464" />
                    <RANKING order="5" place="5" resultid="4968" />
                    <RANKING order="6" place="6" resultid="3377" />
                    <RANKING order="7" place="-1" resultid="3612" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1283" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4058" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1284" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4691" />
                    <RANKING order="2" place="2" resultid="3132" />
                    <RANKING order="3" place="3" resultid="2530" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1285" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1286" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1287" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1288" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1289" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6869" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6870" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6871" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6872" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6873" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6874" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1290" daytime="11:22" gender="F" number="15" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1291" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2417" />
                    <RANKING order="2" place="2" resultid="2061" />
                    <RANKING order="3" place="3" resultid="3658" />
                    <RANKING order="4" place="4" resultid="2524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1292" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2917" />
                    <RANKING order="2" place="2" resultid="3805" />
                    <RANKING order="3" place="3" resultid="2724" />
                    <RANKING order="4" place="4" resultid="4390" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1293" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4831" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1294" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2165" />
                    <RANKING order="2" place="2" resultid="1854" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1295" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2344" />
                    <RANKING order="2" place="2" resultid="2142" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1296" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2471" />
                    <RANKING order="2" place="2" resultid="3079" />
                    <RANKING order="3" place="3" resultid="2733" />
                    <RANKING order="4" place="4" resultid="4172" />
                    <RANKING order="5" place="5" resultid="4977" />
                    <RANKING order="6" place="6" resultid="5038" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1297" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5175" />
                    <RANKING order="2" place="2" resultid="1932" />
                    <RANKING order="3" place="3" resultid="2126" />
                    <RANKING order="4" place="4" resultid="1917" />
                    <RANKING order="5" place="5" resultid="1952" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1298" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3737" />
                    <RANKING order="2" place="2" resultid="4637" />
                    <RANKING order="3" place="3" resultid="5162" />
                    <RANKING order="4" place="-1" resultid="3179" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1299" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2854" />
                    <RANKING order="2" place="2" resultid="3961" />
                    <RANKING order="3" place="3" resultid="2501" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1300" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4962" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1301" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4842" />
                    <RANKING order="2" place="2" resultid="4087" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1302" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2607" />
                    <RANKING order="2" place="2" resultid="4866" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1303" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3104" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1304" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1305" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1306" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6875" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6876" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6877" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6878" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6879" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1307" daytime="11:49" gender="M" number="16" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1308" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2091" />
                    <RANKING order="2" place="2" resultid="5097" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1309" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2329" />
                    <RANKING order="2" place="2" resultid="2951" />
                    <RANKING order="3" place="3" resultid="5052" />
                    <RANKING order="4" place="4" resultid="2741" />
                    <RANKING order="5" place="5" resultid="2425" />
                    <RANKING order="6" place="6" resultid="2940" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1310" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3303" />
                    <RANKING order="2" place="2" resultid="3673" />
                    <RANKING order="3" place="3" resultid="5066" />
                    <RANKING order="4" place="4" resultid="5105" />
                    <RANKING order="5" place="5" resultid="3488" />
                    <RANKING order="6" place="6" resultid="4320" />
                    <RANKING order="7" place="7" resultid="4341" />
                    <RANKING order="8" place="-1" resultid="4148" />
                    <RANKING order="9" place="-1" resultid="6702" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1311" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3419" />
                    <RANKING order="2" place="2" resultid="3512" />
                    <RANKING order="3" place="3" resultid="2681" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1312" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2617" />
                    <RANKING order="2" place="2" resultid="4549" />
                    <RANKING order="3" place="3" resultid="3029" />
                    <RANKING order="4" place="4" resultid="4050" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1313" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2563" />
                    <RANKING order="2" place="2" resultid="4849" />
                    <RANKING order="3" place="3" resultid="2195" />
                    <RANKING order="4" place="4" resultid="1890" />
                    <RANKING order="5" place="5" resultid="4660" />
                    <RANKING order="6" place="6" resultid="5088" />
                    <RANKING order="7" place="-1" resultid="2216" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1314" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2707" />
                    <RANKING order="2" place="2" resultid="4078" />
                    <RANKING order="3" place="3" resultid="3097" />
                    <RANKING order="4" place="4" resultid="5241" />
                    <RANKING order="5" place="5" resultid="3395" />
                    <RANKING order="6" place="6" resultid="3731" />
                    <RANKING order="7" place="7" resultid="5398" />
                    <RANKING order="8" place="-1" resultid="3036" />
                    <RANKING order="9" place="-1" resultid="4890" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1315" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4899" />
                    <RANKING order="2" place="2" resultid="4617" />
                    <RANKING order="3" place="3" resultid="5380" />
                    <RANKING order="4" place="4" resultid="4883" />
                    <RANKING order="5" place="5" resultid="4187" />
                    <RANKING order="6" place="6" resultid="3006" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1316" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2360" />
                    <RANKING order="2" place="2" resultid="3450" />
                    <RANKING order="3" place="3" resultid="2831" />
                    <RANKING order="4" place="4" resultid="4429" />
                    <RANKING order="5" place="5" resultid="4969" />
                    <RANKING order="6" place="6" resultid="2409" />
                    <RANKING order="7" place="7" resultid="3378" />
                    <RANKING order="8" place="8" resultid="3613" />
                    <RANKING order="9" place="9" resultid="3143" />
                    <RANKING order="10" place="-1" resultid="5234" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1317" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5221" />
                    <RANKING order="2" place="2" resultid="5350" />
                    <RANKING order="3" place="-1" resultid="3990" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1318" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2369" />
                    <RANKING order="2" place="2" resultid="2531" />
                    <RANKING order="3" place="3" resultid="4692" />
                    <RANKING order="4" place="-1" resultid="1925" />
                    <RANKING order="5" place="-1" resultid="3605" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1319" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4108" />
                    <RANKING order="2" place="2" resultid="4156" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1320" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1321" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1322" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1323" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6880" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6881" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6882" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6883" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6884" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6885" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6886" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6887" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1324" daytime="12:23" gender="F" number="17" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1392" agemax="96" agemin="80" />
                <AGEGROUP agegroupid="1393" agemax="119" agemin="100">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2971" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1394" agemax="159" agemin="120">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2792" />
                    <RANKING order="2" place="2" resultid="6977" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1395" agemax="199" agemin="160">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2254" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1396" agemax="239" agemin="200">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2245" />
                    <RANKING order="2" place="2" resultid="5295" />
                    <RANKING order="3" place="3" resultid="4983" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1397" agemax="279" agemin="240">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2034" />
                    <RANKING order="2" place="2" resultid="3187" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1398" agemax="319" agemin="280" />
                <AGEGROUP agegroupid="1399" agemax="359" agemin="320" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6979" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1341" daytime="12:31" gender="M" number="18" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1400" agemax="96" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3794" />
                    <RANKING order="2" place="2" resultid="2096" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1401" agemax="119" agemin="100">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2974" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1402" agemax="159" agemin="120">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6982" />
                    <RANKING order="2" place="2" resultid="6660" />
                    <RANKING order="3" place="3" resultid="3528" />
                    <RANKING order="4" place="4" resultid="2793" />
                    <RANKING order="5" place="5" resultid="6981" />
                    <RANKING order="6" place="6" resultid="4405" />
                    <RANKING order="7" place="7" resultid="3878" />
                    <RANKING order="8" place="8" resultid="3685" />
                    <RANKING order="9" place="9" resultid="4404" />
                    <RANKING order="10" place="10" resultid="6661" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1403" agemax="199" agemin="160">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2256" />
                    <RANKING order="2" place="2" resultid="4568" />
                    <RANKING order="3" place="3" resultid="4875" />
                    <RANKING order="4" place="4" resultid="3529" />
                    <RANKING order="5" place="5" resultid="2255" />
                    <RANKING order="6" place="6" resultid="6980" />
                    <RANKING order="7" place="7" resultid="4252" />
                    <RANKING order="8" place="8" resultid="6983" />
                    <RANKING order="9" place="-1" resultid="3042" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1404" agemax="239" agemin="200">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3530" />
                    <RANKING order="2" place="2" resultid="5290" />
                    <RANKING order="3" place="3" resultid="4984" />
                    <RANKING order="4" place="4" resultid="6984" />
                    <RANKING order="5" place="-1" resultid="4570" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1405" agemax="279" agemin="240">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2381" />
                    <RANKING order="2" place="2" resultid="5292" />
                    <RANKING order="3" place="3" resultid="3686" />
                    <RANKING order="4" place="4" resultid="4742" />
                    <RANKING order="5" place="-1" resultid="3189" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1406" agemax="319" agemin="280" />
                <AGEGROUP agegroupid="1407" agemax="359" agemin="320" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6985" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6986" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6987" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6988" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1358" daytime="12:44" gender="F" number="19" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1359" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2418" />
                    <RANKING order="2" place="2" resultid="3659" />
                    <RANKING order="3" place="3" resultid="3270" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1360" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4631" />
                    <RANKING order="2" place="2" resultid="2725" />
                    <RANKING order="3" place="3" resultid="3224" />
                    <RANKING order="4" place="4" resultid="3119" />
                    <RANKING order="5" place="5" resultid="1966" />
                    <RANKING order="6" place="6" resultid="4264" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1361" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3054" />
                    <RANKING order="2" place="2" resultid="2761" />
                    <RANKING order="3" place="3" resultid="2571" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1362" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2837" />
                    <RANKING order="2" place="2" resultid="3985" />
                    <RANKING order="3" place="3" resultid="2166" />
                    <RANKING order="4" place="4" resultid="5373" />
                    <RANKING order="5" place="-1" resultid="1855" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1363" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3823" />
                    <RANKING order="2" place="-1" resultid="3571" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1364" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3320" />
                    <RANKING order="2" place="2" resultid="2991" />
                    <RANKING order="3" place="3" resultid="2158" />
                    <RANKING order="4" place="4" resultid="2472" />
                    <RANKING order="5" place="5" resultid="5039" />
                    <RANKING order="6" place="6" resultid="4165" />
                    <RANKING order="7" place="7" resultid="4278" />
                    <RANKING order="8" place="8" resultid="3276" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1365" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4516" />
                    <RANKING order="2" place="2" resultid="1933" />
                    <RANKING order="3" place="3" resultid="3066" />
                    <RANKING order="4" place="-1" resultid="2491" />
                    <RANKING order="5" place="-1" resultid="3580" />
                    <RANKING order="6" place="-1" resultid="1953" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1366" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4272" />
                    <RANKING order="2" place="2" resultid="4179" />
                    <RANKING order="3" place="3" resultid="4101" />
                    <RANKING order="4" place="4" resultid="3738" />
                    <RANKING order="5" place="5" resultid="2393" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1367" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2675" />
                    <RANKING order="2" place="2" resultid="2502" />
                    <RANKING order="3" place="3" resultid="3213" />
                    <RANKING order="4" place="-1" resultid="4950" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1368" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4957" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1369" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4843" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1370" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4867" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1371" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1372" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1373" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1374" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6894" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6895" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6896" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6897" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6898" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1375" daytime="13:27" gender="M" number="20" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1376" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2440" />
                    <RANKING order="2" place="2" resultid="4916" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1377" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4857" />
                    <RANKING order="2" place="2" resultid="2330" />
                    <RANKING order="3" place="3" resultid="5131" />
                    <RANKING order="4" place="4" resultid="4497" />
                    <RANKING order="5" place="5" resultid="4758" />
                    <RANKING order="6" place="-1" resultid="2769" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1378" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3021" />
                    <RANKING order="2" place="2" resultid="5059" />
                    <RANKING order="3" place="3" resultid="4312" />
                    <RANKING order="4" place="4" resultid="4643" />
                    <RANKING order="5" place="5" resultid="3746" />
                    <RANKING order="6" place="6" resultid="3489" />
                    <RANKING order="7" place="7" resultid="3643" />
                    <RANKING order="8" place="8" resultid="2539" />
                    <RANKING order="9" place="9" resultid="5075" />
                    <RANKING order="10" place="-1" resultid="5067" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1379" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3349" />
                    <RANKING order="2" place="2" resultid="3329" />
                    <RANKING order="3" place="3" resultid="3481" />
                    <RANKING order="4" place="4" resultid="3239" />
                    <RANKING order="5" place="5" resultid="4556" />
                    <RANKING order="6" place="6" resultid="4372" />
                    <RANKING order="7" place="7" resultid="2050" />
                    <RANKING order="8" place="8" resultid="4669" />
                    <RANKING order="9" place="9" resultid="3727" />
                    <RANKING order="10" place="-1" resultid="3902" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1380" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5365" />
                    <RANKING order="2" place="2" resultid="4041" />
                    <RANKING order="3" place="3" resultid="3520" />
                    <RANKING order="4" place="4" resultid="3293" />
                    <RANKING order="5" place="5" resultid="2701" />
                    <RANKING order="6" place="6" resultid="4035" />
                    <RANKING order="7" place="7" resultid="4015" />
                    <RANKING order="8" place="8" resultid="4141" />
                    <RANKING order="9" place="9" resultid="4722" />
                    <RANKING order="10" place="10" resultid="3113" />
                    <RANKING order="11" place="11" resultid="2579" />
                    <RANKING order="12" place="12" resultid="2211" />
                    <RANKING order="13" place="13" resultid="3230" />
                    <RANKING order="14" place="14" resultid="4051" />
                    <RANKING order="15" place="15" resultid="2234" />
                    <RANKING order="16" place="-1" resultid="2513" />
                    <RANKING order="17" place="-1" resultid="4300" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1381" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3702" />
                    <RANKING order="2" place="2" resultid="2519" />
                    <RANKING order="3" place="3" resultid="5089" />
                    <RANKING order="4" place="-1" resultid="3339" />
                    <RANKING order="5" place="-1" resultid="2595" />
                    <RANKING order="6" place="-1" resultid="3286" />
                    <RANKING order="7" place="-1" resultid="5256" />
                    <RANKING order="8" place="-1" resultid="4714" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1382" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3037" />
                    <RANKING order="2" place="2" resultid="5246" />
                    <RANKING order="3" place="3" resultid="3710" />
                    <RANKING order="4" place="4" resultid="4028" />
                    <RANKING order="5" place="5" resultid="2999" />
                    <RANKING order="6" place="6" resultid="3564" />
                    <RANKING order="7" place="7" resultid="4945" />
                    <RANKING order="8" place="8" resultid="2601" />
                    <RANKING order="9" place="-1" resultid="5358" />
                    <RANKING order="10" place="-1" resultid="3467" />
                    <RANKING order="11" place="-1" resultid="3896" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1383" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2008" />
                    <RANKING order="2" place="2" resultid="4067" />
                    <RANKING order="3" place="3" resultid="2810" />
                    <RANKING order="4" place="4" resultid="2826" />
                    <RANKING order="5" place="5" resultid="2353" />
                    <RANKING order="6" place="6" resultid="3366" />
                    <RANKING order="7" place="7" resultid="4926" />
                    <RANKING order="8" place="8" resultid="3403" />
                    <RANKING order="9" place="9" resultid="4779" />
                    <RANKING order="10" place="10" resultid="3387" />
                    <RANKING order="11" place="11" resultid="3754" />
                    <RANKING order="12" place="12" resultid="4771" />
                    <RANKING order="13" place="-1" resultid="3151" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1384" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4006" />
                    <RANKING order="2" place="2" resultid="2361" />
                    <RANKING order="3" place="3" resultid="3451" />
                    <RANKING order="4" place="4" resultid="3718" />
                    <RANKING order="5" place="5" resultid="4505" />
                    <RANKING order="6" place="6" resultid="2465" />
                    <RANKING order="7" place="7" resultid="4700" />
                    <RANKING order="8" place="-1" resultid="4753" />
                    <RANKING order="9" place="-1" resultid="5118" />
                    <RANKING order="10" place="-1" resultid="5429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1385" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2646" />
                    <RANKING order="2" place="-1" resultid="3991" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1386" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3999" />
                    <RANKING order="2" place="-1" resultid="3127" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1387" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4109" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1388" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4611" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1389" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4199" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1390" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1391" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6899" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6900" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6901" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6902" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6903" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6904" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6905" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6906" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6907" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6908" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6909" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2011-11-19" daytime="15:30" number="3">
          <EVENTS>
            <EVENT eventid="1409" daytime="15:30" gender="F" number="21" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1413" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2525" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1414" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2121" />
                    <RANKING order="2" place="2" resultid="2662" />
                    <RANKING order="3" place="3" resultid="4391" />
                    <RANKING order="4" place="4" resultid="4397" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1415" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2755" />
                    <RANKING order="2" place="2" resultid="3667" />
                    <RANKING order="3" place="3" resultid="2572" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1416" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2838" />
                    <RANKING order="2" place="2" resultid="2625" />
                    <RANKING order="3" place="3" resultid="5188" />
                    <RANKING order="4" place="4" resultid="1947" />
                    <RANKING order="5" place="-1" resultid="2783" />
                    <RANKING order="6" place="-1" resultid="1856" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1417" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3824" />
                    <RANKING order="2" place="2" resultid="4730" />
                    <RANKING order="3" place="-1" resultid="3497" />
                    <RANKING order="4" place="-1" resultid="4652" />
                    <RANKING order="5" place="-1" resultid="2143" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1418" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2613" />
                    <RANKING order="2" place="2" resultid="4279" />
                    <RANKING order="3" place="3" resultid="3173" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1419" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2151" />
                    <RANKING order="2" place="2" resultid="1954" />
                    <RANKING order="3" place="3" resultid="2001" />
                    <RANKING order="4" place="4" resultid="3298" />
                    <RANKING order="5" place="-1" resultid="4082" />
                    <RANKING order="6" place="-1" resultid="1941" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1420" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2017" />
                    <RANKING order="2" place="2" resultid="1994" />
                    <RANKING order="3" place="-1" resultid="3180" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1421" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2487" />
                    <RANKING order="2" place="2" resultid="3962" />
                    <RANKING order="3" place="3" resultid="2116" />
                    <RANKING order="4" place="4" resultid="3165" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1422" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2848" />
                    <RANKING order="2" place="2" resultid="1987" />
                    <RANKING order="3" place="3" resultid="4963" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1423" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1424" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3325" />
                    <RANKING order="2" place="2" resultid="4862" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1425" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3105" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1426" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2023" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1427" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1428" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6997" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6998" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6999" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7000" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7001" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1411" daytime="16:01" gender="M" number="22" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1429" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2967" />
                    <RANKING order="2" place="2" resultid="3787" />
                    <RANKING order="3" place="3" resultid="1870" />
                    <RANKING order="4" place="-1" resultid="3816" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1430" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2905" />
                    <RANKING order="2" place="2" resultid="2669" />
                    <RANKING order="3" place="3" resultid="2912" />
                    <RANKING order="4" place="4" resultid="4498" />
                    <RANKING order="5" place="5" resultid="2695" />
                    <RANKING order="6" place="6" resultid="2435" />
                    <RANKING order="7" place="-1" resultid="2737" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1431" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5139" />
                    <RANKING order="2" place="2" resultid="4348" />
                    <RANKING order="3" place="3" resultid="4644" />
                    <RANKING order="4" place="4" resultid="3444" />
                    <RANKING order="5" place="5" resultid="3490" />
                    <RANKING order="6" place="6" resultid="5106" />
                    <RANKING order="7" place="7" resultid="4327" />
                    <RANKING order="8" place="-1" resultid="4149" />
                    <RANKING order="9" place="-1" resultid="2653" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1432" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3513" />
                    <RANKING order="2" place="2" resultid="2240" />
                    <RANKING order="3" place="3" resultid="3436" />
                    <RANKING order="4" place="-1" resultid="3072" />
                    <RANKING order="5" place="-1" resultid="3852" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1433" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2296" />
                    <RANKING order="2" place="2" resultid="5386" />
                    <RANKING order="3" place="3" resultid="3358" />
                    <RANKING order="4" place="4" resultid="3742" />
                    <RANKING order="5" place="5" resultid="4142" />
                    <RANKING order="6" place="6" resultid="3460" />
                    <RANKING order="7" place="7" resultid="2635" />
                    <RANKING order="8" place="8" resultid="4627" />
                    <RANKING order="9" place="9" resultid="3030" />
                    <RANKING order="10" place="-1" resultid="5082" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1434" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3594" />
                    <RANKING order="2" place="2" resultid="5257" />
                    <RANKING order="3" place="3" resultid="4489" />
                    <RANKING order="4" place="4" resultid="4661" />
                    <RANKING order="5" place="5" resultid="4537" />
                    <RANKING order="6" place="6" resultid="3310" />
                    <RANKING order="7" place="7" resultid="3340" />
                    <RANKING order="8" place="8" resultid="2631" />
                    <RANKING order="9" place="-1" resultid="2217" />
                    <RANKING order="10" place="-1" resultid="2551" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1435" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5393" />
                    <RANKING order="2" place="2" resultid="4825" />
                    <RANKING order="3" place="3" resultid="3098" />
                    <RANKING order="4" place="4" resultid="3475" />
                    <RANKING order="5" place="5" resultid="5330" />
                    <RANKING order="6" place="6" resultid="2602" />
                    <RANKING order="7" place="-1" resultid="4227" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1436" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3061" />
                    <RANKING order="2" place="2" resultid="4188" />
                    <RANKING order="3" place="3" resultid="4686" />
                    <RANKING order="4" place="4" resultid="4939" />
                    <RANKING order="5" place="5" resultid="2009" />
                    <RANKING order="6" place="6" resultid="2402" />
                    <RANKING order="7" place="7" resultid="3626" />
                    <RANKING order="8" place="8" resultid="3388" />
                    <RANKING order="9" place="9" resultid="3404" />
                    <RANKING order="10" place="10" resultid="3007" />
                    <RANKING order="11" place="11" resultid="3152" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1437" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4194" />
                    <RANKING order="2" place="2" resultid="2715" />
                    <RANKING order="3" place="3" resultid="5228" />
                    <RANKING order="4" place="4" resultid="3452" />
                    <RANKING order="5" place="5" resultid="3952" />
                    <RANKING order="6" place="6" resultid="4701" />
                    <RANKING order="7" place="7" resultid="3833" />
                    <RANKING order="8" place="8" resultid="2410" />
                    <RANKING order="9" place="9" resultid="3614" />
                    <RANKING order="10" place="10" resultid="2230" />
                    <RANKING order="11" place="-1" resultid="2430" />
                    <RANKING order="12" place="-1" resultid="2466" />
                    <RANKING order="13" place="-1" resultid="5119" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1438" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5351" />
                    <RANKING order="2" place="2" resultid="3619" />
                    <RANKING order="3" place="3" resultid="3282" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1439" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2843" />
                    <RANKING order="2" place="2" resultid="1926" />
                    <RANKING order="3" place="3" resultid="3133" />
                    <RANKING order="4" place="4" resultid="4508" />
                    <RANKING order="5" place="5" resultid="2532" />
                    <RANKING order="6" place="-1" resultid="4118" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1440" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3947" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1441" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1442" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1443" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1444" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7002" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7003" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7004" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7005" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7006" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7007" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7008" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7009" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7010" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7011" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1445" daytime="16:47" gender="F" number="23" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1446" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4872" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1447" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1877" />
                    <RANKING order="2" place="2" resultid="2957" />
                    <RANKING order="3" place="3" resultid="1967" />
                    <RANKING order="4" place="4" resultid="2962" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1448" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4809" />
                    <RANKING order="2" place="2" resultid="3973" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1449" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="1450" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3572" />
                    <RANKING order="2" place="-1" resultid="4591" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1451" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2992" />
                    <RANKING order="2" place="2" resultid="2159" />
                    <RANKING order="3" place="3" resultid="3277" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1452" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4517" />
                    <RANKING order="2" place="2" resultid="1975" />
                    <RANKING order="3" place="3" resultid="2127" />
                    <RANKING order="4" place="4" resultid="2002" />
                    <RANKING order="5" place="5" resultid="3411" />
                    <RANKING order="6" place="-1" resultid="1934" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1453" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2018" />
                    <RANKING order="2" place="2" resultid="5163" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1454" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3957" />
                    <RANKING order="2" place="-1" resultid="4951" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1455" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2849" />
                    <RANKING order="2" place="2" resultid="4958" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1456" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1457" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1458" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1459" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1460" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1461" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7012" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7013" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7014" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1462" daytime="16:56" gender="M" number="24" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1463" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3791" />
                    <RANKING order="2" place="2" resultid="4917" />
                    <RANKING order="3" place="3" resultid="2069" />
                    <RANKING order="4" place="4" resultid="2077" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1464" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4414" />
                    <RANKING order="2" place="2" resultid="3874" />
                    <RANKING order="3" place="3" resultid="1883" />
                    <RANKING order="4" place="4" resultid="5053" />
                    <RANKING order="5" place="5" resultid="3245" />
                    <RANKING order="6" place="6" resultid="2928" />
                    <RANKING order="7" place="7" resultid="5132" />
                    <RANKING order="8" place="8" resultid="2770" />
                    <RANKING order="9" place="9" resultid="3207" />
                    <RANKING order="10" place="-1" resultid="4213" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1465" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2544" />
                    <RANKING order="2" place="2" resultid="4379" />
                    <RANKING order="3" place="3" resultid="5060" />
                    <RANKING order="4" place="4" resultid="5068" />
                    <RANKING order="5" place="5" resultid="2748" />
                    <RANKING order="6" place="6" resultid="3644" />
                    <RANKING order="7" place="7" resultid="5076" />
                    <RANKING order="8" place="-1" resultid="3747" />
                    <RANKING order="9" place="-1" resultid="4313" />
                    <RANKING order="10" place="-1" resultid="4353" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1466" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3428" />
                    <RANKING order="2" place="2" resultid="2203" />
                    <RANKING order="3" place="3" resultid="3240" />
                    <RANKING order="4" place="4" resultid="3482" />
                    <RANKING order="5" place="5" resultid="5278" />
                    <RANKING order="6" place="6" resultid="5343" />
                    <RANKING order="7" place="7" resultid="2316" />
                    <RANKING order="8" place="8" resultid="4670" />
                    <RANKING order="9" place="-1" resultid="1959" />
                    <RANKING order="10" place="-1" resultid="4421" />
                    <RANKING order="11" place="-1" resultid="4557" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1467" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2618" />
                    <RANKING order="2" place="2" resultid="3219" />
                    <RANKING order="3" place="3" resultid="2173" />
                    <RANKING order="4" place="4" resultid="2297" />
                    <RANKING order="5" place="5" resultid="3521" />
                    <RANKING order="6" place="6" resultid="5336" />
                    <RANKING order="7" place="7" resultid="3862" />
                    <RANKING order="8" place="8" resultid="4016" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1468" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3287" />
                    <RANKING order="2" place="2" resultid="3087" />
                    <RANKING order="3" place="3" resultid="2196" />
                    <RANKING order="4" place="4" resultid="5032" />
                    <RANKING order="5" place="5" resultid="4715" />
                    <RANKING order="6" place="-1" resultid="2552" />
                    <RANKING order="7" place="-1" resultid="4220" />
                    <RANKING order="8" place="-1" resultid="3937" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1469" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4206" />
                    <RANKING order="2" place="2" resultid="3913" />
                    <RANKING order="3" place="3" resultid="3711" />
                    <RANKING order="4" place="4" resultid="3565" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1470" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2354" />
                    <RANKING order="2" place="2" resultid="5381" />
                    <RANKING order="3" place="3" resultid="4819" />
                    <RANKING order="4" place="4" resultid="2339" />
                    <RANKING order="5" place="5" resultid="2811" />
                    <RANKING order="6" place="6" resultid="3367" />
                    <RANKING order="7" place="7" resultid="3632" />
                    <RANKING order="8" place="8" resultid="2403" />
                    <RANKING order="9" place="9" resultid="3681" />
                    <RANKING order="10" place="-1" resultid="4780" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1471" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2362" />
                    <RANKING order="2" place="2" resultid="4430" />
                    <RANKING order="3" place="3" resultid="4970" />
                    <RANKING order="4" place="4" resultid="3379" />
                    <RANKING order="5" place="5" resultid="3144" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1472" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4059" />
                    <RANKING order="2" place="-1" resultid="3992" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1473" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3134" />
                    <RANKING order="2" place="2" resultid="4693" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1474" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1475" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1476" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1477" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1478" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7015" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7016" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7017" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7018" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7019" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7020" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7021" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7022" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7023" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1479" daytime="17:14" gender="F" number="25" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1480" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2419" />
                    <RANKING order="2" place="2" resultid="2062" />
                    <RANKING order="3" place="3" resultid="2056" />
                    <RANKING order="4" place="4" resultid="2526" />
                    <RANKING order="5" place="5" resultid="3979" />
                    <RANKING order="6" place="6" resultid="2031" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1481" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3889" />
                    <RANKING order="2" place="2" resultid="2918" />
                    <RANKING order="3" place="3" resultid="3806" />
                    <RANKING order="4" place="4" resultid="2726" />
                    <RANKING order="5" place="5" resultid="3120" />
                    <RANKING order="6" place="6" resultid="4265" />
                    <RANKING order="7" place="-1" resultid="1968" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1482" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3252" />
                    <RANKING order="2" place="2" resultid="3256" />
                    <RANKING order="3" place="3" resultid="4385" />
                    <RANKING order="4" place="4" resultid="2640" />
                    <RANKING order="5" place="5" resultid="4832" />
                    <RANKING order="6" place="6" resultid="3668" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1483" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2302" />
                    <RANKING order="2" place="2" resultid="2687" />
                    <RANKING order="3" place="3" resultid="2167" />
                    <RANKING order="4" place="4" resultid="5284" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1484" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4592" />
                    <RANKING order="2" place="2" resultid="2345" />
                    <RANKING order="3" place="3" resultid="2144" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1485" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2109" />
                    <RANKING order="2" place="2" resultid="4173" />
                    <RANKING order="3" place="3" resultid="3080" />
                    <RANKING order="4" place="4" resultid="2473" />
                    <RANKING order="5" place="5" resultid="4978" />
                    <RANKING order="6" place="6" resultid="4280" />
                    <RANKING order="7" place="7" resultid="3174" />
                    <RANKING order="8" place="-1" resultid="5040" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1486" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3014" />
                    <RANKING order="2" place="2" resultid="5176" />
                    <RANKING order="3" place="3" resultid="2152" />
                    <RANKING order="4" place="4" resultid="1918" />
                    <RANKING order="5" place="5" resultid="2459" />
                    <RANKING order="6" place="6" resultid="2492" />
                    <RANKING order="7" place="-1" resultid="4678" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1487" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4180" />
                    <RANKING order="2" place="2" resultid="3966" />
                    <RANKING order="3" place="3" resultid="4102" />
                    <RANKING order="4" place="4" resultid="4638" />
                    <RANKING order="5" place="5" resultid="2394" />
                    <RANKING order="6" place="-1" resultid="3181" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1488" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2855" />
                    <RANKING order="2" place="2" resultid="2503" />
                    <RANKING order="3" place="3" resultid="5152" />
                    <RANKING order="4" place="4" resultid="3166" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1489" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2876" />
                    <RANKING order="2" place="2" resultid="2027" />
                    <RANKING order="3" place="3" resultid="2863" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1490" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4844" />
                    <RANKING order="2" place="2" resultid="4088" />
                    <RANKING order="3" place="3" resultid="4094" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1491" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4868" />
                    <RANKING order="2" place="2" resultid="2608" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1492" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1493" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3158" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1494" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1495" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7024" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7025" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7026" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7027" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7028" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7029" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7030" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7031" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1496" daytime="17:25" gender="M" number="26" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1497" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4234" />
                    <RANKING order="2" place="2" resultid="2070" />
                    <RANKING order="3" place="3" resultid="3841" />
                    <RANKING order="4" place="4" resultid="5098" />
                    <RANKING order="5" place="5" resultid="2092" />
                    <RANKING order="6" place="6" resultid="5019" />
                    <RANKING order="7" place="-1" resultid="5452" />
                    <RANKING order="8" place="-1" resultid="5454" />
                    <RANKING order="9" place="-1" resultid="2085" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1498" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2952" />
                    <RANKING order="2" place="2" resultid="2934" />
                    <RANKING order="3" place="3" resultid="2742" />
                    <RANKING order="4" place="4" resultid="5126" />
                    <RANKING order="5" place="5" resultid="3246" />
                    <RANKING order="6" place="6" resultid="1884" />
                    <RANKING order="7" place="7" resultid="2426" />
                    <RANKING order="8" place="8" resultid="4130" />
                    <RANKING order="9" place="-1" resultid="2941" />
                    <RANKING order="10" place="-1" resultid="3599" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1499" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2545" />
                    <RANKING order="2" place="2" resultid="3304" />
                    <RANKING order="3" place="3" resultid="4765" />
                    <RANKING order="4" place="4" resultid="5107" />
                    <RANKING order="5" place="5" resultid="4564" />
                    <RANKING order="6" place="6" resultid="4321" />
                    <RANKING order="7" place="7" resultid="4342" />
                    <RANKING order="8" place="8" resultid="3674" />
                    <RANKING order="9" place="9" resultid="4332" />
                    <RANKING order="10" place="-1" resultid="3022" />
                    <RANKING order="11" place="-1" resultid="3638" />
                    <RANKING order="12" place="-1" resultid="3652" />
                    <RANKING order="13" place="-1" resultid="4796" />
                    <RANKING order="14" place="-1" resultid="6703" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1500" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3420" />
                    <RANKING order="2" place="2" resultid="3073" />
                    <RANKING order="3" place="3" resultid="5279" />
                    <RANKING order="4" place="4" resultid="2224" />
                    <RANKING order="5" place="5" resultid="4373" />
                    <RANKING order="6" place="6" resultid="4422" />
                    <RANKING order="7" place="7" resultid="2311" />
                    <RANKING order="8" place="-1" resultid="2682" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1501" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2182" />
                    <RANKING order="2" place="2" resultid="4485" />
                    <RANKING order="3" place="3" resultid="2307" />
                    <RANKING order="4" place="4" resultid="5457" />
                    <RANKING order="5" place="5" resultid="3461" />
                    <RANKING order="6" place="6" resultid="5337" />
                    <RANKING order="7" place="7" resultid="5263" />
                    <RANKING order="8" place="8" resultid="4301" />
                    <RANKING order="9" place="-1" resultid="3231" />
                    <RANKING order="10" place="-1" resultid="4550" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1502" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3264" />
                    <RANKING order="2" place="2" resultid="4850" />
                    <RANKING order="3" place="3" resultid="2564" />
                    <RANKING order="4" place="4" resultid="1891" />
                    <RANKING order="5" place="5" resultid="2197" />
                    <RANKING order="6" place="6" resultid="4662" />
                    <RANKING order="7" place="7" resultid="5404" />
                    <RANKING order="8" place="8" resultid="2632" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1503" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2708" />
                    <RANKING order="2" place="2" resultid="3038" />
                    <RANKING order="3" place="3" resultid="2479" />
                    <RANKING order="4" place="4" resultid="4079" />
                    <RANKING order="5" place="5" resultid="5242" />
                    <RANKING order="6" place="6" resultid="3396" />
                    <RANKING order="7" place="7" resultid="3732" />
                    <RANKING order="8" place="8" resultid="4241" />
                    <RANKING order="9" place="-1" resultid="4207" />
                    <RANKING order="10" place="-1" resultid="4891" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1504" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4900" />
                    <RANKING order="2" place="2" resultid="4618" />
                    <RANKING order="3" place="3" resultid="4884" />
                    <RANKING order="4" place="4" resultid="2827" />
                    <RANKING order="5" place="5" resultid="3008" />
                    <RANKING order="6" place="6" resultid="2776" />
                    <RANKING order="7" place="7" resultid="3755" />
                    <RANKING order="8" place="8" resultid="4772" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1505" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4294" />
                    <RANKING order="2" place="2" resultid="4007" />
                    <RANKING order="3" place="3" resultid="5235" />
                    <RANKING order="4" place="4" resultid="2832" />
                    <RANKING order="5" place="5" resultid="6211" />
                    <RANKING order="6" place="6" resultid="2884" />
                    <RANKING order="7" place="7" resultid="2585" />
                    <RANKING order="8" place="-1" resultid="2890" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1506" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2869" />
                    <RANKING order="2" place="2" resultid="5222" />
                    <RANKING order="3" place="3" resultid="5213" />
                    <RANKING order="4" place="4" resultid="5210" />
                    <RANKING order="5" place="5" resultid="3620" />
                    <RANKING order="6" place="-1" resultid="2647" />
                    <RANKING order="7" place="-1" resultid="3993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1507" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2370" />
                    <RANKING order="2" place="2" resultid="5201" />
                    <RANKING order="3" place="3" resultid="5205" />
                    <RANKING order="4" place="4" resultid="3606" />
                    <RANKING order="5" place="5" resultid="4708" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1508" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4110" />
                    <RANKING order="2" place="2" resultid="5197" />
                    <RANKING order="3" place="3" resultid="1981" />
                    <RANKING order="4" place="4" resultid="4157" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1509" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2447" />
                    <RANKING order="2" place="2" resultid="2323" />
                    <RANKING order="3" place="3" resultid="4910" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1510" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1511" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1512" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7032" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7033" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7034" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7035" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7036" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7037" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7038" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7039" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7040" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7041" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7042" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7043" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1513" daytime="17:42" gender="F" number="27" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1643" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3919" />
                    <RANKING order="2" place="2" resultid="5015" />
                    <RANKING order="3" place="3" resultid="3929" />
                    <RANKING order="4" place="4" resultid="3927" />
                    <RANKING order="5" place="5" resultid="5423" />
                    <RANKING order="6" place="6" resultid="3931" />
                    <RANKING order="7" place="7" resultid="7266" />
                    <RANKING order="8" place="8" resultid="5421" />
                    <RANKING order="9" place="-1" resultid="5443" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7044" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1530" daytime="17:45" gender="M" number="28" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1644" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3921" />
                    <RANKING order="2" place="2" resultid="5020" />
                    <RANKING order="3" place="3" resultid="4975" />
                    <RANKING order="4" place="4" resultid="3925" />
                    <RANKING order="5" place="5" resultid="5448" />
                    <RANKING order="6" place="6" resultid="5449" />
                    <RANKING order="7" place="6" resultid="3923" />
                    <RANKING order="8" place="8" resultid="2376" />
                    <RANKING order="9" place="9" resultid="5453" />
                    <RANKING order="10" place="10" resultid="5419" />
                    <RANKING order="11" place="11" resultid="5407" />
                    <RANKING order="12" place="12" resultid="5409" />
                    <RANKING order="13" place="-1" resultid="5451" />
                    <RANKING order="14" place="-1" resultid="5415" />
                    <RANKING order="15" place="-1" resultid="5441" />
                    <RANKING order="16" place="-1" resultid="3344" />
                    <RANKING order="17" place="-1" resultid="5413" />
                    <RANKING order="18" place="-1" resultid="5417" />
                    <RANKING order="19" place="-1" resultid="5411" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7045" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7046" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7047" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1547" daytime="17:49" gender="F" number="29" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1548" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3333" />
                    <RANKING order="2" place="2" resultid="2420" />
                    <RANKING order="3" place="3" resultid="3660" />
                    <RANKING order="4" place="4" resultid="3980" />
                    <RANKING order="5" place="5" resultid="3271" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1549" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4632" />
                    <RANKING order="2" place="2" resultid="2923" />
                    <RANKING order="3" place="3" resultid="3225" />
                    <RANKING order="4" place="4" resultid="3121" />
                    <RANKING order="5" place="5" resultid="4266" />
                    <RANKING order="6" place="6" resultid="4398" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1550" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3055" />
                    <RANKING order="2" place="2" resultid="4833" />
                    <RANKING order="3" place="3" resultid="2641" />
                    <RANKING order="4" place="-1" resultid="2762" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1551" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2839" />
                    <RANKING order="2" place="2" resultid="2688" />
                    <RANKING order="3" place="3" resultid="2784" />
                    <RANKING order="4" place="4" resultid="2134" />
                    <RANKING order="5" place="-1" resultid="5285" />
                    <RANKING order="6" place="-1" resultid="5374" />
                    <RANKING order="7" place="-1" resultid="3986" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1552" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3825" />
                    <RANKING order="2" place="2" resultid="4731" />
                    <RANKING order="3" place="-1" resultid="4653" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1553" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3321" />
                    <RANKING order="2" place="2" resultid="2110" />
                    <RANKING order="3" place="3" resultid="2160" />
                    <RANKING order="4" place="4" resultid="2474" />
                    <RANKING order="5" place="5" resultid="5041" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1554" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3015" />
                    <RANKING order="2" place="2" resultid="3067" />
                    <RANKING order="3" place="3" resultid="3412" />
                    <RANKING order="4" place="4" resultid="2493" />
                    <RANKING order="5" place="-1" resultid="4679" />
                    <RANKING order="6" place="-1" resultid="1942" />
                    <RANKING order="7" place="-1" resultid="1935" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1555" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4273" />
                    <RANKING order="2" place="2" resultid="2395" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1556" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5157" />
                    <RANKING order="2" place="2" resultid="2657" />
                    <RANKING order="3" place="3" resultid="2676" />
                    <RANKING order="4" place="4" resultid="3214" />
                    <RANKING order="5" place="-1" resultid="2504" />
                    <RANKING order="6" place="-1" resultid="2820" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1557" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2451" />
                    <RANKING order="2" place="2" resultid="4964" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1558" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4095" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1559" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1560" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3106" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1561" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1562" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1563" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7048" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7049" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7050" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7051" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7052" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7053" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1564" daytime="18:14" gender="M" number="30" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1565" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2441" />
                    <RANKING order="2" place="2" resultid="4918" />
                    <RANKING order="3" place="3" resultid="2078" />
                    <RANKING order="4" place="4" resultid="3811" />
                    <RANKING order="5" place="-1" resultid="2086" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1566" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4415" />
                    <RANKING order="2" place="2" resultid="3770" />
                    <RANKING order="3" place="3" resultid="4858" />
                    <RANKING order="4" place="4" resultid="2935" />
                    <RANKING order="5" place="5" resultid="2331" />
                    <RANKING order="6" place="6" resultid="2771" />
                    <RANKING order="7" place="7" resultid="4131" />
                    <RANKING order="8" place="8" resultid="4759" />
                    <RANKING order="9" place="9" resultid="4492" />
                    <RANKING order="10" place="-1" resultid="2743" />
                    <RANKING order="11" place="-1" resultid="3875" />
                    <RANKING order="12" place="-1" resultid="5136" />
                    <RANKING order="13" place="-1" resultid="4499" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1567" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2590" />
                    <RANKING order="2" place="2" resultid="3653" />
                    <RANKING order="3" place="3" resultid="3023" />
                    <RANKING order="4" place="4" resultid="5061" />
                    <RANKING order="5" place="5" resultid="4366" />
                    <RANKING order="6" place="6" resultid="3645" />
                    <RANKING order="7" place="7" resultid="2540" />
                    <RANKING order="8" place="8" resultid="5077" />
                    <RANKING order="9" place="9" resultid="4073" />
                    <RANKING order="10" place="-1" resultid="3748" />
                    <RANKING order="11" place="-1" resultid="4337" />
                    <RANKING order="12" place="-1" resultid="4363" />
                    <RANKING order="13" place="-1" resultid="5402" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1568" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3429" />
                    <RANKING order="2" place="2" resultid="3350" />
                    <RANKING order="3" place="3" resultid="3330" />
                    <RANKING order="4" place="4" resultid="3483" />
                    <RANKING order="5" place="5" resultid="3903" />
                    <RANKING order="6" place="6" resultid="3241" />
                    <RANKING order="7" place="7" resultid="4558" />
                    <RANKING order="8" place="8" resultid="5344" />
                    <RANKING order="9" place="9" resultid="1960" />
                    <RANKING order="10" place="-1" resultid="3853" />
                    <RANKING order="11" place="-1" resultid="3728" />
                    <RANKING order="12" place="-1" resultid="4374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1569" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2514" />
                    <RANKING order="2" place="2" resultid="5366" />
                    <RANKING order="3" place="3" resultid="3359" />
                    <RANKING order="4" place="4" resultid="3522" />
                    <RANKING order="5" place="5" resultid="4042" />
                    <RANKING order="6" place="6" resultid="3294" />
                    <RANKING order="7" place="7" resultid="4036" />
                    <RANKING order="8" place="8" resultid="2702" />
                    <RANKING order="9" place="9" resultid="4302" />
                    <RANKING order="10" place="10" resultid="3505" />
                    <RANKING order="11" place="11" resultid="2580" />
                    <RANKING order="12" place="12" resultid="2189" />
                    <RANKING order="13" place="13" resultid="4723" />
                    <RANKING order="14" place="14" resultid="4143" />
                    <RANKING order="15" place="15" resultid="3232" />
                    <RANKING order="16" place="16" resultid="2212" />
                    <RANKING order="17" place="-1" resultid="2619" />
                    <RANKING order="18" place="-1" resultid="4052" />
                    <RANKING order="19" place="-1" resultid="3114" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1570" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3288" />
                    <RANKING order="2" place="2" resultid="5047" />
                    <RANKING order="3" place="3" resultid="4851" />
                    <RANKING order="4" place="4" resultid="4543" />
                    <RANKING order="5" place="5" resultid="5258" />
                    <RANKING order="6" place="6" resultid="2520" />
                    <RANKING order="7" place="7" resultid="5033" />
                    <RANKING order="8" place="8" resultid="5090" />
                    <RANKING order="9" place="-1" resultid="3703" />
                    <RANKING order="10" place="-1" resultid="2596" />
                    <RANKING order="11" place="-1" resultid="3938" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1571" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3468" />
                    <RANKING order="2" place="2" resultid="4029" />
                    <RANKING order="3" place="3" resultid="3000" />
                    <RANKING order="4" place="4" resultid="3566" />
                    <RANKING order="5" place="5" resultid="5359" />
                    <RANKING order="6" place="6" resultid="2603" />
                    <RANKING order="7" place="7" resultid="5399" />
                    <RANKING order="8" place="-1" resultid="2558" />
                    <RANKING order="9" place="-1" resultid="3039" />
                    <RANKING order="10" place="-1" resultid="3897" />
                    <RANKING order="11" place="-1" resultid="4892" />
                    <RANKING order="12" place="-1" resultid="4946" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1572" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4901" />
                    <RANKING order="2" place="2" resultid="3586" />
                    <RANKING order="3" place="3" resultid="2355" />
                    <RANKING order="4" place="4" resultid="2828" />
                    <RANKING order="5" place="5" resultid="4068" />
                    <RANKING order="6" place="6" resultid="2010" />
                    <RANKING order="7" place="7" resultid="4927" />
                    <RANKING order="8" place="8" resultid="3389" />
                    <RANKING order="9" place="9" resultid="4773" />
                    <RANKING order="10" place="-1" resultid="5382" />
                    <RANKING order="11" place="-1" resultid="3405" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1573" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4008" />
                    <RANKING order="2" place="2" resultid="2363" />
                    <RANKING order="3" place="3" resultid="3719" />
                    <RANKING order="4" place="4" resultid="4702" />
                    <RANKING order="5" place="5" resultid="3615" />
                    <RANKING order="6" place="-1" resultid="3834" />
                    <RANKING order="7" place="-1" resultid="5120" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1574" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2870" />
                    <RANKING order="2" place="2" resultid="2648" />
                    <RANKING order="3" place="3" resultid="2455" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1575" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4000" />
                    <RANKING order="2" place="2" resultid="2371" />
                    <RANKING order="3" place="3" resultid="3607" />
                    <RANKING order="4" place="4" resultid="4119" />
                    <RANKING order="5" place="5" resultid="3128" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1576" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4111" />
                    <RANKING order="2" place="2" resultid="4158" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1577" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2324" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1578" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4200" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1579" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1580" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7054" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7055" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7056" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7057" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7058" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7059" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7060" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7061" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7062" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7063" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7064" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7065" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7066" number="13" order="13" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1581" daytime="18:59" gender="F" number="31" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1582" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2057" />
                    <RANKING order="2" place="2" resultid="3661" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1583" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2727" />
                    <RANKING order="2" place="2" resultid="2663" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1584" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2763" />
                    <RANKING order="2" place="2" resultid="3974" />
                    <RANKING order="3" place="-1" resultid="2573" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1585" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2168" />
                    <RANKING order="2" place="2" resultid="1857" />
                    <RANKING order="3" place="3" resultid="1948" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1586" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3573" />
                    <RANKING order="2" place="2" resultid="3498" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1587" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2993" />
                    <RANKING order="2" place="2" resultid="3081" />
                    <RANKING order="3" place="3" resultid="4166" />
                    <RANKING order="4" place="4" resultid="4979" />
                    <RANKING order="5" place="5" resultid="3278" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1588" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2128" />
                    <RANKING order="2" place="2" resultid="1976" />
                    <RANKING order="3" place="3" resultid="1919" />
                    <RANKING order="4" place="4" resultid="3581" />
                    <RANKING order="5" place="5" resultid="2507" />
                    <RANKING order="6" place="-1" resultid="4518" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1589" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4181" />
                    <RANKING order="2" place="2" resultid="3967" />
                    <RANKING order="3" place="3" resultid="4103" />
                    <RANKING order="4" place="4" resultid="1995" />
                    <RANKING order="5" place="-1" resultid="5164" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1590" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="2856" />
                    <RANKING order="2" place="-1" resultid="4952" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1591" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="4959" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1592" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1593" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1594" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1595" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1596" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1597" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7067" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7068" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7069" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7070" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1598" daytime="19:19" gender="M" number="32" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1599" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3774" />
                    <RANKING order="2" place="2" resultid="2093" />
                    <RANKING order="3" place="3" resultid="1864" />
                    <RANKING order="4" place="4" resultid="1871" />
                    <RANKING order="5" place="-1" resultid="3817" />
                    <RANKING order="6" place="-1" resultid="5099" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1600" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2332" />
                    <RANKING order="2" place="2" resultid="2906" />
                    <RANKING order="3" place="3" resultid="2953" />
                    <RANKING order="4" place="4" resultid="4214" />
                    <RANKING order="5" place="5" resultid="2946" />
                    <RANKING order="6" place="-1" resultid="4760" />
                    <RANKING order="7" place="-1" resultid="5054" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1601" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2591" />
                    <RANKING order="2" place="2" resultid="4380" />
                    <RANKING order="3" place="3" resultid="4314" />
                    <RANKING order="4" place="4" resultid="5069" />
                    <RANKING order="5" place="5" resultid="3675" />
                    <RANKING order="6" place="6" resultid="3491" />
                    <RANKING order="7" place="7" resultid="3445" />
                    <RANKING order="8" place="-1" resultid="4645" />
                    <RANKING order="9" place="-1" resultid="2749" />
                    <RANKING order="10" place="-1" resultid="4349" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1602" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3514" />
                    <RANKING order="2" place="2" resultid="3351" />
                    <RANKING order="3" place="3" resultid="3421" />
                    <RANKING order="4" place="4" resultid="2225" />
                    <RANKING order="5" place="-1" resultid="2312" />
                    <RANKING order="6" place="-1" resultid="3437" />
                    <RANKING order="7" place="-1" resultid="4671" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1603" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5367" />
                    <RANKING order="2" place="2" resultid="3506" />
                    <RANKING order="3" place="3" resultid="4724" />
                    <RANKING order="4" place="4" resultid="3863" />
                    <RANKING order="5" place="5" resultid="2235" />
                    <RANKING order="6" place="-1" resultid="4017" />
                    <RANKING order="7" place="-1" resultid="2515" />
                    <RANKING order="8" place="-1" resultid="3031" />
                    <RANKING order="9" place="-1" resultid="5264" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1604" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3265" />
                    <RANKING order="2" place="2" resultid="3088" />
                    <RANKING order="3" place="3" resultid="4716" />
                    <RANKING order="4" place="4" resultid="4221" />
                    <RANKING order="5" place="-1" resultid="2218" />
                    <RANKING order="6" place="-1" resultid="2565" />
                    <RANKING order="7" place="-1" resultid="3311" />
                    <RANKING order="8" place="-1" resultid="5091" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1605" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3469" />
                    <RANKING order="2" place="2" resultid="3099" />
                    <RANKING order="3" place="3" resultid="3914" />
                    <RANKING order="4" place="4" resultid="3712" />
                    <RANKING order="5" place="5" resultid="5394" />
                    <RANKING order="6" place="6" resultid="3397" />
                    <RANKING order="7" place="-1" resultid="2709" />
                    <RANKING order="8" place="-1" resultid="4826" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1606" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4619" />
                    <RANKING order="2" place="2" resultid="5238" />
                    <RANKING order="3" place="3" resultid="4940" />
                    <RANKING order="4" place="4" resultid="2812" />
                    <RANKING order="5" place="5" resultid="4189" />
                    <RANKING order="6" place="6" resultid="3633" />
                    <RANKING order="7" place="7" resultid="4885" />
                    <RANKING order="8" place="8" resultid="4781" />
                    <RANKING order="9" place="9" resultid="3756" />
                    <RANKING order="10" place="10" resultid="3153" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1607" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3453" />
                    <RANKING order="2" place="2" resultid="5229" />
                    <RANKING order="3" place="3" resultid="4431" />
                    <RANKING order="4" place="4" resultid="2467" />
                    <RANKING order="5" place="5" resultid="4971" />
                    <RANKING order="6" place="6" resultid="2411" />
                    <RANKING order="7" place="7" resultid="3380" />
                    <RANKING order="8" place="8" resultid="3145" />
                    <RANKING order="9" place="-1" resultid="2377" />
                    <RANKING order="10" place="-1" resultid="4295" />
                    <RANKING order="11" place="-1" resultid="5430" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1608" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4060" />
                    <RANKING order="2" place="2" resultid="5352" />
                    <RANKING order="3" place="-1" resultid="5223" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1609" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1927" />
                    <RANKING order="2" place="2" resultid="4694" />
                    <RANKING order="3" place="3" resultid="2533" />
                    <RANKING order="4" place="-1" resultid="3129" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1610" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1611" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4612" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1612" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1613" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1614" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7071" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7072" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7073" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7074" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7075" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7076" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7077" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7078" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7079" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7080" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1615" daytime="19:57" gender="X" number="33" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1632" agemax="96" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="2097" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1633" agemax="119" agemin="100">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2975" />
                    <RANKING order="2" place="2" resultid="2789" />
                    <RANKING order="3" place="3" resultid="4408" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1634" agemax="159" agemin="120">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4876" />
                    <RANKING order="2" place="2" resultid="7268" />
                    <RANKING order="3" place="3" resultid="2243" />
                    <RANKING order="4" place="-1" resultid="4744" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1635" agemax="199" agemin="160">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2251" />
                    <RANKING order="2" place="2" resultid="5296" />
                    <RANKING order="3" place="3" resultid="2787" />
                    <RANKING order="4" place="-1" resultid="7269" />
                    <RANKING order="5" place="-1" resultid="4305" />
                    <RANKING order="6" place="-1" resultid="5424" />
                    <RANKING order="7" place="-1" resultid="7270" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1636" agemax="239" agemin="200">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2253" />
                    <RANKING order="2" place="2" resultid="5298" />
                    <RANKING order="3" place="3" resultid="3184" />
                    <RANKING order="4" place="-1" resultid="3044" />
                    <RANKING order="5" place="-1" resultid="4986" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1637" agemax="279" agemin="240">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2900" />
                    <RANKING order="2" place="-1" resultid="5300" />
                    <RANKING order="3" place="-1" resultid="4985" />
                    <RANKING order="4" place="-1" resultid="7271" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1638" agemax="319" agemin="280">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7267" />
                    <RANKING order="2" place="2" resultid="3190" />
                    <RANKING order="3" place="-1" resultid="6664" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1639" agemax="359" agemin="320" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7440" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7441" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7442" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7443" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2011-11-20" daytime="09:30" number="4">
          <EVENTS>
            <EVENT eventid="1641" daytime="09:30" gender="F" number="34" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1647" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4873" />
                    <RANKING order="2" place="2" resultid="2058" />
                    <RANKING order="3" place="3" resultid="2063" />
                    <RANKING order="4" place="4" resultid="3662" />
                    <RANKING order="5" place="-1" resultid="5013" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1648" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1878" />
                    <RANKING order="2" place="2" resultid="3890" />
                    <RANKING order="3" place="3" resultid="2958" />
                    <RANKING order="4" place="4" resultid="2728" />
                    <RANKING order="5" place="5" resultid="1969" />
                    <RANKING order="6" place="6" resultid="2664" />
                    <RANKING order="7" place="7" resultid="3122" />
                    <RANKING order="8" place="8" resultid="2963" />
                    <RANKING order="9" place="-1" resultid="2924" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1649" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4810" />
                    <RANKING order="2" place="2" resultid="3056" />
                    <RANKING order="3" place="3" resultid="4834" />
                    <RANKING order="4" place="4" resultid="3669" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1650" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2303" />
                    <RANKING order="2" place="2" resultid="5286" />
                    <RANKING order="3" place="-1" resultid="2135" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1651" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3574" />
                    <RANKING order="2" place="2" resultid="3499" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1652" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2994" />
                    <RANKING order="2" place="2" resultid="2161" />
                    <RANKING order="3" place="3" resultid="3082" />
                    <RANKING order="4" place="4" resultid="4174" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1653" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3016" />
                    <RANKING order="2" place="2" resultid="1977" />
                    <RANKING order="3" place="3" resultid="4680" />
                    <RANKING order="4" place="4" resultid="2129" />
                    <RANKING order="5" place="5" resultid="3413" />
                    <RANKING order="6" place="6" resultid="1920" />
                    <RANKING order="7" place="7" resultid="3582" />
                    <RANKING order="8" place="8" resultid="2508" />
                    <RANKING order="9" place="-1" resultid="2460" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1654" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4182" />
                    <RANKING order="2" place="2" resultid="2019" />
                    <RANKING order="3" place="3" resultid="5165" />
                    <RANKING order="4" place="4" resultid="2396" />
                    <RANKING order="5" place="5" resultid="1996" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1655" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3958" />
                    <RANKING order="2" place="2" resultid="2821" />
                    <RANKING order="3" place="3" resultid="3167" />
                    <RANKING order="4" place="-1" resultid="4953" />
                    <RANKING order="5" place="-1" resultid="5158" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1656" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2850" />
                    <RANKING order="2" place="2" resultid="1988" />
                    <RANKING order="3" place="-1" resultid="2877" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1657" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1658" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1659" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1660" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1661" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1662" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7275" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7276" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7277" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7278" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7279" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7280" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1645" daytime="09:38" gender="M" number="35" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1663" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3792" />
                    <RANKING order="2" place="2" resultid="4235" />
                    <RANKING order="3" place="3" resultid="1894" />
                    <RANKING order="4" place="4" resultid="2442" />
                    <RANKING order="5" place="5" resultid="3782" />
                    <RANKING order="6" place="6" resultid="2079" />
                    <RANKING order="7" place="7" resultid="2071" />
                    <RANKING order="8" place="8" resultid="1865" />
                    <RANKING order="9" place="9" resultid="3906" />
                    <RANKING order="10" place="-1" resultid="3818" />
                    <RANKING order="11" place="-1" resultid="5021" />
                    <RANKING order="12" place="-1" resultid="4919" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1664" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4416" />
                    <RANKING order="2" place="2" resultid="3600" />
                    <RANKING order="3" place="3" resultid="4859" />
                    <RANKING order="4" place="4" resultid="1885" />
                    <RANKING order="5" place="5" resultid="2936" />
                    <RANKING order="6" place="6" resultid="5112" />
                    <RANKING order="7" place="7" resultid="4215" />
                    <RANKING order="8" place="8" resultid="2929" />
                    <RANKING order="9" place="9" resultid="5127" />
                    <RANKING order="10" place="10" resultid="5055" />
                    <RANKING order="11" place="11" resultid="2947" />
                    <RANKING order="12" place="12" resultid="3208" />
                    <RANKING order="13" place="13" resultid="3869" />
                    <RANKING order="14" place="14" resultid="4132" />
                    <RANKING order="15" place="-1" resultid="2942" />
                    <RANKING order="16" place="-1" resultid="3247" />
                    <RANKING order="17" place="-1" resultid="4761" />
                    <RANKING order="18" place="-1" resultid="3876" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1665" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2546" />
                    <RANKING order="2" place="2" resultid="3305" />
                    <RANKING order="3" place="3" resultid="5145" />
                    <RANKING order="4" place="4" resultid="4354" />
                    <RANKING order="5" place="5" resultid="5062" />
                    <RANKING order="6" place="6" resultid="3024" />
                    <RANKING order="7" place="7" resultid="2750" />
                    <RANKING order="8" place="8" resultid="3676" />
                    <RANKING order="9" place="9" resultid="4367" />
                    <RANKING order="10" place="10" resultid="4565" />
                    <RANKING order="11" place="11" resultid="4333" />
                    <RANKING order="12" place="12" resultid="4338" />
                    <RANKING order="13" place="13" resultid="4315" />
                    <RANKING order="14" place="14" resultid="3646" />
                    <RANKING order="15" place="15" resultid="2720" />
                    <RANKING order="16" place="16" resultid="3749" />
                    <RANKING order="17" place="-1" resultid="4074" />
                    <RANKING order="18" place="-1" resultid="4381" />
                    <RANKING order="19" place="-1" resultid="5108" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1666" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3430" />
                    <RANKING order="2" place="2" resultid="5280" />
                    <RANKING order="3" place="3" resultid="3074" />
                    <RANKING order="4" place="4" resultid="2226" />
                    <RANKING order="5" place="5" resultid="4423" />
                    <RANKING order="6" place="6" resultid="3484" />
                    <RANKING order="7" place="7" resultid="2204" />
                    <RANKING order="8" place="8" resultid="2313" />
                    <RANKING order="9" place="9" resultid="1961" />
                    <RANKING order="10" place="10" resultid="4559" />
                    <RANKING order="11" place="11" resultid="5345" />
                    <RANKING order="12" place="12" resultid="4672" />
                    <RANKING order="13" place="-1" resultid="3242" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1667" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2620" />
                    <RANKING order="2" place="2" resultid="3220" />
                    <RANKING order="3" place="3" resultid="2174" />
                    <RANKING order="4" place="4" resultid="3360" />
                    <RANKING order="5" place="5" resultid="5338" />
                    <RANKING order="6" place="6" resultid="4303" />
                    <RANKING order="7" place="7" resultid="4023" />
                    <RANKING order="8" place="8" resultid="3462" />
                    <RANKING order="9" place="9" resultid="2190" />
                    <RANKING order="10" place="10" resultid="4018" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1668" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3266" />
                    <RANKING order="2" place="2" resultid="3289" />
                    <RANKING order="3" place="3" resultid="3089" />
                    <RANKING order="4" place="4" resultid="2198" />
                    <RANKING order="5" place="5" resultid="4538" />
                    <RANKING order="6" place="6" resultid="4717" />
                    <RANKING order="7" place="7" resultid="5034" />
                    <RANKING order="8" place="-1" resultid="3704" />
                    <RANKING order="9" place="-1" resultid="3939" />
                    <RANKING order="10" place="-1" resultid="4222" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1669" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2710" />
                    <RANKING order="2" place="2" resultid="3040" />
                    <RANKING order="3" place="3" resultid="4208" />
                    <RANKING order="4" place="4" resultid="3713" />
                    <RANKING order="5" place="5" resultid="4247" />
                    <RANKING order="6" place="6" resultid="3001" />
                    <RANKING order="7" place="7" resultid="2604" />
                    <RANKING order="8" place="8" resultid="3733" />
                    <RANKING order="9" place="9" resultid="5360" />
                    <RANKING order="10" place="-1" resultid="4030" />
                    <RANKING order="11" place="-1" resultid="3898" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1670" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3587" />
                    <RANKING order="2" place="2" resultid="4820" />
                    <RANKING order="3" place="3" resultid="3634" />
                    <RANKING order="4" place="4" resultid="2356" />
                    <RANKING order="5" place="5" resultid="2340" />
                    <RANKING order="6" place="6" resultid="3682" />
                    <RANKING order="7" place="7" resultid="2777" />
                    <RANKING order="8" place="8" resultid="3757" />
                    <RANKING order="9" place="9" resultid="3154" />
                    <RANKING order="10" place="-1" resultid="3062" />
                    <RANKING order="11" place="-1" resultid="2813" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1671" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4296" />
                    <RANKING order="2" place="2" resultid="2891" />
                    <RANKING order="3" place="3" resultid="5251" />
                    <RANKING order="4" place="4" resultid="2586" />
                    <RANKING order="5" place="5" resultid="2716" />
                    <RANKING order="6" place="6" resultid="2885" />
                    <RANKING order="7" place="7" resultid="2378" />
                    <RANKING order="8" place="8" resultid="3381" />
                    <RANKING order="9" place="9" resultid="2412" />
                    <RANKING order="10" place="10" resultid="3146" />
                    <RANKING order="11" place="-1" resultid="5431" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1672" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4061" />
                    <RANKING order="2" place="2" resultid="2349" />
                    <RANKING order="3" place="-1" resultid="3994" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1673" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2498" />
                    <RANKING order="2" place="2" resultid="3135" />
                    <RANKING order="3" place="3" resultid="4001" />
                    <RANKING order="4" place="-1" resultid="4120" />
                    <RANKING order="5" place="-1" resultid="4125" />
                    <RANKING order="6" place="-1" resultid="5202" />
                    <RANKING order="7" place="-1" resultid="5206" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1674" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1675" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1676" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1677" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1678" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7281" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7282" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7283" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7284" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7285" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7286" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7287" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7288" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7289" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7290" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7291" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7292" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7293" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7294" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1679" daytime="09:56" gender="F" number="36" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1680" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="5014" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1681" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2122" />
                    <RANKING order="2" place="2" resultid="2665" />
                    <RANKING order="3" place="3" resultid="4267" />
                    <RANKING order="4" place="4" resultid="4399" />
                    <RANKING order="5" place="5" resultid="4392" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1682" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2756" />
                    <RANKING order="2" place="2" resultid="3670" />
                    <RANKING order="3" place="3" resultid="2574" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1683" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2840" />
                    <RANKING order="2" place="2" resultid="2626" />
                    <RANKING order="3" place="3" resultid="5189" />
                    <RANKING order="4" place="4" resultid="5375" />
                    <RANKING order="5" place="5" resultid="1949" />
                    <RANKING order="6" place="6" resultid="2785" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1684" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3575" />
                    <RANKING order="2" place="2" resultid="3500" />
                    <RANKING order="3" place="3" resultid="3826" />
                    <RANKING order="4" place="4" resultid="4732" />
                    <RANKING order="5" place="-1" resultid="4654" />
                    <RANKING order="6" place="-1" resultid="2145" />
                    <RANKING order="7" place="-1" resultid="4593" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1685" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2614" />
                    <RANKING order="2" place="2" resultid="4167" />
                    <RANKING order="3" place="3" resultid="4281" />
                    <RANKING order="4" place="4" resultid="3175" />
                    <RANKING order="5" place="5" resultid="4933" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1686" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2153" />
                    <RANKING order="2" place="2" resultid="2003" />
                    <RANKING order="3" place="3" resultid="1955" />
                    <RANKING order="4" place="4" resultid="3299" />
                    <RANKING order="5" place="5" resultid="2139" />
                    <RANKING order="6" place="6" resultid="1943" />
                    <RANKING order="7" place="-1" resultid="4083" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1687" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2020" />
                    <RANKING order="2" place="2" resultid="3968" />
                    <RANKING order="3" place="3" resultid="4104" />
                    <RANKING order="4" place="-1" resultid="3182" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1688" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2881" />
                    <RANKING order="2" place="2" resultid="2488" />
                    <RANKING order="3" place="3" resultid="2117" />
                    <RANKING order="4" place="4" resultid="3215" />
                    <RANKING order="5" place="-1" resultid="5153" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1689" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2864" />
                    <RANKING order="2" place="2" resultid="2851" />
                    <RANKING order="3" place="3" resultid="1989" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1690" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1691" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3326" />
                    <RANKING order="2" place="2" resultid="4863" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1692" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3107" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1693" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2024" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1694" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1695" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7295" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7296" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7297" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7298" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7299" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7300" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1696" daytime="10:14" gender="M" number="37" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1697" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3842" />
                    <RANKING order="2" place="2" resultid="2968" />
                    <RANKING order="3" place="3" resultid="3788" />
                    <RANKING order="4" place="4" resultid="3819" />
                    <RANKING order="5" place="5" resultid="1872" />
                    <RANKING order="6" place="6" resultid="4906" />
                    <RANKING order="7" place="-1" resultid="2087" />
                    <RANKING order="8" place="-1" resultid="5442" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1698" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2907" />
                    <RANKING order="2" place="2" resultid="2670" />
                    <RANKING order="3" place="3" resultid="2913" />
                    <RANKING order="4" place="4" resultid="4500" />
                    <RANKING order="5" place="5" resultid="2436" />
                    <RANKING order="6" place="-1" resultid="5447" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1699" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5140" />
                    <RANKING order="2" place="2" resultid="4350" />
                    <RANKING order="3" place="3" resultid="3446" />
                    <RANKING order="4" place="4" resultid="4646" />
                    <RANKING order="5" place="5" resultid="4322" />
                    <RANKING order="6" place="6" resultid="3492" />
                    <RANKING order="7" place="7" resultid="4328" />
                    <RANKING order="8" place="-1" resultid="4150" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1700" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3515" />
                    <RANKING order="2" place="2" resultid="3485" />
                    <RANKING order="3" place="3" resultid="3438" />
                    <RANKING order="4" place="4" resultid="2241" />
                    <RANKING order="5" place="5" resultid="2317" />
                    <RANKING order="6" place="-1" resultid="3854" />
                    <RANKING order="7" place="-1" resultid="3352" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1701" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2298" />
                    <RANKING order="2" place="2" resultid="5387" />
                    <RANKING order="3" place="3" resultid="3743" />
                    <RANKING order="4" place="4" resultid="2636" />
                    <RANKING order="5" place="5" resultid="4144" />
                    <RANKING order="6" place="6" resultid="5083" />
                    <RANKING order="7" place="7" resultid="3233" />
                    <RANKING order="8" place="-1" resultid="3864" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1702" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3595" />
                    <RANKING order="2" place="2" resultid="5259" />
                    <RANKING order="3" place="3" resultid="4544" />
                    <RANKING order="4" place="4" resultid="4539" />
                    <RANKING order="5" place="5" resultid="4663" />
                    <RANKING order="6" place="-1" resultid="2219" />
                    <RANKING order="7" place="-1" resultid="2553" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1703" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5395" />
                    <RANKING order="2" place="2" resultid="4827" />
                    <RANKING order="3" place="3" resultid="3476" />
                    <RANKING order="4" place="4" resultid="3915" />
                    <RANKING order="5" place="5" resultid="5331" />
                    <RANKING order="6" place="6" resultid="4228" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1704" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3063" />
                    <RANKING order="2" place="2" resultid="4190" />
                    <RANKING order="3" place="3" resultid="4941" />
                    <RANKING order="4" place="4" resultid="4687" />
                    <RANKING order="5" place="5" resultid="3390" />
                    <RANKING order="6" place="6" resultid="3627" />
                    <RANKING order="7" place="7" resultid="2404" />
                    <RANKING order="8" place="8" resultid="3406" />
                    <RANKING order="9" place="9" resultid="3683" />
                    <RANKING order="10" place="10" resultid="3758" />
                    <RANKING order="11" place="11" resultid="3155" />
                    <RANKING order="12" place="12" resultid="2778" />
                    <RANKING order="13" place="13" resultid="4774" />
                    <RANKING order="14" place="-1" resultid="2011" />
                    <RANKING order="15" place="-1" resultid="3765" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1705" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4195" />
                    <RANKING order="2" place="2" resultid="5230" />
                    <RANKING order="3" place="3" resultid="3953" />
                    <RANKING order="4" place="4" resultid="3835" />
                    <RANKING order="5" place="5" resultid="4703" />
                    <RANKING order="6" place="6" resultid="2431" />
                    <RANKING order="7" place="7" resultid="2413" />
                    <RANKING order="8" place="8" resultid="3616" />
                    <RANKING order="9" place="-1" resultid="5121" />
                    <RANKING order="10" place="-1" resultid="2231" />
                    <RANKING order="11" place="-1" resultid="6212" />
                    <RANKING order="12" place="-1" resultid="2468" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1706" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2871" />
                    <RANKING order="2" place="2" resultid="5353" />
                    <RANKING order="3" place="3" resultid="3621" />
                    <RANKING order="4" place="4" resultid="3283" />
                    <RANKING order="5" place="5" resultid="5217" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1707" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2844" />
                    <RANKING order="2" place="2" resultid="1928" />
                    <RANKING order="3" place="3" resultid="3136" />
                    <RANKING order="4" place="4" resultid="4509" />
                    <RANKING order="5" place="5" resultid="4121" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1708" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3948" />
                    <RANKING order="2" place="2" resultid="4112" />
                    <RANKING order="3" place="3" resultid="1982" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1709" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1710" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1711" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1712" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7301" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7302" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7303" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7304" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7305" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7306" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7307" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7308" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7309" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7310" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7311" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1713" daytime="10:38" gender="F" number="38" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1714" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2064" />
                    <RANKING order="2" place="2" resultid="2421" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1715" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2919" />
                    <RANKING order="2" place="2" resultid="3807" />
                    <RANKING order="3" place="3" resultid="2729" />
                    <RANKING order="4" place="4" resultid="1970" />
                    <RANKING order="5" place="5" resultid="4393" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1716" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3253" />
                    <RANKING order="2" place="2" resultid="3257" />
                    <RANKING order="3" place="3" resultid="4835" />
                    <RANKING order="4" place="4" resultid="3057" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1717" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2169" />
                    <RANKING order="2" place="2" resultid="5184" />
                    <RANKING order="3" place="3" resultid="1858" />
                    <RANKING order="4" place="4" resultid="5287" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1718" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4594" />
                    <RANKING order="2" place="2" resultid="2346" />
                    <RANKING order="3" place="3" resultid="2146" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1719" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3322" />
                    <RANKING order="2" place="2" resultid="2111" />
                    <RANKING order="3" place="3" resultid="3083" />
                    <RANKING order="4" place="4" resultid="2475" />
                    <RANKING order="5" place="5" resultid="4980" />
                    <RANKING order="6" place="6" resultid="5042" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1720" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5177" />
                    <RANKING order="2" place="2" resultid="1936" />
                    <RANKING order="3" place="3" resultid="1921" />
                    <RANKING order="4" place="4" resultid="1956" />
                    <RANKING order="5" place="-1" resultid="2494" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1721" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4639" />
                    <RANKING order="2" place="2" resultid="5166" />
                    <RANKING order="3" place="3" resultid="3739" />
                    <RANKING order="4" place="-1" resultid="3183" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1722" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2857" />
                    <RANKING order="2" place="2" resultid="3959" />
                    <RANKING order="3" place="3" resultid="2505" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1723" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2029" />
                    <RANKING order="2" place="2" resultid="4965" />
                    <RANKING order="3" place="-1" resultid="4960" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1724" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4845" />
                    <RANKING order="2" place="2" resultid="4089" />
                    <RANKING order="3" place="3" resultid="4096" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1725" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4869" />
                    <RANKING order="2" place="2" resultid="2609" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1726" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1727" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3159" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1728" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1729" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7312" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7313" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7314" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7315" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7316" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7317" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1730" daytime="10:55" gender="M" number="39" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1731" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4236" />
                    <RANKING order="2" place="2" resultid="2072" />
                    <RANKING order="3" place="3" resultid="2094" />
                    <RANKING order="4" place="4" resultid="5100" />
                    <RANKING order="5" place="-1" resultid="5022" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1732" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2333" />
                    <RANKING order="2" place="2" resultid="2954" />
                    <RANKING order="3" place="3" resultid="5056" />
                    <RANKING order="4" place="4" resultid="3248" />
                    <RANKING order="5" place="5" resultid="2427" />
                    <RANKING order="6" place="6" resultid="2943" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1733" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2547" />
                    <RANKING order="2" place="2" resultid="3654" />
                    <RANKING order="3" place="3" resultid="5070" />
                    <RANKING order="4" place="4" resultid="4343" />
                    <RANKING order="5" place="4" resultid="3677" />
                    <RANKING order="6" place="6" resultid="2541" />
                    <RANKING order="7" place="7" resultid="5078" />
                    <RANKING order="8" place="-1" resultid="4151" />
                    <RANKING order="9" place="-1" resultid="6704" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1734" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3422" />
                    <RANKING order="2" place="2" resultid="2683" />
                    <RANKING order="3" place="3" resultid="3075" />
                    <RANKING order="4" place="4" resultid="5281" />
                    <RANKING order="5" place="5" resultid="3243" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1735" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2621" />
                    <RANKING order="2" place="2" resultid="2308" />
                    <RANKING order="3" place="3" resultid="3507" />
                    <RANKING order="4" place="4" resultid="4053" />
                    <RANKING order="5" place="-1" resultid="4551" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1736" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2566" />
                    <RANKING order="2" place="2" resultid="4852" />
                    <RANKING order="3" place="3" resultid="4664" />
                    <RANKING order="4" place="4" resultid="5035" />
                    <RANKING order="5" place="5" resultid="5092" />
                    <RANKING order="6" place="-1" resultid="2199" />
                    <RANKING order="7" place="-1" resultid="5405" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1737" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2711" />
                    <RANKING order="2" place="2" resultid="3041" />
                    <RANKING order="3" place="3" resultid="2480" />
                    <RANKING order="4" place="4" resultid="4080" />
                    <RANKING order="5" place="5" resultid="5243" />
                    <RANKING order="6" place="6" resultid="3100" />
                    <RANKING order="7" place="7" resultid="3398" />
                    <RANKING order="8" place="8" resultid="3734" />
                    <RANKING order="9" place="9" resultid="5400" />
                    <RANKING order="10" place="-1" resultid="4893" />
                    <RANKING order="11" place="-1" resultid="4209" />
                    <RANKING order="12" place="-1" resultid="3470" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1738" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4902" />
                    <RANKING order="2" place="2" resultid="4620" />
                    <RANKING order="3" place="3" resultid="5383" />
                    <RANKING order="4" place="4" resultid="4886" />
                    <RANKING order="5" place="5" resultid="4782" />
                    <RANKING order="6" place="6" resultid="3009" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1739" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4009" />
                    <RANKING order="2" place="2" resultid="2364" />
                    <RANKING order="3" place="3" resultid="5236" />
                    <RANKING order="4" place="4" resultid="3454" />
                    <RANKING order="5" place="5" resultid="2833" />
                    <RANKING order="6" place="6" resultid="4432" />
                    <RANKING order="7" place="7" resultid="4972" />
                    <RANKING order="8" place="8" resultid="3147" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1740" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5224" />
                    <RANKING order="2" place="2" resultid="5354" />
                    <RANKING order="3" place="3" resultid="2649" />
                    <RANKING order="4" place="4" resultid="3622" />
                    <RANKING order="5" place="-1" resultid="3995" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1741" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2372" />
                    <RANKING order="2" place="2" resultid="4695" />
                    <RANKING order="3" place="3" resultid="2534" />
                    <RANKING order="4" place="4" resultid="3608" />
                    <RANKING order="5" place="5" resultid="4709" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1742" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4113" />
                    <RANKING order="2" place="2" resultid="1983" />
                    <RANKING order="3" place="3" resultid="4159" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1743" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2325" />
                    <RANKING order="2" place="2" resultid="4911" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1744" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1745" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1746" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7318" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7319" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7320" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7321" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7322" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7323" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7324" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7325" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7326" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1747" daytime="11:16" gender="F" number="40" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1748" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3334" />
                    <RANKING order="2" place="2" resultid="2059" />
                    <RANKING order="3" place="3" resultid="3981" />
                    <RANKING order="4" place="4" resultid="2032" />
                    <RANKING order="5" place="5" resultid="3272" />
                    <RANKING order="6" place="-1" resultid="4874" />
                    <RANKING order="7" place="-1" resultid="5016" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1749" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1879" />
                    <RANKING order="2" place="2" resultid="3891" />
                    <RANKING order="3" place="3" resultid="2925" />
                    <RANKING order="4" place="4" resultid="4633" />
                    <RANKING order="5" place="5" resultid="3808" />
                    <RANKING order="6" place="6" resultid="4268" />
                    <RANKING order="7" place="7" resultid="3123" />
                    <RANKING order="8" place="-1" resultid="2959" />
                    <RANKING order="9" place="-1" resultid="2964" />
                    <RANKING order="10" place="-1" resultid="4400" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1750" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4811" />
                    <RANKING order="2" place="2" resultid="3258" />
                    <RANKING order="3" place="3" resultid="2642" />
                    <RANKING order="4" place="4" resultid="4386" />
                    <RANKING order="5" place="-1" resultid="2757" />
                    <RANKING order="6" place="-1" resultid="2764" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1751" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2304" />
                    <RANKING order="2" place="2" resultid="5376" />
                    <RANKING order="3" place="3" resultid="2627" />
                    <RANKING order="4" place="4" resultid="2690" />
                    <RANKING order="5" place="5" resultid="2786" />
                    <RANKING order="6" place="6" resultid="5185" />
                    <RANKING order="7" place="7" resultid="2136" />
                    <RANKING order="8" place="-1" resultid="5194" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1752" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4733" />
                    <RANKING order="2" place="-1" resultid="4655" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1753" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2112" />
                    <RANKING order="2" place="2" resultid="2162" />
                    <RANKING order="3" place="3" resultid="4175" />
                    <RANKING order="4" place="4" resultid="4168" />
                    <RANKING order="5" place="5" resultid="5043" />
                    <RANKING order="6" place="6" resultid="4282" />
                    <RANKING order="7" place="7" resultid="3176" />
                    <RANKING order="8" place="8" resultid="4934" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1754" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3017" />
                    <RANKING order="2" place="2" resultid="4681" />
                    <RANKING order="3" place="3" resultid="5178" />
                    <RANKING order="4" place="4" resultid="2154" />
                    <RANKING order="5" place="5" resultid="1978" />
                    <RANKING order="6" place="6" resultid="3414" />
                    <RANKING order="7" place="7" resultid="3068" />
                    <RANKING order="8" place="8" resultid="5171" />
                    <RANKING order="9" place="9" resultid="3583" />
                    <RANKING order="10" place="10" resultid="2495" />
                    <RANKING order="11" place="11" resultid="2461" />
                    <RANKING order="12" place="12" resultid="4921" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1755" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4105" />
                    <RANKING order="2" place="2" resultid="4274" />
                    <RANKING order="3" place="3" resultid="4183" />
                    <RANKING order="4" place="4" resultid="2397" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1756" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5159" />
                    <RANKING order="2" place="2" resultid="2658" />
                    <RANKING order="3" place="3" resultid="2822" />
                    <RANKING order="4" place="4" resultid="2882" />
                    <RANKING order="5" place="5" resultid="2677" />
                    <RANKING order="6" place="6" resultid="3168" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1757" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2878" />
                    <RANKING order="2" place="2" resultid="2028" />
                    <RANKING order="3" place="3" resultid="2452" />
                    <RANKING order="4" place="4" resultid="4966" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1758" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4097" />
                    <RANKING order="2" place="2" resultid="4090" />
                    <RANKING order="3" place="-1" resultid="5149" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1759" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4870" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1760" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3108" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1761" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3160" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1762" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1763" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7327" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7328" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7329" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7330" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7331" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7332" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7333" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7334" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7335" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1764" daytime="11:26" gender="M" number="41" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1765" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7491" />
                    <RANKING order="2" place="2" resultid="1895" />
                    <RANKING order="3" place="3" resultid="3843" />
                    <RANKING order="4" place="4" resultid="1866" />
                    <RANKING order="5" place="5" resultid="2443" />
                    <RANKING order="6" place="6" resultid="3783" />
                    <RANKING order="7" place="7" resultid="3812" />
                    <RANKING order="8" place="8" resultid="3789" />
                    <RANKING order="9" place="9" resultid="2080" />
                    <RANKING order="10" place="10" resultid="5101" />
                    <RANKING order="11" place="11" resultid="2088" />
                    <RANKING order="12" place="-1" resultid="5023" />
                    <RANKING order="13" place="-1" resultid="3907" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1766" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4417" />
                    <RANKING order="2" place="2" resultid="3771" />
                    <RANKING order="3" place="3" resultid="3601" />
                    <RANKING order="4" place="4" resultid="2937" />
                    <RANKING order="5" place="5" resultid="2908" />
                    <RANKING order="6" place="6" resultid="5128" />
                    <RANKING order="7" place="7" resultid="1886" />
                    <RANKING order="8" place="8" resultid="2930" />
                    <RANKING order="9" place="9" resultid="3857" />
                    <RANKING order="10" place="9" resultid="5113" />
                    <RANKING order="11" place="11" resultid="2948" />
                    <RANKING order="12" place="12" resultid="3870" />
                    <RANKING order="13" place="13" resultid="2671" />
                    <RANKING order="14" place="14" resultid="4501" />
                    <RANKING order="15" place="15" resultid="3209" />
                    <RANKING order="16" place="16" resultid="4133" />
                    <RANKING order="17" place="17" resultid="2772" />
                    <RANKING order="18" place="-1" resultid="4762" />
                    <RANKING order="19" place="-1" resultid="5115" />
                    <RANKING order="20" place="-1" resultid="5137" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1767" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4766" />
                    <RANKING order="2" place="2" resultid="3306" />
                    <RANKING order="3" place="3" resultid="2592" />
                    <RANKING order="4" place="4" resultid="3639" />
                    <RANKING order="5" place="5" resultid="3847" />
                    <RANKING order="6" place="6" resultid="3655" />
                    <RANKING order="7" place="6" resultid="4566" />
                    <RANKING order="8" place="8" resultid="5146" />
                    <RANKING order="9" place="9" resultid="4334" />
                    <RANKING order="10" place="10" resultid="4355" />
                    <RANKING order="11" place="11" resultid="3025" />
                    <RANKING order="12" place="12" resultid="5063" />
                    <RANKING order="13" place="13" resultid="2751" />
                    <RANKING order="14" place="13" resultid="4368" />
                    <RANKING order="15" place="15" resultid="4323" />
                    <RANKING order="16" place="16" resultid="4647" />
                    <RANKING order="17" place="16" resultid="4316" />
                    <RANKING order="18" place="18" resultid="4359" />
                    <RANKING order="19" place="19" resultid="4344" />
                    <RANKING order="20" place="20" resultid="3647" />
                    <RANKING order="21" place="21" resultid="2542" />
                    <RANKING order="22" place="22" resultid="2721" />
                    <RANKING order="23" place="23" resultid="4364" />
                    <RANKING order="24" place="-1" resultid="3750" />
                    <RANKING order="25" place="-1" resultid="4075" />
                    <RANKING order="26" place="-1" resultid="4797" />
                    <RANKING order="27" place="-1" resultid="5109" />
                    <RANKING order="28" place="-1" resultid="5141" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1768" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3431" />
                    <RANKING order="2" place="2" resultid="3423" />
                    <RANKING order="3" place="3" resultid="2684" />
                    <RANKING order="4" place="4" resultid="3374" />
                    <RANKING order="5" place="5" resultid="4424" />
                    <RANKING order="6" place="6" resultid="4375" />
                    <RANKING order="7" place="7" resultid="2314" />
                    <RANKING order="8" place="8" resultid="4560" />
                    <RANKING order="9" place="9" resultid="1962" />
                    <RANKING order="10" place="10" resultid="5086" />
                    <RANKING order="11" place="11" resultid="5346" />
                    <RANKING order="12" place="12" resultid="2318" />
                    <RANKING order="13" place="-1" resultid="2227" />
                    <RANKING order="14" place="-1" resultid="3855" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1769" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5368" />
                    <RANKING order="2" place="2" resultid="2183" />
                    <RANKING order="3" place="3" resultid="3221" />
                    <RANKING order="4" place="4" resultid="3361" />
                    <RANKING order="5" place="5" resultid="3523" />
                    <RANKING order="6" place="6" resultid="2309" />
                    <RANKING order="7" place="7" resultid="7495" />
                    <RANKING order="8" place="8" resultid="3032" />
                    <RANKING order="9" place="9" resultid="3295" />
                    <RANKING order="10" place="10" resultid="4304" />
                    <RANKING order="11" place="11" resultid="3463" />
                    <RANKING order="12" place="12" resultid="4024" />
                    <RANKING order="13" place="13" resultid="5458" />
                    <RANKING order="14" place="14" resultid="2191" />
                    <RANKING order="15" place="15" resultid="3508" />
                    <RANKING order="16" place="16" resultid="2637" />
                    <RANKING order="17" place="17" resultid="4725" />
                    <RANKING order="18" place="18" resultid="4019" />
                    <RANKING order="19" place="19" resultid="3115" />
                    <RANKING order="20" place="20" resultid="3234" />
                    <RANKING order="21" place="21" resultid="2236" />
                    <RANKING order="22" place="-1" resultid="2703" />
                    <RANKING order="23" place="-1" resultid="4037" />
                    <RANKING order="24" place="-1" resultid="5388" />
                    <RANKING order="25" place="-1" resultid="4552" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1770" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3596" />
                    <RANKING order="2" place="2" resultid="5048" />
                    <RANKING order="3" place="3" resultid="3267" />
                    <RANKING order="4" place="4" resultid="4545" />
                    <RANKING order="5" place="5" resultid="3090" />
                    <RANKING order="6" place="6" resultid="2567" />
                    <RANKING order="7" place="7" resultid="4853" />
                    <RANKING order="8" place="8" resultid="5274" />
                    <RANKING order="9" place="9" resultid="4718" />
                    <RANKING order="10" place="10" resultid="2208" />
                    <RANKING order="11" place="-1" resultid="2554" />
                    <RANKING order="12" place="-1" resultid="2597" />
                    <RANKING order="13" place="-1" resultid="3940" />
                    <RANKING order="14" place="-1" resultid="4250" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1771" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2559" />
                    <RANKING order="2" place="2" resultid="2481" />
                    <RANKING order="3" place="3" resultid="4031" />
                    <RANKING order="4" place="4" resultid="3899" />
                    <RANKING order="5" place="5" resultid="3477" />
                    <RANKING order="6" place="6" resultid="4248" />
                    <RANKING order="7" place="7" resultid="2605" />
                    <RANKING order="8" place="8" resultid="5361" />
                    <RANKING order="9" place="9" resultid="4242" />
                    <RANKING order="10" place="-1" resultid="4894" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1772" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4903" />
                    <RANKING order="2" place="2" resultid="3588" />
                    <RANKING order="3" place="3" resultid="2829" />
                    <RANKING order="4" place="4" resultid="4942" />
                    <RANKING order="5" place="5" resultid="3635" />
                    <RANKING order="6" place="6" resultid="2341" />
                    <RANKING order="7" place="7" resultid="4821" />
                    <RANKING order="8" place="8" resultid="2357" />
                    <RANKING order="9" place="9" resultid="3391" />
                    <RANKING order="10" place="10" resultid="4928" />
                    <RANKING order="11" place="11" resultid="4775" />
                    <RANKING order="12" place="-1" resultid="2012" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1773" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4297" />
                    <RANKING order="2" place="2" resultid="2892" />
                    <RANKING order="3" place="3" resultid="4010" />
                    <RANKING order="4" place="4" resultid="6213" />
                    <RANKING order="5" place="5" resultid="2587" />
                    <RANKING order="6" place="6" resultid="2886" />
                    <RANKING order="7" place="7" resultid="2379" />
                    <RANKING order="8" place="8" resultid="3836" />
                    <RANKING order="9" place="9" resultid="2432" />
                    <RANKING order="10" place="10" resultid="5122" />
                    <RANKING order="11" place="-1" resultid="2860" />
                    <RANKING order="12" place="-1" resultid="4754" />
                    <RANKING order="13" place="-1" resultid="5252" />
                    <RANKING order="14" place="-1" resultid="5432" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1774" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4062" />
                    <RANKING order="2" place="2" resultid="2872" />
                    <RANKING order="3" place="3" resultid="2456" />
                    <RANKING order="4" place="4" resultid="2650" />
                    <RANKING order="5" place="5" resultid="5211" />
                    <RANKING order="6" place="6" resultid="5218" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1775" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2373" />
                    <RANKING order="2" place="2" resultid="2499" />
                    <RANKING order="3" place="3" resultid="1929" />
                    <RANKING order="4" place="4" resultid="4126" />
                    <RANKING order="5" place="5" resultid="4710" />
                    <RANKING order="6" place="-1" resultid="3609" />
                    <RANKING order="7" place="-1" resultid="5203" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1776" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5198" />
                    <RANKING order="2" place="2" resultid="4160" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1777" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4613" />
                    <RANKING order="2" place="2" resultid="2448" />
                    <RANKING order="3" place="3" resultid="3944" />
                    <RANKING order="4" place="4" resultid="2326" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1778" agemax="89" agemin="85">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4201" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1779" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1780" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7336" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7337" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7338" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7339" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7340" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7341" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7342" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7343" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="7344" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="7345" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="7346" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="7347" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="7348" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="7349" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="7350" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="7351" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="7352" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="7353" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="7354" number="19" order="19" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1781" daytime="11:50" gender="F" number="42" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1782" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2422" />
                    <RANKING order="2" place="2" resultid="3663" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1783" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="1784" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2765" />
                    <RANKING order="2" place="2" resultid="2575" />
                    <RANKING order="3" place="3" resultid="3975" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1785" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2170" />
                    <RANKING order="2" place="2" resultid="1859" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1786" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3827" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1787" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2995" />
                    <RANKING order="2" place="2" resultid="3279" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1788" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2130" />
                    <RANKING order="2" place="2" resultid="1937" />
                    <RANKING order="3" place="3" resultid="2004" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1789" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1997" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1790" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="1791" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1792" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1793" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1794" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1795" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1796" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1797" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7355" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7356" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1798" daytime="12:09" gender="M" number="43" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1799" agemax="24" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3775" />
                    <RANKING order="2" place="2" resultid="1873" />
                    <RANKING order="3" place="-1" resultid="4920" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1800" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2334" />
                    <RANKING order="2" place="2" resultid="5133" />
                    <RANKING order="3" place="3" resultid="4216" />
                    <RANKING order="4" place="4" resultid="2914" />
                    <RANKING order="5" place="-1" resultid="2773" />
                    <RANKING order="6" place="-1" resultid="2696" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1801" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4382" />
                    <RANKING order="2" place="2" resultid="3447" />
                    <RANKING order="3" place="3" resultid="3493" />
                    <RANKING order="4" place="4" resultid="5079" />
                    <RANKING order="5" place="-1" resultid="5071" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1802" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3353" />
                    <RANKING order="2" place="2" resultid="2205" />
                    <RANKING order="3" place="3" resultid="3439" />
                    <RANKING order="4" place="4" resultid="4673" />
                    <RANKING order="5" place="-1" resultid="3516" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1803" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5369" />
                    <RANKING order="2" place="2" resultid="2299" />
                    <RANKING order="3" place="3" resultid="3524" />
                    <RANKING order="4" place="4" resultid="4043" />
                    <RANKING order="5" place="5" resultid="3033" />
                    <RANKING order="6" place="6" resultid="5339" />
                    <RANKING order="7" place="7" resultid="4145" />
                    <RANKING order="8" place="8" resultid="3865" />
                    <RANKING order="9" place="9" resultid="4726" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1804" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3705" />
                    <RANKING order="2" place="2" resultid="3312" />
                    <RANKING order="3" place="3" resultid="4223" />
                    <RANKING order="4" place="-1" resultid="5093" />
                    <RANKING order="5" place="-1" resultid="2220" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1805" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5247" />
                    <RANKING order="2" place="2" resultid="3471" />
                    <RANKING order="3" place="3" resultid="3101" />
                    <RANKING order="4" place="4" resultid="3714" />
                    <RANKING order="5" place="5" resultid="3916" />
                    <RANKING order="6" place="6" resultid="3567" />
                    <RANKING order="7" place="7" resultid="3002" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1806" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5239" />
                    <RANKING order="2" place="2" resultid="3368" />
                    <RANKING order="3" place="3" resultid="2814" />
                    <RANKING order="4" place="4" resultid="4191" />
                    <RANKING order="5" place="5" resultid="4887" />
                    <RANKING order="6" place="6" resultid="2405" />
                    <RANKING order="7" place="7" resultid="4929" />
                    <RANKING order="8" place="8" resultid="4783" />
                    <RANKING order="9" place="9" resultid="3407" />
                    <RANKING order="10" place="10" resultid="3010" />
                    <RANKING order="11" place="-1" resultid="4069" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1807" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2365" />
                    <RANKING order="2" place="2" resultid="3455" />
                    <RANKING order="3" place="3" resultid="5231" />
                    <RANKING order="4" place="4" resultid="3954" />
                    <RANKING order="5" place="5" resultid="4704" />
                    <RANKING order="6" place="6" resultid="4433" />
                    <RANKING order="7" place="7" resultid="4973" />
                    <RANKING order="8" place="8" resultid="3720" />
                    <RANKING order="9" place="9" resultid="3382" />
                    <RANKING order="10" place="-1" resultid="2717" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1808" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1809" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4696" />
                    <RANKING order="2" place="2" resultid="2535" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1810" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1811" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="1812" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="1813" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="1814" agemax="99" agemin="95" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7358" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7359" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="7360" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="7361" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="7362" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="7363" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="7364" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1815" daytime="13:13" gender="X" number="44" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1832" agemax="96" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2098" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1833" agemax="119" agemin="100">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2976" />
                    <RANKING order="2" place="2" resultid="2969" />
                    <RANKING order="3" place="3" resultid="4407" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1834" agemax="159" agemin="120">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7499" />
                    <RANKING order="2" place="2" resultid="2242" />
                    <RANKING order="3" place="3" resultid="7500" />
                    <RANKING order="4" place="-1" resultid="4745" />
                    <RANKING order="5" place="-1" resultid="2794" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1835" agemax="199" agemin="160">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2250" />
                    <RANKING order="2" place="-1" resultid="5425" />
                    <RANKING order="3" place="-1" resultid="3045" />
                    <RANKING order="4" place="-1" resultid="2788" />
                    <RANKING order="5" place="-1" resultid="4306" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1836" agemax="239" agemin="200">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5297" />
                    <RANKING order="2" place="2" resultid="2252" />
                    <RANKING order="3" place="-1" resultid="4988" />
                    <RANKING order="4" place="-1" resultid="3185" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1837" agemax="279" agemin="240">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5299" />
                    <RANKING order="2" place="-1" resultid="4987" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1838" agemax="319" agemin="280">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7498" />
                    <RANKING order="2" place="-1" resultid="2035" />
                    <RANKING order="3" place="-1" resultid="3191" />
                    <RANKING order="4" place="-1" resultid="6665" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1839" agemax="359" agemin="320" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="7502" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="7503" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="7504" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="NESTA" name="Miedzyszkolny Klub Sportowy &quot;Neptun&quot;" nation="POL" region="SZ">
          <CONTACT city="Stargard Szcz." email="prezes@mksneptun.pl" name="Ireneusz Drozd" phone="602731410" state="ZACHO" street="Os. Zachód B15" zip="73-110" />
          <ATHLETES>
            <ATHLETE birthdate="1973-01-19" firstname="Katarzyna" gender="F" lastname="Sawicka" nation="POL" athleteid="1852">
              <RESULTS>
                <RESULT eventid="1290" points="169" reactiontime="+74" swimtime="00:03:46.50" resultid="1854" lane="1" heatid="6877" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.27" />
                    <SPLIT distance="50" swimtime="00:00:48.55" />
                    <SPLIT distance="75" swimtime="00:01:15.81" />
                    <SPLIT distance="100" swimtime="00:01:43.84" />
                    <SPLIT distance="125" swimtime="00:02:13.83" />
                    <SPLIT distance="150" swimtime="00:02:44.36" />
                    <SPLIT distance="175" swimtime="00:03:16.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1781" points="201" reactiontime="+99" swimtime="00:07:39.43" resultid="1859" lane="6" heatid="7355">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.08" />
                    <SPLIT distance="50" swimtime="00:00:45.61" />
                    <SPLIT distance="75" swimtime="00:01:15.37" />
                    <SPLIT distance="100" swimtime="00:01:45.34" />
                    <SPLIT distance="125" swimtime="00:02:17.05" />
                    <SPLIT distance="150" swimtime="00:02:46.99" />
                    <SPLIT distance="175" swimtime="00:03:17.29" />
                    <SPLIT distance="200" swimtime="00:03:46.82" />
                    <SPLIT distance="225" swimtime="00:04:17.34" />
                    <SPLIT distance="250" swimtime="00:04:46.62" />
                    <SPLIT distance="275" swimtime="00:05:17.70" />
                    <SPLIT distance="300" swimtime="00:05:48.47" />
                    <SPLIT distance="325" swimtime="00:06:16.12" />
                    <SPLIT distance="350" swimtime="00:06:43.93" />
                    <SPLIT distance="375" swimtime="00:07:12.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1581" points="210" reactiontime="+90" swimtime="00:03:35.91" resultid="1857" lane="2" heatid="7068" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.52" />
                    <SPLIT distance="50" swimtime="00:00:43.92" />
                    <SPLIT distance="75" swimtime="00:01:13.26" />
                    <SPLIT distance="100" swimtime="00:01:42.23" />
                    <SPLIT distance="125" swimtime="00:02:12.78" />
                    <SPLIT distance="150" swimtime="00:02:43.60" />
                    <SPLIT distance="175" swimtime="00:03:10.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="192" reactiontime="+74" swimtime="00:01:41.84" resultid="1858" lane="3" heatid="7314" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.71" />
                    <SPLIT distance="50" swimtime="00:00:48.04" />
                    <SPLIT distance="75" swimtime="00:01:15.02" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="przekroczenie limitu 14:20:00" eventid="1058" status="DSQ" swimtime="00:14:53.04" resultid="1853" lane="5" heatid="6713" />
                <RESULT eventid="1358" status="DNS" swimtime="00:00:00.00" resultid="1855" lane="2" heatid="6895" entrytime="00:06:50.00" />
                <RESULT eventid="1409" status="DNS" swimtime="00:00:00.00" resultid="1856" lane="2" heatid="6999" entrytime="00:03:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-11-01" firstname="Oskar" gender="M" lastname="Wróblewski" nation="POL" license="S00116200598" athleteid="1860">
              <RESULTS>
                <RESULT eventid="1598" points="358" reactiontime="+74" swimtime="00:02:40.73" resultid="1864" lane="2" heatid="7079" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.28" />
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                    <SPLIT distance="75" swimtime="00:00:53.05" />
                    <SPLIT distance="100" swimtime="00:01:13.29" />
                    <SPLIT distance="125" swimtime="00:01:38.38" />
                    <SPLIT distance="150" swimtime="00:02:04.84" />
                    <SPLIT distance="175" swimtime="00:02:24.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="617" reactiontime="+72" swimtime="00:00:24.99" resultid="1866" lane="5" heatid="7353" entrytime="00:00:25.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="572" reactiontime="+77" swimtime="00:00:56.67" resultid="1862" lane="5" heatid="6845" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.55" />
                    <SPLIT distance="50" swimtime="00:00:26.62" />
                    <SPLIT distance="75" swimtime="00:00:41.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="473" reactiontime="+77" swimtime="00:00:34.88" resultid="1863" lane="7" heatid="6861" entrytime="00:00:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="462" reactiontime="+75" swimtime="00:00:29.68" resultid="1865" lane="1" heatid="7292" entrytime="00:00:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="411" reactiontime="+76" swimtime="00:01:08.76" resultid="1861" lane="7" heatid="6743" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.41" />
                    <SPLIT distance="50" swimtime="00:00:31.25" />
                    <SPLIT distance="75" swimtime="00:00:52.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-11-01" firstname="Michał" gender="M" lastname="Draczyński" nation="POL" license="S00816200080" athleteid="1867">
              <RESULTS>
                <RESULT eventid="1273" points="221" reactiontime="+90" swimtime="00:03:05.14" resultid="1869" lane="8" heatid="6874" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.34" />
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                    <SPLIT distance="75" swimtime="00:00:55.84" />
                    <SPLIT distance="100" swimtime="00:01:19.61" />
                    <SPLIT distance="125" swimtime="00:01:45.45" />
                    <SPLIT distance="150" swimtime="00:02:11.17" />
                    <SPLIT distance="175" swimtime="00:02:38.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="352" reactiontime="+87" swimtime="00:05:45.17" resultid="1873" lane="3" heatid="7363" entrytime="00:05:57.31">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.64" />
                    <SPLIT distance="50" swimtime="00:00:35.03" />
                    <SPLIT distance="75" swimtime="00:00:55.21" />
                    <SPLIT distance="100" swimtime="00:01:18.86" />
                    <SPLIT distance="125" swimtime="00:01:43.47" />
                    <SPLIT distance="150" swimtime="00:02:06.52" />
                    <SPLIT distance="175" swimtime="00:02:29.53" />
                    <SPLIT distance="200" swimtime="00:02:52.44" />
                    <SPLIT distance="225" swimtime="00:03:16.64" />
                    <SPLIT distance="250" swimtime="00:03:40.77" />
                    <SPLIT distance="275" swimtime="00:04:05.13" />
                    <SPLIT distance="300" swimtime="00:04:28.46" />
                    <SPLIT distance="325" swimtime="00:04:49.82" />
                    <SPLIT distance="350" swimtime="00:05:09.50" />
                    <SPLIT distance="375" swimtime="00:05:28.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="375" reactiontime="+83" swimtime="00:02:56.67" resultid="1870" lane="2" heatid="7010" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.79" />
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                    <SPLIT distance="75" swimtime="00:01:00.36" />
                    <SPLIT distance="100" swimtime="00:01:23.01" />
                    <SPLIT distance="125" swimtime="00:01:46.62" />
                    <SPLIT distance="150" swimtime="00:02:10.01" />
                    <SPLIT distance="175" swimtime="00:02:33.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="322" reactiontime="+87" swimtime="00:02:46.60" resultid="1871" lane="5" heatid="7079" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.55" />
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                    <SPLIT distance="75" swimtime="00:00:56.44" />
                    <SPLIT distance="100" swimtime="00:01:17.93" />
                    <SPLIT distance="125" swimtime="00:01:41.66" />
                    <SPLIT distance="150" swimtime="00:02:05.22" />
                    <SPLIT distance="175" swimtime="00:02:25.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="403" reactiontime="+86" swimtime="00:01:19.73" resultid="1872" lane="4" heatid="7310" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.30" />
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                    <SPLIT distance="75" swimtime="00:00:58.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="425" reactiontime="+83" swimtime="00:01:02.54" resultid="1868" lane="8" heatid="6845" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.20" />
                    <SPLIT distance="50" swimtime="00:00:29.70" />
                    <SPLIT distance="75" swimtime="00:00:46.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AZWAW" name="Azs Awf Warszawa" nation="POL">
          <CONTACT city="Warszawa" name="Gołębiowska" phone="504-794-417" street="Marymoncka 34" zip="01-813" />
          <ATHLETES>
            <ATHLETE birthdate="1982-02-23" firstname="Joanna" gender="F" lastname="Gołębiowska" nation="POL" license="S00114100002" athleteid="1875">
              <RESULTS>
                <RESULT comment="Rekord Polski " eventid="1187" points="722" reactiontime="+71" swimtime="00:00:58.93" resultid="1876" lane="4" heatid="6828" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.48" />
                    <SPLIT distance="50" swimtime="00:00:28.57" />
                    <SPLIT distance="75" swimtime="00:00:43.92" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1445" points="693" reactiontime="+69" swimtime="00:01:03.95" resultid="1877" lane="4" heatid="7014" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.68" />
                    <SPLIT distance="50" swimtime="00:00:30.05" />
                    <SPLIT distance="75" swimtime="00:00:47.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="668" reactiontime="+68" swimtime="00:00:29.12" resultid="1878" lane="4" heatid="7280" entrytime="00:00:29.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.62" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1747" points="677" reactiontime="+68" swimtime="00:00:27.29" resultid="1879" lane="4" heatid="7335" entrytime="00:00:28.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Małgorzata" gender="F" lastname="Młyńczak" nation="POL" athleteid="5011">
              <RESULTS>
                <RESULT eventid="1513" points="307" reactiontime="+96" swimtime="00:00:35.52" resultid="5015" lane="3" heatid="7044" entrytime="00:00:36.33">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="280" reactiontime="+87" swimtime="00:00:46.31" resultid="5012" heatid="6851" entrytime="00:00:46.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" status="DNS" swimtime="00:00:00.00" resultid="5013" heatid="7278" entrytime="00:00:42.55" />
                <RESULT eventid="1679" status="DNS" swimtime="00:00:00.00" resultid="5014" lane="5" heatid="7298" entrytime="00:01:43.80" />
                <RESULT eventid="1747" status="DNS" swimtime="00:00:00.00" resultid="5016" lane="4" heatid="7331" entrytime="00:00:36.33" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-01-01" firstname="Łukasz" gender="M" lastname="Stąpor" nation="POL" athleteid="5017">
              <RESULTS>
                <RESULT eventid="1530" points="397" reactiontime="+90" swimtime="00:00:28.93" resultid="5020" lane="3" heatid="7047" entrytime="00:00:33.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="321" reactiontime="+80" swimtime="00:00:35.71" resultid="5019" lane="6" heatid="7038" entrytime="00:00:35.56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="5021" lane="7" heatid="7286" entrytime="00:00:34.50" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="5018" lane="3" heatid="6839" entrytime="00:01:06.50" />
                <RESULT eventid="1730" status="DNS" swimtime="00:00:00.00" resultid="5022" lane="4" heatid="7323" entrytime="00:01:18.00" />
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="5023" lane="6" heatid="7340" entrytime="00:00:33.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CIPOZ" name="CitiZen Poznań" nation="POL" region="WIE">
          <CONTACT email="sport@cityzenclub.pl" />
          <ATHLETES>
            <ATHLETE birthdate="1985-01-01" firstname="Tadeusz" gender="M" lastname="Gołembiewski" nation="POL" athleteid="1881">
              <RESULTS>
                <RESULT eventid="1462" points="534" reactiontime="+76" swimtime="00:01:02.09" resultid="1883" lane="7" heatid="7023" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.37" />
                    <SPLIT distance="50" swimtime="00:00:28.65" />
                    <SPLIT distance="75" swimtime="00:00:45.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="590" reactiontime="+74" swimtime="00:00:56.09" resultid="1882" lane="7" heatid="6846" entrytime="00:00:55.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.59" />
                    <SPLIT distance="50" swimtime="00:00:26.31" />
                    <SPLIT distance="75" swimtime="00:00:40.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="547" reactiontime="+76" swimtime="00:00:28.06" resultid="1885" lane="7" heatid="7293" entrytime="00:00:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="454" reactiontime="+71" swimtime="00:00:31.83" resultid="1884" lane="4" heatid="7042" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="554" reactiontime="+75" swimtime="00:00:25.91" resultid="1886" lane="4" heatid="7353" entrytime="00:00:25.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-01-01" firstname="Marco" gender="M" lastname="Foelske" nation="POL" athleteid="1887">
              <RESULTS>
                <RESULT eventid="1496" points="358" reactiontime="+71" swimtime="00:00:34.46" resultid="1891" lane="1" heatid="7040" entrytime="00:00:33.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="289" reactiontime="+72" swimtime="00:02:52.24" resultid="1890" lane="7" heatid="6885" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.45" />
                    <SPLIT distance="50" swimtime="00:00:38.98" />
                    <SPLIT distance="75" swimtime="00:01:00.72" />
                    <SPLIT distance="100" swimtime="00:01:23.20" />
                    <SPLIT distance="125" swimtime="00:01:46.29" />
                    <SPLIT distance="150" swimtime="00:02:09.09" />
                    <SPLIT distance="175" swimtime="00:02:31.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="307" reactiontime="+90" swimtime="00:01:15.78" resultid="1888" lane="5" heatid="6739" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.36" />
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                    <SPLIT distance="75" swimtime="00:00:57.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="337" reactiontime="+96" swimtime="00:00:39.04" resultid="1889" heatid="6861" entrytime="00:00:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Tomasz" gender="M" lastname="Kawicki" nation="POL" athleteid="1892">
              <RESULTS>
                <RESULT eventid="1764" points="628" reactiontime="+69" swimtime="00:00:24.84" resultid="1895" lane="7" heatid="7354" entrytime="00:00:24.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="584" reactiontime="+75" swimtime="00:00:27.46" resultid="1894" lane="6" heatid="7293" entrytime="00:00:27.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="528" swimtime="00:01:03.27" resultid="1893" lane="8" heatid="6745" entrytime="00:01:04.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Mikołaj" gender="M" lastname="Grzesiak" nation="POL" athleteid="1902">
              <RESULTS>
                <RESULT eventid="1143" points="328" swimtime="00:21:07.78" resultid="1903" lane="5" heatid="6751" entrytime="00:22:14.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1177" status="DNS" swimtime="00:00:00.00" resultid="1905" lane="2" heatid="6810" entrytime="00:01:45.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1881" number="1" />
                    <RELAYPOSITION athleteid="1902" number="2" />
                    <RELAYPOSITION athleteid="1892" number="3" />
                    <RELAYPOSITION athleteid="1887" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MAGDY" name="Gdynia Masters" nation="POL">
          <CONTACT email="misiek@am.gdynia.pl" name="Mysiak Katarzyna" />
          <ATHLETES>
            <ATHLETE birthdate="1961-01-01" firstname="Katarzyna" gender="F" lastname="Mysiak" nation="POL" athleteid="1915">
              <RESULTS>
                <RESULT eventid="1058" points="195" swimtime="00:14:12.04" resultid="1916" lane="2" heatid="6714" entrytime="00:14:16.00" />
                <RESULT eventid="1713" points="205" reactiontime="+79" swimtime="00:01:39.51" resultid="1921" lane="1" heatid="7315" entrytime="00:01:39.32">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.62" />
                    <SPLIT distance="50" swimtime="00:00:47.42" />
                    <SPLIT distance="75" swimtime="00:01:14.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1581" points="196" reactiontime="+96" swimtime="00:03:41.00" resultid="1919" lane="8" heatid="7069" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.48" />
                    <SPLIT distance="50" swimtime="00:00:47.44" />
                    <SPLIT distance="75" swimtime="00:01:16.50" />
                    <SPLIT distance="100" swimtime="00:01:43.23" />
                    <SPLIT distance="125" swimtime="00:02:17.28" />
                    <SPLIT distance="150" swimtime="00:02:50.79" />
                    <SPLIT distance="175" swimtime="00:03:17.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="198" reactiontime="+77" swimtime="00:03:34.72" resultid="1917" lane="2" heatid="6877" entrytime="00:03:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.99" />
                    <SPLIT distance="50" swimtime="00:00:47.97" />
                    <SPLIT distance="75" swimtime="00:01:16.36" />
                    <SPLIT distance="100" swimtime="00:01:43.85" />
                    <SPLIT distance="125" swimtime="00:02:11.71" />
                    <SPLIT distance="150" swimtime="00:02:40.91" />
                    <SPLIT distance="175" swimtime="00:03:08.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="246" reactiontime="+72" swimtime="00:00:44.12" resultid="1918" lane="5" heatid="7028" entrytime="00:00:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="193" reactiontime="+97" swimtime="00:00:44.03" resultid="1920" lane="4" heatid="7277" entrytime="00:00:43.18">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1939-01-01" firstname="Andrzej" gender="M" lastname="Skwarło" nation="POL" athleteid="1922">
              <RESULTS>
                <RESULT eventid="1109" points="146" reactiontime="+97" swimtime="00:01:36.98" resultid="1923" lane="2" heatid="6732" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.55" />
                    <SPLIT distance="50" swimtime="00:00:46.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="139" reactiontime="+102" swimtime="00:03:40.21" resultid="1927" lane="6" heatid="7073" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.04" />
                    <SPLIT distance="50" swimtime="00:00:50.18" />
                    <SPLIT distance="75" swimtime="00:01:19.51" />
                    <SPLIT distance="100" swimtime="00:01:46.53" />
                    <SPLIT distance="125" swimtime="00:02:18.29" />
                    <SPLIT distance="150" swimtime="00:02:49.17" />
                    <SPLIT distance="175" swimtime="00:03:15.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="165" reactiontime="+107" swimtime="00:03:52.28" resultid="1926" lane="5" heatid="7004" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.99" />
                    <SPLIT distance="50" swimtime="00:00:50.34" />
                    <SPLIT distance="75" swimtime="00:01:20.10" />
                    <SPLIT distance="100" swimtime="00:01:50.53" />
                    <SPLIT distance="125" swimtime="00:02:21.97" />
                    <SPLIT distance="150" swimtime="00:02:53.14" />
                    <SPLIT distance="175" swimtime="00:03:23.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="243" reactiontime="+103" swimtime="00:00:43.50" resultid="1924" lane="5" heatid="6857" entrytime="00:00:42.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="213" reactiontime="+105" swimtime="00:01:38.52" resultid="1928" lane="2" heatid="7305" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.46" />
                    <SPLIT distance="50" swimtime="00:00:45.53" />
                    <SPLIT distance="75" swimtime="00:01:11.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="178" reactiontime="+79" swimtime="00:00:37.80" resultid="1929" lane="1" heatid="7338" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.24" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G 7" eventid="1307" reactiontime="+96" status="DSQ" swimtime="00:03:47.58" resultid="1925" lane="7" heatid="6882" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.71" />
                    <SPLIT distance="50" swimtime="00:00:49.30" />
                    <SPLIT distance="75" swimtime="00:01:17.57" />
                    <SPLIT distance="100" swimtime="00:01:46.19" />
                    <SPLIT distance="125" swimtime="00:02:19.48" />
                    <SPLIT distance="150" swimtime="00:02:48.66" />
                    <SPLIT distance="175" swimtime="00:03:18.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Renata" gender="F" lastname="Polańczyk" nation="POL" athleteid="1930">
              <RESULTS>
                <RESULT eventid="1781" points="174" reactiontime="+115" swimtime="00:08:02.22" resultid="1937" lane="5" heatid="7355" entrytime="00:08:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.68" />
                    <SPLIT distance="50" swimtime="00:00:52.21" />
                    <SPLIT distance="75" swimtime="00:01:22.87" />
                    <SPLIT distance="100" swimtime="00:01:53.69" />
                    <SPLIT distance="125" swimtime="00:02:22.34" />
                    <SPLIT distance="150" swimtime="00:02:50.09" />
                    <SPLIT distance="175" swimtime="00:03:17.31" />
                    <SPLIT distance="200" swimtime="00:03:44.42" />
                    <SPLIT distance="225" swimtime="00:04:22.50" />
                    <SPLIT distance="250" swimtime="00:05:00.21" />
                    <SPLIT distance="275" swimtime="00:05:38.54" />
                    <SPLIT distance="300" swimtime="00:06:16.15" />
                    <SPLIT distance="325" swimtime="00:06:44.11" />
                    <SPLIT distance="350" swimtime="00:07:11.08" />
                    <SPLIT distance="375" swimtime="00:07:37.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="200" reactiontime="+112" swimtime="00:06:52.46" resultid="1933" lane="4" heatid="6895" entrytime="00:06:46.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.30" />
                    <SPLIT distance="50" swimtime="00:00:44.23" />
                    <SPLIT distance="75" swimtime="00:01:08.88" />
                    <SPLIT distance="100" swimtime="00:01:34.70" />
                    <SPLIT distance="125" swimtime="00:02:01.39" />
                    <SPLIT distance="150" swimtime="00:02:27.71" />
                    <SPLIT distance="175" swimtime="00:02:54.25" />
                    <SPLIT distance="200" swimtime="00:03:20.49" />
                    <SPLIT distance="225" swimtime="00:03:47.71" />
                    <SPLIT distance="250" swimtime="00:04:14.27" />
                    <SPLIT distance="275" swimtime="00:04:41.04" />
                    <SPLIT distance="300" swimtime="00:05:07.91" />
                    <SPLIT distance="325" swimtime="00:05:34.80" />
                    <SPLIT distance="350" swimtime="00:06:02.06" />
                    <SPLIT distance="375" swimtime="00:06:28.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="209" reactiontime="+76" swimtime="00:01:38.98" resultid="1936" lane="2" heatid="7315" entrytime="00:01:36.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.01" />
                    <SPLIT distance="50" swimtime="00:00:48.11" />
                    <SPLIT distance="75" swimtime="00:01:14.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="215" reactiontime="+80" swimtime="00:03:28.92" resultid="1932" lane="5" heatid="6877" entrytime="00:03:31.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.56" />
                    <SPLIT distance="50" swimtime="00:00:48.59" />
                    <SPLIT distance="75" swimtime="00:01:14.93" />
                    <SPLIT distance="100" swimtime="00:01:41.46" />
                    <SPLIT distance="125" swimtime="00:02:08.73" />
                    <SPLIT distance="150" swimtime="00:02:36.10" />
                    <SPLIT distance="175" swimtime="00:03:03.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1058" points="190" swimtime="00:14:19.37" resultid="1931" lane="5" heatid="6714" entrytime="00:13:38.00" />
                <RESULT eventid="1445" status="DNS" swimtime="00:00:00.00" resultid="1934" lane="7" heatid="7013" entrytime="00:01:47.20" />
                <RESULT eventid="1547" status="DNS" swimtime="00:00:00.00" resultid="1935" lane="7" heatid="7050" entrytime="00:03:31.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-01-01" firstname="Zuzanna" gender="F" lastname="Drążkiewicz" nation="POL" athleteid="1938">
              <RESULTS>
                <RESULT eventid="1679" points="49" reactiontime="+118" swimtime="00:02:56.99" resultid="1943" lane="6" heatid="7295">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:40.64" />
                    <SPLIT distance="50" swimtime="00:01:25.95" />
                    <SPLIT distance="75" swimtime="00:02:12.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="48" reactiontime="+109" swimtime="00:01:23.03" resultid="1940" lane="3" heatid="6847">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:38.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="46" reactiontime="+191" swimtime="00:02:26.73" resultid="1939" lane="5" heatid="6821">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.64" />
                    <SPLIT distance="50" swimtime="00:01:03.13" />
                    <SPLIT distance="75" swimtime="00:01:42.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="68" reactiontime="+105" swimtime="00:00:58.56" resultid="4921" lane="5" heatid="7327">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1409" status="DNS" swimtime="00:00:00.00" resultid="1941" lane="1" heatid="6997" />
                <RESULT eventid="1547" status="DNS" swimtime="00:00:00.00" resultid="1942" lane="2" heatid="7048" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-01" firstname="Maja" gender="F" lastname="Szaduro" nation="POL" athleteid="1944">
              <RESULTS>
                <RESULT eventid="1222" points="317" reactiontime="+102" swimtime="00:00:44.41" resultid="1946" lane="2" heatid="6851" entrytime="00:00:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1581" points="194" reactiontime="+107" swimtime="00:03:41.83" resultid="1948" lane="4" heatid="7068" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.13" />
                    <SPLIT distance="50" swimtime="00:00:47.58" />
                    <SPLIT distance="75" swimtime="00:01:15.81" />
                    <SPLIT distance="100" swimtime="00:01:46.17" />
                    <SPLIT distance="125" swimtime="00:02:15.59" />
                    <SPLIT distance="150" swimtime="00:02:44.89" />
                    <SPLIT distance="175" swimtime="00:03:12.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1409" points="292" reactiontime="+106" swimtime="00:03:31.31" resultid="1947" heatid="7000" entrytime="00:03:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.06" />
                    <SPLIT distance="50" swimtime="00:00:47.52" />
                    <SPLIT distance="75" swimtime="00:01:13.54" />
                    <SPLIT distance="100" swimtime="00:01:41.06" />
                    <SPLIT distance="125" swimtime="00:02:09.17" />
                    <SPLIT distance="150" swimtime="00:02:36.91" />
                    <SPLIT distance="175" swimtime="00:03:03.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="292" reactiontime="+112" swimtime="00:01:38.07" resultid="1949" lane="4" heatid="7298" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.63" />
                    <SPLIT distance="50" swimtime="00:00:46.23" />
                    <SPLIT distance="75" swimtime="00:01:11.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="217" reactiontime="+106" swimtime="00:01:37.76" resultid="1945" lane="8" heatid="6726" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.43" />
                    <SPLIT distance="50" swimtime="00:00:45.81" />
                    <SPLIT distance="75" swimtime="00:01:11.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-01" firstname="Anna" gender="F" lastname="Krzysztofik" nation="POL" athleteid="1950">
              <RESULTS>
                <RESULT eventid="1409" points="235" reactiontime="+99" swimtime="00:03:47.07" resultid="1954" lane="4" heatid="6999" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.97" />
                    <SPLIT distance="50" swimtime="00:00:51.35" />
                    <SPLIT distance="75" swimtime="00:01:19.23" />
                    <SPLIT distance="100" swimtime="00:01:47.64" />
                    <SPLIT distance="125" swimtime="00:02:17.33" />
                    <SPLIT distance="150" swimtime="00:02:47.15" />
                    <SPLIT distance="175" swimtime="00:03:16.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="219" reactiontime="+118" swimtime="00:01:47.96" resultid="1955" heatid="7299" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.85" />
                    <SPLIT distance="50" swimtime="00:00:50.90" />
                    <SPLIT distance="75" swimtime="00:01:18.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="158" reactiontime="+86" swimtime="00:01:48.55" resultid="1956" heatid="7315" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.75" />
                    <SPLIT distance="50" swimtime="00:00:53.90" />
                    <SPLIT distance="75" swimtime="00:01:21.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1058" points="140" swimtime="00:15:50.66" resultid="1951" heatid="6714" entrytime="00:15:30.00" />
                <RESULT eventid="1290" points="180" reactiontime="+85" swimtime="00:03:41.52" resultid="1952" lane="6" heatid="6877" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.78" />
                    <SPLIT distance="50" swimtime="00:00:52.30" />
                    <SPLIT distance="75" swimtime="00:01:19.26" />
                    <SPLIT distance="100" swimtime="00:01:47.89" />
                    <SPLIT distance="125" swimtime="00:02:16.01" />
                    <SPLIT distance="150" swimtime="00:02:45.41" />
                    <SPLIT distance="175" swimtime="00:03:14.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" status="DNS" swimtime="00:00:00.00" resultid="1953" heatid="6895" entrytime="00:07:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-01" firstname="Kamil" gender="M" lastname="Plata" nation="POL" athleteid="1957">
              <RESULTS>
                <RESULT eventid="1645" points="322" reactiontime="+94" swimtime="00:00:33.49" resultid="1961" lane="3" heatid="7286" entrytime="00:00:34.28">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="267" reactiontime="+95" swimtime="00:02:39.71" resultid="1960" lane="3" heatid="7060" entrytime="00:02:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.27" />
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                    <SPLIT distance="75" swimtime="00:00:54.53" />
                    <SPLIT distance="100" swimtime="00:01:15.23" />
                    <SPLIT distance="125" swimtime="00:01:36.46" />
                    <SPLIT distance="150" swimtime="00:01:57.91" />
                    <SPLIT distance="175" swimtime="00:02:20.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="344" reactiontime="+93" swimtime="00:00:30.35" resultid="1962" lane="8" heatid="7344" entrytime="00:00:30.19">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="320" reactiontime="+89" swimtime="00:01:08.76" resultid="1958" lane="3" heatid="6837" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.95" />
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                    <SPLIT distance="75" swimtime="00:00:49.74" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="04 " eventid="1462" reactiontime="+84" status="DSQ" swimtime="00:00:00.00" resultid="1959" lane="6" heatid="7018" entrytime="00:01:25.23">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.14" />
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                    <SPLIT distance="75" swimtime="00:00:57.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-01" firstname="Beata" gender="F" lastname="Niewiadomska" nation="POL" athleteid="1963">
              <RESULTS>
                <RESULT eventid="1256" points="306" reactiontime="+98" swimtime="00:03:04.25" resultid="1965" lane="3" heatid="6868" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.53" />
                    <SPLIT distance="50" swimtime="00:00:40.20" />
                    <SPLIT distance="75" swimtime="00:01:02.92" />
                    <SPLIT distance="100" swimtime="00:01:26.58" />
                    <SPLIT distance="125" swimtime="00:01:51.08" />
                    <SPLIT distance="150" swimtime="00:02:15.23" />
                    <SPLIT distance="175" swimtime="00:02:40.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1445" points="337" reactiontime="+95" swimtime="00:01:21.29" resultid="1967" lane="7" heatid="7014" entrytime="00:01:19.56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.53" />
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                    <SPLIT distance="75" swimtime="00:00:59.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1058" points="308" swimtime="00:12:11.57" resultid="1964" lane="6" heatid="6715" entrytime="00:11:50.00" />
                <RESULT eventid="1713" points="338" reactiontime="+68" swimtime="00:01:24.36" resultid="1970" lane="8" heatid="7317" entrytime="00:01:21.86">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.91" />
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                    <SPLIT distance="75" swimtime="00:01:02.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="336" reactiontime="+94" swimtime="00:05:47.10" resultid="1966" lane="4" heatid="6897" entrytime="00:05:40.21">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.44" />
                    <SPLIT distance="50" swimtime="00:00:38.67" />
                    <SPLIT distance="75" swimtime="00:00:59.14" />
                    <SPLIT distance="100" swimtime="00:01:20.25" />
                    <SPLIT distance="125" swimtime="00:01:41.43" />
                    <SPLIT distance="150" swimtime="00:02:03.12" />
                    <SPLIT distance="175" swimtime="00:02:24.67" />
                    <SPLIT distance="200" swimtime="00:02:46.94" />
                    <SPLIT distance="225" swimtime="00:03:08.95" />
                    <SPLIT distance="250" swimtime="00:03:31.37" />
                    <SPLIT distance="275" swimtime="00:03:53.64" />
                    <SPLIT distance="300" swimtime="00:04:16.29" />
                    <SPLIT distance="325" swimtime="00:04:39.10" />
                    <SPLIT distance="350" swimtime="00:05:01.95" />
                    <SPLIT distance="375" swimtime="00:05:24.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="365" reactiontime="+87" swimtime="00:00:35.61" resultid="1969" lane="4" heatid="7279" entrytime="00:00:34.16">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="1968" lane="3" heatid="7029" entrytime="00:00:39.14" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Katarzyna" gender="F" lastname="Mazurek" nation="POL" athleteid="1971">
              <RESULTS>
                <RESULT eventid="1222" points="379" reactiontime="+87" swimtime="00:00:41.85" resultid="1974" lane="2" heatid="6852" entrytime="00:00:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1445" points="211" reactiontime="+96" swimtime="00:01:35.00" resultid="1975" lane="5" heatid="7013" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.06" />
                    <SPLIT distance="50" swimtime="00:00:42.84" />
                    <SPLIT distance="75" swimtime="00:01:08.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1581" points="204" reactiontime="+95" swimtime="00:03:38.09" resultid="1976" lane="3" heatid="7068" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.54" />
                    <SPLIT distance="50" swimtime="00:00:45.88" />
                    <SPLIT distance="75" swimtime="00:02:14.31" />
                    <SPLIT distance="100" swimtime="00:01:44.64" />
                    <SPLIT distance="125" swimtime="00:03:12.49" />
                    <SPLIT distance="150" swimtime="00:02:44.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="253" reactiontime="+95" swimtime="00:00:40.22" resultid="1977" lane="7" heatid="7278" entrytime="00:00:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="268" reactiontime="+97" swimtime="00:01:31.09" resultid="1972" lane="6" heatid="6727" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.72" />
                    <SPLIT distance="50" swimtime="00:00:42.98" />
                    <SPLIT distance="75" swimtime="00:01:08.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="256" reactiontime="+94" swimtime="00:01:23.24" resultid="1973" lane="2" heatid="6825" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.09" />
                    <SPLIT distance="50" swimtime="00:00:38.79" />
                    <SPLIT distance="75" swimtime="00:01:00.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="303" reactiontime="+81" swimtime="00:00:35.67" resultid="1978" lane="3" heatid="7332" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1934-01-01" firstname="Józef" gender="M" lastname="Kwias" nation="POL" athleteid="1979">
              <RESULTS>
                <RESULT eventid="1730" points="41" reactiontime="+93" swimtime="00:02:31.32" resultid="1983" lane="6" heatid="7319" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.38" />
                    <SPLIT distance="50" swimtime="00:01:13.28" />
                    <SPLIT distance="75" swimtime="00:01:53.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="55" swimtime="00:02:34.17" resultid="1982" lane="4" heatid="7302" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.37" />
                    <SPLIT distance="50" swimtime="00:01:12.73" />
                    <SPLIT distance="75" swimtime="00:01:54.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="41" reactiontime="+98" swimtime="00:01:10.59" resultid="1981" heatid="7033" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:33.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="60" swimtime="00:01:09.39" resultid="1980" lane="5" heatid="6854" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:33.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-01-01" firstname="Stefania" gender="F" lastname="Kowalska" nation="POL" athleteid="1984">
              <RESULTS>
                <RESULT eventid="1222" points="127" reactiontime="+91" swimtime="00:01:00.18" resultid="1986" lane="3" heatid="6848" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1409" points="90" reactiontime="+101" swimtime="00:05:12.38" resultid="1987" lane="7" heatid="6998" entrytime="00:04:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:33.48" />
                    <SPLIT distance="50" swimtime="00:01:11.28" />
                    <SPLIT distance="75" swimtime="00:01:51.74" />
                    <SPLIT distance="100" swimtime="00:02:33.05" />
                    <SPLIT distance="125" swimtime="00:03:15.29" />
                    <SPLIT distance="150" swimtime="00:03:57.65" />
                    <SPLIT distance="175" swimtime="00:04:38.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="62" reactiontime="+97" swimtime="00:01:04.03" resultid="1988" lane="2" heatid="7275" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="86" reactiontime="+124" swimtime="00:02:13.14" resultid="1985" lane="4" heatid="6723" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.29" />
                    <SPLIT distance="50" swimtime="00:01:07.24" />
                    <SPLIT distance="75" swimtime="00:01:41.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="109" reactiontime="+98" swimtime="00:02:16.20" resultid="1989" lane="7" heatid="7296" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.68" />
                    <SPLIT distance="50" swimtime="00:01:06.57" />
                    <SPLIT distance="75" swimtime="00:01:43.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-01" firstname="Barbara" gender="F" lastname="Chomicka" nation="POL" athleteid="1990">
              <RESULTS>
                <RESULT eventid="1781" points="130" reactiontime="+105" swimtime="00:08:51.68" resultid="1997" lane="2" heatid="7355" entrytime="00:09:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.04" />
                    <SPLIT distance="50" swimtime="00:00:59.64" />
                    <SPLIT distance="75" swimtime="00:01:34.41" />
                    <SPLIT distance="100" swimtime="00:02:10.42" />
                    <SPLIT distance="125" swimtime="00:02:45.10" />
                    <SPLIT distance="150" swimtime="00:03:19.95" />
                    <SPLIT distance="175" swimtime="00:03:54.57" />
                    <SPLIT distance="200" swimtime="00:04:29.93" />
                    <SPLIT distance="225" swimtime="00:05:05.23" />
                    <SPLIT distance="250" swimtime="00:05:41.30" />
                    <SPLIT distance="275" swimtime="00:06:16.32" />
                    <SPLIT distance="300" swimtime="00:06:51.48" />
                    <SPLIT distance="325" swimtime="00:07:22.69" />
                    <SPLIT distance="350" swimtime="00:07:54.32" />
                    <SPLIT distance="375" swimtime="00:08:25.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="101" reactiontime="+102" swimtime="00:04:26.11" resultid="1993" lane="5" heatid="6867" entrytime="00:04:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.00" />
                    <SPLIT distance="50" swimtime="00:00:59.79" />
                    <SPLIT distance="75" swimtime="00:01:33.47" />
                    <SPLIT distance="100" swimtime="00:02:07.99" />
                    <SPLIT distance="125" swimtime="00:02:43.27" />
                    <SPLIT distance="150" swimtime="00:03:17.74" />
                    <SPLIT distance="175" swimtime="00:03:52.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1409" points="168" reactiontime="+104" swimtime="00:04:13.70" resultid="1994" lane="5" heatid="6998" entrytime="00:04:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.75" />
                    <SPLIT distance="50" swimtime="00:00:57.11" />
                    <SPLIT distance="75" swimtime="00:01:28.75" />
                    <SPLIT distance="100" swimtime="00:02:01.14" />
                    <SPLIT distance="125" swimtime="00:02:33.82" />
                    <SPLIT distance="150" swimtime="00:03:07.22" />
                    <SPLIT distance="175" swimtime="00:03:40.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1581" points="133" reactiontime="+112" swimtime="00:04:11.25" resultid="1995" lane="3" heatid="7067" entrytime="00:04:24.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.32" />
                    <SPLIT distance="50" swimtime="00:00:57.74" />
                    <SPLIT distance="75" swimtime="00:01:30.60" />
                    <SPLIT distance="100" swimtime="00:02:04.13" />
                    <SPLIT distance="125" swimtime="00:02:39.11" />
                    <SPLIT distance="150" swimtime="00:03:14.33" />
                    <SPLIT distance="175" swimtime="00:03:43.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="83" reactiontime="+105" swimtime="00:00:58.23" resultid="1996" lane="4" heatid="7275" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="152" reactiontime="+101" swimtime="00:01:50.15" resultid="1991" lane="8" heatid="6724" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.40" />
                    <SPLIT distance="50" swimtime="00:00:51.08" />
                    <SPLIT distance="75" swimtime="00:01:23.00" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K 11" eventid="1222" reactiontime="+104" status="DSQ" swimtime="00:00:53.95" resultid="1992" lane="7" heatid="6849" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-01" firstname="Danuta" gender="F" lastname="Radkowiak" nation="POL" athleteid="1998">
              <RESULTS>
                <RESULT eventid="1679" points="227" reactiontime="+103" swimtime="00:01:46.60" resultid="2003" lane="8" heatid="7298" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.66" />
                    <SPLIT distance="50" swimtime="00:00:50.81" />
                    <SPLIT distance="75" swimtime="00:01:18.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1409" points="222" reactiontime="+100" swimtime="00:03:51.48" resultid="2001" lane="5" heatid="6999" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.48" />
                    <SPLIT distance="50" swimtime="00:00:52.76" />
                    <SPLIT distance="75" swimtime="00:01:22.11" />
                    <SPLIT distance="100" swimtime="00:01:51.16" />
                    <SPLIT distance="125" swimtime="00:02:21.12" />
                    <SPLIT distance="150" swimtime="00:02:51.88" />
                    <SPLIT distance="175" swimtime="00:03:21.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1781" points="160" reactiontime="+105" swimtime="00:08:15.87" resultid="2004" lane="3" heatid="7355" entrytime="00:08:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.21" />
                    <SPLIT distance="50" swimtime="00:00:54.73" />
                    <SPLIT distance="75" swimtime="00:01:25.08" />
                    <SPLIT distance="100" swimtime="00:01:56.75" />
                    <SPLIT distance="125" swimtime="00:02:32.98" />
                    <SPLIT distance="150" swimtime="00:03:06.69" />
                    <SPLIT distance="175" swimtime="00:03:39.51" />
                    <SPLIT distance="200" swimtime="00:04:13.43" />
                    <SPLIT distance="225" swimtime="00:04:45.82" />
                    <SPLIT distance="250" swimtime="00:05:18.12" />
                    <SPLIT distance="275" swimtime="00:05:50.79" />
                    <SPLIT distance="300" swimtime="00:06:23.33" />
                    <SPLIT distance="325" swimtime="00:06:52.40" />
                    <SPLIT distance="350" swimtime="00:07:20.42" />
                    <SPLIT distance="375" swimtime="00:07:48.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="135" reactiontime="+113" swimtime="00:04:01.59" resultid="2000" lane="3" heatid="6867" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.19" />
                    <SPLIT distance="50" swimtime="00:00:54.11" />
                    <SPLIT distance="75" swimtime="00:01:24.43" />
                    <SPLIT distance="100" swimtime="00:01:54.76" />
                    <SPLIT distance="125" swimtime="00:02:26.08" />
                    <SPLIT distance="150" swimtime="00:02:57.54" />
                    <SPLIT distance="175" swimtime="00:03:30.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1445" points="137" reactiontime="+96" swimtime="00:01:49.63" resultid="2002" lane="5" heatid="7012" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.19" />
                    <SPLIT distance="50" swimtime="00:00:51.84" />
                    <SPLIT distance="75" swimtime="00:01:21.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" status="DNS" swimtime="00:00:00.00" resultid="1999" lane="3" heatid="6850" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:56.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Leszek" gender="M" lastname="Kubicki" nation="POL" athleteid="2005">
              <RESULTS>
                <RESULT eventid="1375" points="285" reactiontime="+99" swimtime="00:05:34.32" resultid="2008" lane="8" heatid="6909" entrytime="00:04:46.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.33" />
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="75" swimtime="00:00:54.87" />
                    <SPLIT distance="100" swimtime="00:01:15.10" />
                    <SPLIT distance="125" swimtime="00:01:36.71" />
                    <SPLIT distance="150" swimtime="00:01:58.02" />
                    <SPLIT distance="175" swimtime="00:02:19.72" />
                    <SPLIT distance="200" swimtime="00:02:41.54" />
                    <SPLIT distance="225" swimtime="00:03:03.58" />
                    <SPLIT distance="250" swimtime="00:03:25.30" />
                    <SPLIT distance="275" swimtime="00:03:47.37" />
                    <SPLIT distance="300" swimtime="00:04:09.16" />
                    <SPLIT distance="325" swimtime="00:04:30.90" />
                    <SPLIT distance="350" swimtime="00:04:52.79" />
                    <SPLIT distance="375" swimtime="00:05:13.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="272" swimtime="00:22:29.27" resultid="2006" lane="3" heatid="6750" entrytime="00:23:18.00" />
                <RESULT eventid="1411" points="243" reactiontime="+99" swimtime="00:03:24.13" resultid="2009" lane="8" heatid="7007" entrytime="00:03:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.82" />
                    <SPLIT distance="50" swimtime="00:00:45.19" />
                    <SPLIT distance="75" swimtime="00:01:10.76" />
                    <SPLIT distance="100" swimtime="00:01:37.39" />
                    <SPLIT distance="125" swimtime="00:02:04.26" />
                    <SPLIT distance="150" swimtime="00:02:31.25" />
                    <SPLIT distance="175" swimtime="00:02:57.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="260" reactiontime="+99" swimtime="00:02:41.11" resultid="2010" lane="8" heatid="7060" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.02" />
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                    <SPLIT distance="75" swimtime="00:00:54.14" />
                    <SPLIT distance="100" swimtime="00:01:15.12" />
                    <SPLIT distance="125" swimtime="00:01:36.65" />
                    <SPLIT distance="150" swimtime="00:01:58.42" />
                    <SPLIT distance="175" swimtime="00:02:20.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="263" reactiontime="+102" swimtime="00:01:13.40" resultid="2007" lane="7" heatid="6835" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.39" />
                    <SPLIT distance="75" swimtime="00:00:54.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" status="DNS" swimtime="00:00:00.00" resultid="2011" lane="7" heatid="7306" entrytime="00:01:35.00" />
                <RESULT eventid="1764" reactiontime="+96" status="DNS" swimtime="00:00:00.00" resultid="2012" lane="2" heatid="7341" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-01-01" firstname="Hanka" gender="F" lastname="Kania" nation="POL" athleteid="2013">
              <RESULTS>
                <RESULT eventid="1409" points="187" reactiontime="+104" swimtime="00:04:05.06" resultid="2017" heatid="7001" entrytime="00:03:19.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.20" />
                    <SPLIT distance="50" swimtime="00:00:51.13" />
                    <SPLIT distance="75" swimtime="00:01:19.96" />
                    <SPLIT distance="100" swimtime="00:01:51.86" />
                    <SPLIT distance="125" swimtime="00:02:26.02" />
                    <SPLIT distance="150" swimtime="00:03:00.00" />
                    <SPLIT distance="175" swimtime="00:03:33.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="204" reactiontime="+93" swimtime="00:01:50.46" resultid="2020" lane="4" heatid="7297" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.55" />
                    <SPLIT distance="50" swimtime="00:00:52.67" />
                    <SPLIT distance="75" swimtime="00:01:21.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1445" points="135" reactiontime="+104" swimtime="00:01:50.10" resultid="2018" lane="3" heatid="7013" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.99" />
                    <SPLIT distance="50" swimtime="00:00:49.71" />
                    <SPLIT distance="75" swimtime="00:01:19.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="226" reactiontime="+90" swimtime="00:00:49.74" resultid="2016" lane="7" heatid="6850" entrytime="00:00:51.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="168" reactiontime="+109" swimtime="00:00:46.05" resultid="2019" lane="7" heatid="7277" entrytime="00:00:47.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="208" reactiontime="+109" swimtime="00:01:39.13" resultid="2014" lane="6" heatid="6725" entrytime="00:01:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.78" />
                    <SPLIT distance="50" swimtime="00:00:46.27" />
                    <SPLIT distance="75" swimtime="00:01:15.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="2015" lane="1" heatid="6824" entrytime="00:01:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1923-01-01" firstname="Danuta" gender="F" lastname="Kowalewska" nation="POL" athleteid="2021">
              <RESULTS>
                <RESULT eventid="1679" points="14" swimtime="00:04:24.81" resultid="2024" lane="3" heatid="7295" entrytime="00:04:00.77">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:01:06.36" />
                    <SPLIT distance="50" swimtime="00:02:17.07" />
                    <SPLIT distance="75" swimtime="00:03:26.51" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1409" points="13" swimtime="00:09:41.85" resultid="2023" lane="3" heatid="6997" entrytime="00:09:47.74">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:01:07.83" />
                    <SPLIT distance="50" swimtime="00:02:25.32" />
                    <SPLIT distance="75" swimtime="00:03:43.47" />
                    <SPLIT distance="100" swimtime="00:04:58.34" />
                    <SPLIT distance="125" swimtime="00:06:10.98" />
                    <SPLIT distance="150" swimtime="00:07:25.24" />
                    <SPLIT distance="175" swimtime="00:08:36.24" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1222" points="21" swimtime="00:01:48.37" resultid="2022" lane="8" heatid="6848" entrytime="00:01:49.32" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-01-01" firstname="Anna" gender="F" lastname="Walczak" nation="POL" athleteid="2025">
              <RESULTS>
                <RESULT eventid="1713" points="158" reactiontime="+69" swimtime="00:01:48.64" resultid="2029" lane="2" heatid="7314" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.64" />
                    <SPLIT distance="50" swimtime="00:00:54.05" />
                    <SPLIT distance="75" swimtime="00:01:22.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="131" reactiontime="+102" swimtime="00:01:43.97" resultid="2026" lane="7" heatid="6823" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.00" />
                    <SPLIT distance="50" swimtime="00:00:47.66" />
                    <SPLIT distance="75" swimtime="00:01:15.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="135" reactiontime="+102" swimtime="00:00:46.72" resultid="2028" lane="2" heatid="7329" entrytime="00:00:47.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="181" reactiontime="+65" swimtime="00:00:48.83" resultid="2027" lane="1" heatid="7027" entrytime="00:00:49.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Magdalena" gender="F" lastname="Majewska" nation="POL" athleteid="2030">
              <RESULTS>
                <RESULT eventid="1747" points="215" reactiontime="+102" swimtime="00:00:40.00" resultid="2032" lane="1" heatid="7330" entrytime="00:00:40.82">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="166" reactiontime="+63" swimtime="00:00:50.31" resultid="2031" lane="4" heatid="7027" entrytime="00:00:45.23">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1324" points="149" reactiontime="+66" swimtime="00:03:24.07" resultid="2034" lane="7" heatid="6979" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.79" />
                    <SPLIT distance="50" swimtime="00:00:49.31" />
                    <SPLIT distance="75" swimtime="00:01:17.11" />
                    <SPLIT distance="100" swimtime="00:01:10.24" />
                    <SPLIT distance="125" swimtime="00:02:14.49" />
                    <SPLIT distance="150" swimtime="00:01:48.61" />
                    <SPLIT distance="175" swimtime="00:03:04.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2025" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="1990" number="2" reactiontime="+69" />
                    <RELAYPOSITION athleteid="1984" number="3" />
                    <RELAYPOSITION athleteid="1971" number="4" reactiontime="+76" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="319" agemin="280" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1815" status="DNS" swimtime="00:00:00.00" resultid="2035" lane="8" heatid="7503" entrytime="00:04:00.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1984" number="1" />
                    <RELAYPOSITION athleteid="1979" number="2" />
                    <RELAYPOSITION athleteid="1922" number="3" />
                    <RELAYPOSITION athleteid="2025" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="GRKOZ" name="Grot Koziegłowy" nation="POL" region="WIE">
          <CONTACT name="JERSZYŃSKI" phone="500276047" />
          <ATHLETES>
            <ATHLETE birthdate="1975-08-24" firstname="Adam" gender="M" lastname="Witkowski" nation="POL" athleteid="2048">
              <RESULTS>
                <RESULT eventid="1075" points="220" swimtime="00:12:39.66" resultid="2049" lane="6" heatid="6719" entrytime="00:12:20.00" />
                <RESULT eventid="1375" points="244" reactiontime="+104" swimtime="00:05:52.15" resultid="2050" lane="6" heatid="6905" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.47" />
                    <SPLIT distance="50" swimtime="00:00:38.39" />
                    <SPLIT distance="75" swimtime="00:00:59.50" />
                    <SPLIT distance="100" swimtime="00:01:21.47" />
                    <SPLIT distance="125" swimtime="00:01:42.69" />
                    <SPLIT distance="150" swimtime="00:02:04.89" />
                    <SPLIT distance="175" swimtime="00:02:27.40" />
                    <SPLIT distance="200" swimtime="00:02:50.80" />
                    <SPLIT distance="225" swimtime="00:03:13.42" />
                    <SPLIT distance="250" swimtime="00:03:36.22" />
                    <SPLIT distance="275" swimtime="00:03:59.43" />
                    <SPLIT distance="300" swimtime="00:04:22.50" />
                    <SPLIT distance="325" swimtime="00:04:45.45" />
                    <SPLIT distance="350" swimtime="00:05:08.71" />
                    <SPLIT distance="375" swimtime="00:05:31.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TRCZE" name="UKS TRÓJKA Częstochowa" nation="POL" region="SLA">
          <CONTACT city="Częstochowa" email="trojkaczestochowa@poczta.onet.pl" name="Gawda Jacek" phone="511181791" state="ŚL" zip="42-200" />
          <ATHLETES>
            <ATHLETE birthdate="1990-02-15" firstname="Manuela" gender="F" lastname="Nawrocka" nation="POL" license="S00111100008" athleteid="2052">
              <RESULTS>
                <RESULT eventid="1581" points="482" reactiontime="+88" swimtime="00:02:43.76" resultid="2057" lane="3" heatid="7070" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.61" />
                    <SPLIT distance="50" swimtime="00:00:37.27" />
                    <SPLIT distance="75" swimtime="00:00:58.35" />
                    <SPLIT distance="100" swimtime="00:01:18.69" />
                    <SPLIT distance="125" swimtime="00:01:42.80" />
                    <SPLIT distance="150" swimtime="00:02:06.89" />
                    <SPLIT distance="175" swimtime="00:02:26.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="489" reactiontime="+93" swimtime="00:01:14.59" resultid="2053" lane="3" heatid="6729" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.89" />
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                    <SPLIT distance="75" swimtime="00:00:57.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="393" reactiontime="+84" swimtime="00:00:34.73" resultid="2058" heatid="7280" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="417" reactiontime="+85" swimtime="00:00:40.56" resultid="2055" heatid="6853" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="506" reactiontime="+85" swimtime="00:01:06.35" resultid="2054" lane="5" heatid="6828" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.10" />
                    <SPLIT distance="50" swimtime="00:00:31.39" />
                    <SPLIT distance="75" swimtime="00:00:48.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="489" reactiontime="+84" swimtime="00:00:30.42" resultid="2059" lane="7" heatid="7335" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="451" reactiontime="+76" swimtime="00:00:36.07" resultid="2056" lane="6" heatid="7031" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-09-11" firstname="Karolina" gender="F" lastname="Wawrzyńczak" nation="POL" license="S00111100007" athleteid="2060">
              <RESULTS>
                <RESULT eventid="1713" points="485" reactiontime="+74" swimtime="00:01:14.80" resultid="2064" lane="5" heatid="7317" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.82" />
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                    <SPLIT distance="75" swimtime="00:00:55.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="414" reactiontime="+75" swimtime="00:02:47.99" resultid="2061" lane="3" heatid="6879" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.23" />
                    <SPLIT distance="50" swimtime="00:00:38.33" />
                    <SPLIT distance="75" swimtime="00:00:58.75" />
                    <SPLIT distance="100" swimtime="00:01:20.05" />
                    <SPLIT distance="125" swimtime="00:01:41.82" />
                    <SPLIT distance="150" swimtime="00:02:04.21" />
                    <SPLIT distance="175" swimtime="00:02:26.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="477" reactiontime="+76" swimtime="00:00:35.39" resultid="2062" lane="5" heatid="7031" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="391" reactiontime="+90" swimtime="00:00:34.80" resultid="2063" lane="6" heatid="7280" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-07-31" firstname="Piotr" gender="M" lastname="Krogulec" nation="POL" license="S00111200006" athleteid="2065">
              <RESULTS>
                <RESULT eventid="1730" points="480" reactiontime="+72" swimtime="00:01:07.08" resultid="2072" lane="1" heatid="7325" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.36" />
                    <SPLIT distance="50" swimtime="00:00:32.06" />
                    <SPLIT distance="75" swimtime="00:00:49.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="503" reactiontime="+78" swimtime="00:00:30.75" resultid="2070" lane="4" heatid="7040" entrytime="00:00:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="484" reactiontime="+78" swimtime="00:01:04.16" resultid="2069" lane="5" heatid="7021" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.48" />
                    <SPLIT distance="50" swimtime="00:00:29.83" />
                    <SPLIT distance="75" swimtime="00:00:46.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="520" reactiontime="+81" swimtime="00:00:33.78" resultid="2068" heatid="6863" entrytime="00:00:36.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="461" reactiontime="+85" swimtime="00:01:06.18" resultid="2066" lane="1" heatid="6742" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.99" />
                    <SPLIT distance="50" swimtime="00:00:29.25" />
                    <SPLIT distance="75" swimtime="00:00:49.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="474" reactiontime="+89" swimtime="00:00:29.43" resultid="2071" lane="2" heatid="7288" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="499" reactiontime="+81" swimtime="00:00:59.28" resultid="2067" lane="4" heatid="6841" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.03" />
                    <SPLIT distance="50" swimtime="00:00:27.99" />
                    <SPLIT distance="75" swimtime="00:00:43.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-10-04" firstname="Jakub" gender="M" lastname="Kowalik" nation="POL" license="S00111200005" athleteid="2073">
              <RESULTS>
                <RESULT eventid="1564" points="424" reactiontime="+82" swimtime="00:02:17.02" resultid="2078" lane="8" heatid="7063" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.11" />
                    <SPLIT distance="50" swimtime="00:00:30.37" />
                    <SPLIT distance="75" swimtime="00:00:47.27" />
                    <SPLIT distance="100" swimtime="00:01:04.79" />
                    <SPLIT distance="125" swimtime="00:01:22.55" />
                    <SPLIT distance="150" swimtime="00:01:40.95" />
                    <SPLIT distance="175" swimtime="00:01:58.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="402" reactiontime="+80" swimtime="00:01:08.25" resultid="2077" lane="6" heatid="7021" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.86" />
                    <SPLIT distance="50" swimtime="00:00:30.37" />
                    <SPLIT distance="75" swimtime="00:00:48.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="437" reactiontime="+77" swimtime="00:00:35.80" resultid="2076" lane="7" heatid="6864" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="489" reactiontime="+79" swimtime="00:00:29.13" resultid="2079" lane="2" heatid="7290" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="513" reactiontime="+81" swimtime="00:00:58.76" resultid="2075" lane="5" heatid="6841" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.13" />
                    <SPLIT distance="50" swimtime="00:00:27.97" />
                    <SPLIT distance="75" swimtime="00:00:43.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="427" reactiontime="+83" swimtime="00:01:07.92" resultid="2074" lane="8" heatid="6743" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.26" />
                    <SPLIT distance="50" swimtime="00:00:30.85" />
                    <SPLIT distance="75" swimtime="00:00:52.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="527" reactiontime="+81" swimtime="00:00:26.33" resultid="2080" lane="5" heatid="7351" entrytime="00:00:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-12-08" firstname="Bartłomiej" gender="M" lastname="Drzewski" nation="POL" athleteid="2081">
              <RESULTS>
                <RESULT eventid="1239" points="401" reactiontime="+76" swimtime="00:00:36.83" resultid="2084" lane="5" heatid="6864" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="422" reactiontime="+70" swimtime="00:00:28.35" resultid="2088" lane="7" heatid="7351" entrytime="00:00:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="2083" lane="4" heatid="6840" entrytime="00:01:05.00" />
                <RESULT eventid="1496" status="DNS" swimtime="00:00:00.00" resultid="2085" lane="4" heatid="7039" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="2086" lane="4" heatid="7062" entrytime="00:02:22.00" />
                <RESULT eventid="1696" status="DNS" swimtime="00:00:00.00" resultid="2087" lane="5" heatid="7309" entrytime="00:01:20.00" />
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="2082" lane="5" heatid="6740" entrytime="00:01:12.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-11-28" firstname="Przemysław" gender="M" lastname="Szczypiński" nation="POL" license="S00111200010" athleteid="2089">
              <RESULTS>
                <RESULT eventid="1307" points="376" reactiontime="+70" swimtime="00:02:37.84" resultid="2091" heatid="6887" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.12" />
                    <SPLIT distance="50" swimtime="00:00:35.77" />
                    <SPLIT distance="75" swimtime="00:00:55.32" />
                    <SPLIT distance="100" swimtime="00:01:15.36" />
                    <SPLIT distance="125" swimtime="00:01:35.78" />
                    <SPLIT distance="150" swimtime="00:01:56.83" />
                    <SPLIT distance="175" swimtime="00:02:17.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="384" reactiontime="+71" swimtime="00:02:37.07" resultid="2093" lane="3" heatid="7079" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.98" />
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                    <SPLIT distance="75" swimtime="00:00:51.41" />
                    <SPLIT distance="100" swimtime="00:01:10.72" />
                    <SPLIT distance="125" swimtime="00:01:35.01" />
                    <SPLIT distance="150" swimtime="00:01:58.92" />
                    <SPLIT distance="175" swimtime="00:02:18.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="392" reactiontime="+71" swimtime="00:01:11.77" resultid="2094" lane="3" heatid="7325" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.57" />
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="75" swimtime="00:00:52.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="411" reactiontime="+73" swimtime="00:00:32.89" resultid="2092" lane="3" heatid="7041" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="369" reactiontime="+75" swimtime="00:01:11.28" resultid="2090" lane="6" heatid="6743" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.68" />
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                    <SPLIT distance="75" swimtime="00:00:53.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="96" agemin="80" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1177" points="518" reactiontime="+76" swimtime="00:01:48.02" resultid="2095" lane="7" heatid="6810" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.34" />
                    <SPLIT distance="50" swimtime="00:00:27.94" />
                    <SPLIT distance="75" swimtime="00:00:40.91" />
                    <SPLIT distance="100" swimtime="00:00:55.66" />
                    <SPLIT distance="125" swimtime="00:01:08.40" />
                    <SPLIT distance="150" swimtime="00:01:21.84" />
                    <SPLIT distance="175" swimtime="00:01:34.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2081" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="2089" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="2073" number="3" reactiontime="+81" />
                    <RELAYPOSITION athleteid="2065" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1341" points="449" reactiontime="+72" swimtime="00:02:04.71" resultid="2096" lane="4" heatid="6987" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.86" />
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                    <SPLIT distance="75" swimtime="00:00:49.37" />
                    <SPLIT distance="100" swimtime="00:01:07.54" />
                    <SPLIT distance="125" swimtime="00:01:20.88" />
                    <SPLIT distance="150" swimtime="00:01:36.61" />
                    <SPLIT distance="175" swimtime="00:01:49.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2089" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="2065" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="2073" number="3" reactiontime="+89" />
                    <RELAYPOSITION athleteid="2081" number="4" reactiontime="+67" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="96" agemin="80" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1615" status="DNS" swimtime="00:00:00.00" resultid="2097" lane="2" heatid="7443" entrytime="00:01:55.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2065" number="1" />
                    <RELAYPOSITION athleteid="2060" number="2" />
                    <RELAYPOSITION athleteid="2052" number="3" />
                    <RELAYPOSITION athleteid="2073" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1815" reactiontime="+74" swimtime="00:02:09.87" resultid="2098" lane="6" heatid="7504" entrytime="00:02:10.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.87" />
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                    <SPLIT distance="75" swimtime="00:00:51.13" />
                    <SPLIT distance="100" swimtime="00:01:09.25" />
                    <SPLIT distance="125" swimtime="00:01:22.53" />
                    <SPLIT distance="150" swimtime="00:01:38.21" />
                    <SPLIT distance="175" swimtime="00:01:53.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2060" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="2065" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="2073" number="3" reactiontime="+80" />
                    <RELAYPOSITION athleteid="2052" number="4" reactiontime="+85" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="KOKRA" name="Masters Korona Kraków" nation="POL">
          <CONTACT city="Kraków" email="masterskorona@wp.pl" internet="www.masterskorona.pl" name="Mariola Kuliś" phone="500677133" state="MAŁ" street="Kalwaryjska 9-15" zip="30-504" />
          <ATHLETES>
            <ATHLETE birthdate="1966-07-27" firstname="Mariola" gender="F" lastname="Kuliś" nation="POL" athleteid="2105">
              <RESULTS>
                <RESULT eventid="1092" points="452" reactiontime="+73" swimtime="00:01:16.59" resultid="2106" lane="1" heatid="6729" entrytime="00:01:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.30" />
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                    <SPLIT distance="75" swimtime="00:00:57.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="435" reactiontime="+77" swimtime="00:01:09.75" resultid="2107" lane="3" heatid="6827" entrytime="00:01:11.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.68" />
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                    <SPLIT distance="75" swimtime="00:00:51.29" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1222" points="493" reactiontime="+74" swimtime="00:00:38.36" resultid="2108" lane="6" heatid="6853" entrytime="00:00:39.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="438" reactiontime="+62" swimtime="00:00:36.41" resultid="2109" lane="4" heatid="7030" entrytime="00:00:36.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="447" reactiontime="+72" swimtime="00:00:31.33" resultid="2112" lane="8" heatid="7335" entrytime="00:00:30.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="361" reactiontime="+90" swimtime="00:02:41.13" resultid="2110" lane="5" heatid="7052" entrytime="00:02:41.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.06" />
                    <SPLIT distance="50" swimtime="00:00:36.04" />
                    <SPLIT distance="75" swimtime="00:00:55.84" />
                    <SPLIT distance="100" swimtime="00:01:16.29" />
                    <SPLIT distance="125" swimtime="00:01:37.33" />
                    <SPLIT distance="150" swimtime="00:01:58.58" />
                    <SPLIT distance="175" swimtime="00:02:20.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="403" reactiontime="+62" swimtime="00:01:19.55" resultid="2111" lane="6" heatid="7315" entrytime="00:01:37.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.06" />
                    <SPLIT distance="50" swimtime="00:00:38.72" />
                    <SPLIT distance="75" swimtime="00:00:59.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-07-26" firstname="Anna" gender="F" lastname="Kożmin" nation="POL" athleteid="2113">
              <RESULTS>
                <RESULT eventid="1222" points="193" reactiontime="+114" swimtime="00:00:52.36" resultid="2115" lane="1" heatid="6849" entrytime="00:00:54.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="168" reactiontime="+115" swimtime="00:01:57.73" resultid="2117" lane="1" heatid="7297" entrytime="00:01:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.19" />
                    <SPLIT distance="50" swimtime="00:00:55.19" />
                    <SPLIT distance="75" swimtime="00:01:26.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1409" points="151" reactiontime="+116" swimtime="00:04:22.96" resultid="2116" lane="3" heatid="6998" entrytime="00:04:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.22" />
                    <SPLIT distance="50" swimtime="00:00:55.96" />
                    <SPLIT distance="75" swimtime="00:01:29.11" />
                    <SPLIT distance="100" swimtime="00:02:03.86" />
                    <SPLIT distance="125" swimtime="00:02:39.46" />
                    <SPLIT distance="150" swimtime="00:03:14.31" />
                    <SPLIT distance="175" swimtime="00:03:48.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="133" reactiontime="+115" swimtime="00:01:54.93" resultid="2114" lane="3" heatid="6724" entrytime="00:01:53.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.51" />
                    <SPLIT distance="50" swimtime="00:00:55.02" />
                    <SPLIT distance="75" swimtime="00:01:26.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-09-12" firstname="Joanna" gender="F" lastname="Kwatera" nation="POL" athleteid="2118">
              <RESULTS>
                <RESULT eventid="1679" points="332" reactiontime="+73" swimtime="00:01:33.94" resultid="2122" lane="4" heatid="7299" entrytime="00:01:34.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.93" />
                    <SPLIT distance="50" swimtime="00:00:44.67" />
                    <SPLIT distance="75" swimtime="00:01:09.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1409" points="362" reactiontime="+84" swimtime="00:03:16.68" resultid="2121" lane="8" heatid="7001" entrytime="00:03:19.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.78" />
                    <SPLIT distance="50" swimtime="00:00:44.32" />
                    <SPLIT distance="75" swimtime="00:01:08.57" />
                    <SPLIT distance="100" swimtime="00:01:33.33" />
                    <SPLIT distance="125" swimtime="00:01:58.89" />
                    <SPLIT distance="150" swimtime="00:02:24.83" />
                    <SPLIT distance="175" swimtime="00:02:51.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="353" reactiontime="+84" swimtime="00:00:42.88" resultid="2120" lane="1" heatid="6852" entrytime="00:00:42.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="245" reactiontime="+86" swimtime="00:01:33.92" resultid="2119" lane="6" heatid="6726" entrytime="00:01:34.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.15" />
                    <SPLIT distance="50" swimtime="00:00:46.77" />
                    <SPLIT distance="75" swimtime="00:01:11.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-09-15" firstname="Mirosława" gender="F" lastname="Legutko" nation="POL" athleteid="2123">
              <RESULTS>
                <RESULT eventid="1781" points="211" reactiontime="+113" swimtime="00:07:32.52" resultid="2130" lane="7" heatid="7356" entrytime="00:07:50.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.42" />
                    <SPLIT distance="50" swimtime="00:00:50.30" />
                    <SPLIT distance="75" swimtime="00:01:19.76" />
                    <SPLIT distance="100" swimtime="00:01:49.79" />
                    <SPLIT distance="125" swimtime="00:02:18.05" />
                    <SPLIT distance="150" swimtime="00:02:46.44" />
                    <SPLIT distance="175" swimtime="00:03:15.79" />
                    <SPLIT distance="200" swimtime="00:03:44.28" />
                    <SPLIT distance="225" swimtime="00:04:17.45" />
                    <SPLIT distance="250" swimtime="00:04:49.80" />
                    <SPLIT distance="275" swimtime="00:05:21.90" />
                    <SPLIT distance="300" swimtime="00:05:54.91" />
                    <SPLIT distance="325" swimtime="00:06:20.16" />
                    <SPLIT distance="350" swimtime="00:06:44.80" />
                    <SPLIT distance="375" swimtime="00:07:09.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1581" points="225" reactiontime="+108" swimtime="00:03:31.10" resultid="2128" lane="7" heatid="7069" entrytime="00:03:30.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.86" />
                    <SPLIT distance="50" swimtime="00:00:46.63" />
                    <SPLIT distance="75" swimtime="00:02:10.95" />
                    <SPLIT distance="100" swimtime="00:01:38.71" />
                    <SPLIT distance="125" swimtime="00:03:08.17" />
                    <SPLIT distance="150" swimtime="00:02:43.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="163" reactiontime="+107" swimtime="00:03:47.28" resultid="2125" lane="1" heatid="6868" entrytime="00:03:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.42" />
                    <SPLIT distance="50" swimtime="00:00:47.29" />
                    <SPLIT distance="75" swimtime="00:01:16.50" />
                    <SPLIT distance="100" swimtime="00:01:46.58" />
                    <SPLIT distance="125" swimtime="00:02:16.65" />
                    <SPLIT distance="150" swimtime="00:02:47.32" />
                    <SPLIT distance="175" swimtime="00:03:17.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="205" reactiontime="+83" swimtime="00:03:32.29" resultid="2126" lane="3" heatid="6877" entrytime="00:03:30.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:01:16.16" />
                    <SPLIT distance="50" swimtime="00:00:50.27" />
                    <SPLIT distance="75" swimtime="00:02:12.43" />
                    <SPLIT distance="100" swimtime="00:01:43.73" />
                    <SPLIT distance="125" swimtime="00:03:07.17" />
                    <SPLIT distance="150" swimtime="00:02:40.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1445" points="175" reactiontime="+106" swimtime="00:01:41.15" resultid="2127" lane="6" heatid="7013" entrytime="00:01:43.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.94" />
                    <SPLIT distance="50" swimtime="00:00:45.04" />
                    <SPLIT distance="75" swimtime="00:01:12.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="255" reactiontime="+103" swimtime="00:01:32.64" resultid="2124" heatid="6726" entrytime="00:01:36.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.82" />
                    <SPLIT distance="50" swimtime="00:00:41.10" />
                    <SPLIT distance="75" swimtime="00:01:09.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="239" reactiontime="+104" swimtime="00:00:40.98" resultid="2129" lane="5" heatid="7277" entrytime="00:00:43.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-04-22" firstname="Alicja" gender="F" lastname="Romańska" nation="POL" athleteid="2131">
              <RESULTS>
                <RESULT eventid="1547" points="150" reactiontime="+111" swimtime="00:03:36.07" resultid="2134" lane="1" heatid="7050" entrytime="00:03:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.48" />
                    <SPLIT distance="50" swimtime="00:00:49.47" />
                    <SPLIT distance="75" swimtime="00:01:15.53" />
                    <SPLIT distance="100" swimtime="00:01:43.90" />
                    <SPLIT distance="125" swimtime="00:02:12.44" />
                    <SPLIT distance="150" swimtime="00:02:41.35" />
                    <SPLIT distance="175" swimtime="00:03:09.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="140" reactiontime="+106" swimtime="00:01:41.62" resultid="2133" lane="4" heatid="6823" entrytime="00:01:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.77" />
                    <SPLIT distance="50" swimtime="00:00:49.94" />
                    <SPLIT distance="75" swimtime="00:01:16.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="145" swimtime="00:00:45.62" resultid="2136" heatid="7330" entrytime="00:00:42.00" entrycourse="SCM" />
                <RESULT comment="Z 2" eventid="1092" reactiontime="+105" status="DSQ" swimtime="00:00:00.00" resultid="2132" lane="7" heatid="6725" entrytime="00:01:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.46" />
                    <SPLIT distance="50" swimtime="00:00:56.81" />
                    <SPLIT distance="75" swimtime="00:01:32.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" status="DNS" swimtime="00:00:00.00" resultid="2135" lane="2" heatid="7276" entrytime="00:00:50.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-04-20" firstname="Małgorzata" gender="F" lastname="Szczygielska- Wertepna" nation="POL" athleteid="2137">
              <RESULTS>
                <RESULT eventid="1679" points="192" reactiontime="+88" swimtime="00:01:52.66" resultid="2139" lane="5" heatid="7297" entrytime="00:01:51.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.58" />
                    <SPLIT distance="50" swimtime="00:00:53.81" />
                    <SPLIT distance="75" swimtime="00:01:23.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="195" reactiontime="+88" swimtime="00:00:52.21" resultid="2138" lane="1" heatid="6850" entrytime="00:00:51.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-05-28" firstname="Marta" gender="F" lastname="Wolska" nation="POL" athleteid="2140">
              <RESULTS>
                <RESULT eventid="1290" points="104" reactiontime="+75" swimtime="00:04:25.89" resultid="2142" lane="2" heatid="6876" entrytime="00:04:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.27" />
                    <SPLIT distance="50" swimtime="00:01:01.09" />
                    <SPLIT distance="75" swimtime="00:01:34.72" />
                    <SPLIT distance="100" swimtime="00:02:09.06" />
                    <SPLIT distance="125" swimtime="00:02:44.87" />
                    <SPLIT distance="150" swimtime="00:03:19.57" />
                    <SPLIT distance="175" swimtime="00:03:52.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="130" reactiontime="+70" swimtime="00:00:54.54" resultid="2144" lane="8" heatid="7027" entrytime="00:00:53.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="109" swimtime="00:02:02.67" resultid="2146" lane="4" heatid="7313" entrytime="00:02:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.28" />
                    <SPLIT distance="75" swimtime="00:01:30.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" status="DNS" swimtime="00:00:00.00" resultid="2141" lane="2" heatid="6848" entrytime="00:01:00.00" entrycourse="SCM" />
                <RESULT eventid="1409" status="DNS" swimtime="00:00:00.00" resultid="2143" lane="6" heatid="6998" entrytime="00:04:40.00" entrycourse="SCM" />
                <RESULT eventid="1679" status="DNS" swimtime="00:00:00.00" resultid="2145" heatid="7296" entrytime="00:02:28.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-26" firstname="Marta" gender="F" lastname="Wysocka" nation="POL" athleteid="2147">
              <RESULTS>
                <RESULT eventid="1409" points="384" reactiontime="+86" swimtime="00:03:12.88" resultid="2151" lane="7" heatid="7001" entrytime="00:03:14.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.72" />
                    <SPLIT distance="50" swimtime="00:00:43.25" />
                    <SPLIT distance="75" swimtime="00:01:07.45" />
                    <SPLIT distance="100" swimtime="00:01:31.53" />
                    <SPLIT distance="125" swimtime="00:01:56.46" />
                    <SPLIT distance="150" swimtime="00:02:21.82" />
                    <SPLIT distance="175" swimtime="00:02:47.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="385" reactiontime="+91" swimtime="00:01:29.44" resultid="2153" lane="7" heatid="7300" entrytime="00:01:30.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.89" />
                    <SPLIT distance="50" swimtime="00:00:42.68" />
                    <SPLIT distance="75" swimtime="00:01:06.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="399" reactiontime="+88" swimtime="00:00:41.17" resultid="2150" lane="4" heatid="6852" entrytime="00:00:40.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="310" swimtime="00:01:26.84" resultid="2148" lane="2" heatid="6727" entrytime="00:01:26.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.49" />
                    <SPLIT distance="50" swimtime="00:00:43.64" />
                    <SPLIT distance="75" swimtime="00:01:06.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="311" reactiontime="+89" swimtime="00:01:17.97" resultid="2149" lane="2" heatid="6826" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.37" />
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                    <SPLIT distance="75" swimtime="00:00:57.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="267" reactiontime="+79" swimtime="00:00:42.95" resultid="2152" heatid="7029" entrytime="00:00:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="314" reactiontime="+87" swimtime="00:00:35.24" resultid="2154" lane="7" heatid="7333" entrytime="00:00:34.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-21" firstname="Klaudia" gender="F" lastname="Wysocka" nation="POL" athleteid="2155">
              <RESULTS>
                <RESULT eventid="1747" points="365" reactiontime="+86" swimtime="00:00:33.54" resultid="2162" lane="5" heatid="7333" entrytime="00:00:33.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="403" reactiontime="+88" swimtime="00:01:19.58" resultid="2156" lane="6" heatid="6728" entrytime="00:01:22.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.13" />
                    <SPLIT distance="50" swimtime="00:00:37.46" />
                    <SPLIT distance="75" swimtime="00:01:00.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="373" reactiontime="+91" swimtime="00:01:13.40" resultid="2157" lane="4" heatid="6826" entrytime="00:01:14.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.43" />
                    <SPLIT distance="50" swimtime="00:00:36.04" />
                    <SPLIT distance="75" swimtime="00:00:55.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1445" points="388" reactiontime="+92" swimtime="00:01:17.61" resultid="2159" lane="2" heatid="7014" entrytime="00:01:16.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.66" />
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                    <SPLIT distance="75" swimtime="00:00:56.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="408" reactiontime="+86" swimtime="00:00:34.32" resultid="2161" lane="2" heatid="7280" entrytime="00:00:33.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="362" reactiontime="+98" swimtime="00:05:38.71" resultid="2158" lane="3" heatid="6897" entrytime="00:05:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.47" />
                    <SPLIT distance="50" swimtime="00:00:38.70" />
                    <SPLIT distance="75" swimtime="00:00:59.17" />
                    <SPLIT distance="100" swimtime="00:01:19.92" />
                    <SPLIT distance="125" swimtime="00:01:40.89" />
                    <SPLIT distance="150" swimtime="00:02:02.21" />
                    <SPLIT distance="175" swimtime="00:02:23.49" />
                    <SPLIT distance="200" swimtime="00:02:45.43" />
                    <SPLIT distance="225" swimtime="00:03:06.91" />
                    <SPLIT distance="250" swimtime="00:03:28.34" />
                    <SPLIT distance="275" swimtime="00:03:50.13" />
                    <SPLIT distance="300" swimtime="00:04:12.17" />
                    <SPLIT distance="325" swimtime="00:04:34.20" />
                    <SPLIT distance="350" swimtime="00:04:56.01" />
                    <SPLIT distance="375" swimtime="00:05:18.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="359" reactiontime="+96" swimtime="00:02:41.52" resultid="2160" lane="2" heatid="7052" entrytime="00:02:42.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.12" />
                    <SPLIT distance="50" swimtime="00:00:37.95" />
                    <SPLIT distance="75" swimtime="00:00:57.87" />
                    <SPLIT distance="100" swimtime="00:01:18.24" />
                    <SPLIT distance="125" swimtime="00:01:39.29" />
                    <SPLIT distance="150" swimtime="00:02:00.42" />
                    <SPLIT distance="175" swimtime="00:02:21.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-12-23" firstname="Anna" gender="F" lastname="Janeczko" nation="POL" athleteid="2163">
              <RESULTS>
                <RESULT eventid="1290" points="252" reactiontime="+92" swimtime="00:03:18.06" resultid="2165" lane="7" heatid="6878" entrytime="00:03:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.47" />
                    <SPLIT distance="50" swimtime="00:00:44.52" />
                    <SPLIT distance="75" swimtime="00:01:08.88" />
                    <SPLIT distance="100" swimtime="00:01:33.98" />
                    <SPLIT distance="125" swimtime="00:02:00.77" />
                    <SPLIT distance="150" swimtime="00:02:28.06" />
                    <SPLIT distance="175" swimtime="00:02:53.84" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1126" points="225" swimtime="00:25:47.97" resultid="2164" lane="7" heatid="6747" entrytime="00:26:30.00" entrycourse="SCM" />
                <RESULT eventid="1581" points="255" reactiontime="+103" swimtime="00:03:22.39" resultid="2168" lane="2" heatid="7069" entrytime="00:03:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.79" />
                    <SPLIT distance="50" swimtime="00:00:48.64" />
                    <SPLIT distance="75" swimtime="00:01:14.84" />
                    <SPLIT distance="100" swimtime="00:01:40.46" />
                    <SPLIT distance="125" swimtime="00:02:09.95" />
                    <SPLIT distance="150" swimtime="00:02:38.84" />
                    <SPLIT distance="175" swimtime="00:03:02.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="284" reactiontime="+84" swimtime="00:01:29.39" resultid="2169" lane="7" heatid="7315" entrytime="00:01:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.45" />
                    <SPLIT distance="50" swimtime="00:00:43.78" />
                    <SPLIT distance="75" swimtime="00:01:06.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1781" points="228" reactiontime="+102" swimtime="00:07:20.55" resultid="2170" lane="8" heatid="7356" entrytime="00:07:58.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.55" />
                    <SPLIT distance="50" swimtime="00:00:55.12" />
                    <SPLIT distance="75" swimtime="00:01:26.87" />
                    <SPLIT distance="100" swimtime="00:02:00.11" />
                    <SPLIT distance="125" swimtime="00:02:27.54" />
                    <SPLIT distance="150" swimtime="00:02:54.43" />
                    <SPLIT distance="175" swimtime="00:03:21.15" />
                    <SPLIT distance="200" swimtime="00:03:47.10" />
                    <SPLIT distance="225" swimtime="00:04:17.64" />
                    <SPLIT distance="250" swimtime="00:04:47.99" />
                    <SPLIT distance="275" swimtime="00:05:17.64" />
                    <SPLIT distance="300" swimtime="00:05:47.38" />
                    <SPLIT distance="325" swimtime="00:06:12.53" />
                    <SPLIT distance="350" swimtime="00:06:36.09" />
                    <SPLIT distance="375" swimtime="00:06:59.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="244" reactiontime="+115" swimtime="00:06:26.24" resultid="2166" lane="2" heatid="6896" entrytime="00:06:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.42" />
                    <SPLIT distance="50" swimtime="00:00:43.08" />
                    <SPLIT distance="75" swimtime="00:01:05.93" />
                    <SPLIT distance="100" swimtime="00:01:30.03" />
                    <SPLIT distance="125" swimtime="00:01:53.88" />
                    <SPLIT distance="150" swimtime="00:02:19.09" />
                    <SPLIT distance="175" swimtime="00:02:43.33" />
                    <SPLIT distance="200" swimtime="00:03:08.84" />
                    <SPLIT distance="225" swimtime="00:03:33.66" />
                    <SPLIT distance="250" swimtime="00:03:59.31" />
                    <SPLIT distance="275" swimtime="00:04:24.10" />
                    <SPLIT distance="300" swimtime="00:04:50.11" />
                    <SPLIT distance="325" swimtime="00:05:14.84" />
                    <SPLIT distance="350" swimtime="00:05:39.78" />
                    <SPLIT distance="375" swimtime="00:06:03.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="286" reactiontime="+82" swimtime="00:00:41.96" resultid="2167" lane="6" heatid="7027" entrytime="00:00:49.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-03-07" firstname="Robert" gender="M" lastname="Grela" nation="POL" athleteid="2171">
              <RESULTS>
                <RESULT eventid="1273" points="311" reactiontime="+78" swimtime="00:02:45.22" resultid="2172" heatid="6874" entrytime="00:02:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.89" />
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                    <SPLIT distance="75" swimtime="00:00:50.45" />
                    <SPLIT distance="100" swimtime="00:01:09.60" />
                    <SPLIT distance="125" swimtime="00:01:29.39" />
                    <SPLIT distance="150" swimtime="00:01:51.64" />
                    <SPLIT distance="175" swimtime="00:02:17.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="405" reactiontime="+76" swimtime="00:01:08.10" resultid="2173" lane="6" heatid="7022" entrytime="00:01:07.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.66" />
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                    <SPLIT distance="75" swimtime="00:00:49.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="454" reactiontime="+71" swimtime="00:00:29.86" resultid="2174" lane="2" heatid="7292" entrytime="00:00:28.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-03-15" firstname="Mariusz" gender="M" lastname="Kaliszyk" nation="POL" athleteid="2180">
              <RESULTS>
                <RESULT eventid="1496" points="472" reactiontime="+59" swimtime="00:00:31.42" resultid="2182" heatid="7039" entrytime="00:00:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="515" reactiontime="+78" swimtime="00:00:26.54" resultid="2183" lane="7" heatid="7344" entrytime="00:00:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="469" reactiontime="+84" swimtime="00:01:00.52" resultid="2181" lane="7" heatid="6840" entrytime="00:01:06.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.60" />
                    <SPLIT distance="50" swimtime="00:00:28.96" />
                    <SPLIT distance="75" swimtime="00:00:44.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-11-02" firstname="Piotr" gender="M" lastname="Klimczak" nation="POL" athleteid="2184">
              <RESULTS>
                <RESULT eventid="1205" points="293" reactiontime="+94" swimtime="00:01:10.77" resultid="2185" lane="7" heatid="6837" entrytime="00:01:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.92" />
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                    <SPLIT distance="75" swimtime="00:00:51.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-08-16" firstname="Marek" gender="M" lastname="Nawieśniak" nation="POL" athleteid="2186">
              <RESULTS>
                <RESULT eventid="1109" points="260" reactiontime="+74" swimtime="00:01:20.07" resultid="2187" lane="6" heatid="6736" entrytime="00:01:22.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.97" />
                    <SPLIT distance="50" swimtime="00:00:36.69" />
                    <SPLIT distance="75" swimtime="00:01:01.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="265" reactiontime="+89" swimtime="00:00:35.74" resultid="2190" lane="6" heatid="7287" entrytime="00:00:33.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="260" reactiontime="+70" swimtime="00:02:41.18" resultid="2189" lane="4" heatid="7059" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.81" />
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                    <SPLIT distance="75" swimtime="00:00:55.50" />
                    <SPLIT distance="100" swimtime="00:01:15.84" />
                    <SPLIT distance="125" swimtime="00:01:36.45" />
                    <SPLIT distance="150" swimtime="00:01:58.14" />
                    <SPLIT distance="175" swimtime="00:02:19.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="370" reactiontime="+94" swimtime="00:00:29.63" resultid="2191" lane="1" heatid="7344" entrytime="00:00:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="329" reactiontime="+69" swimtime="00:01:08.11" resultid="2188" lane="8" heatid="6837" entrytime="00:01:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.45" />
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                    <SPLIT distance="75" swimtime="00:00:48.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-11-10" firstname="Waldemar" gender="M" lastname="Piszczek" nation="POL" athleteid="2192">
              <RESULTS>
                <RESULT eventid="1462" points="314" reactiontime="+92" swimtime="00:01:14.13" resultid="2196" lane="5" heatid="7020" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.61" />
                    <SPLIT distance="50" swimtime="00:00:32.73" />
                    <SPLIT distance="75" swimtime="00:00:52.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="304" reactiontime="+88" swimtime="00:02:49.38" resultid="2195" lane="3" heatid="6885" entrytime="00:02:47.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.34" />
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                    <SPLIT distance="75" swimtime="00:00:59.06" />
                    <SPLIT distance="100" swimtime="00:01:20.90" />
                    <SPLIT distance="125" swimtime="00:01:42.74" />
                    <SPLIT distance="150" swimtime="00:02:05.64" />
                    <SPLIT distance="175" swimtime="00:02:28.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="401" reactiontime="+99" swimtime="00:00:31.13" resultid="2198" lane="8" heatid="7290" entrytime="00:00:31.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="334" reactiontime="+77" swimtime="00:00:35.24" resultid="2197" heatid="7040" entrytime="00:00:34.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="329" reactiontime="+91" swimtime="00:01:14.02" resultid="2193" lane="7" heatid="6740" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.13" />
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                    <SPLIT distance="75" swimtime="00:00:55.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="396" reactiontime="+95" swimtime="00:00:37.01" resultid="2194" lane="1" heatid="6859" entrytime="00:00:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" status="DNS" swimtime="00:00:00.00" resultid="2199" lane="6" heatid="7324" entrytime="00:01:15.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-04-22" firstname="Szymon" gender="M" lastname="Pyrć" nation="POL" athleteid="2200">
              <RESULTS>
                <RESULT eventid="1143" points="383" swimtime="00:20:04.18" resultid="2201" lane="2" heatid="6751" entrytime="00:22:22.00" entrycourse="SCM" />
                <RESULT eventid="1273" points="413" reactiontime="+79" swimtime="00:02:30.36" resultid="2202" lane="7" heatid="6874" entrytime="00:02:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.79" />
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                    <SPLIT distance="75" swimtime="00:00:51.47" />
                    <SPLIT distance="100" swimtime="00:01:10.74" />
                    <SPLIT distance="125" swimtime="00:01:30.55" />
                    <SPLIT distance="150" swimtime="00:01:50.32" />
                    <SPLIT distance="175" swimtime="00:02:10.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="380" reactiontime="+76" swimtime="00:05:36.39" resultid="2205" heatid="7363" entrytime="00:06:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.77" />
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                    <SPLIT distance="75" swimtime="00:00:50.90" />
                    <SPLIT distance="100" swimtime="00:01:10.14" />
                    <SPLIT distance="125" swimtime="00:01:34.51" />
                    <SPLIT distance="150" swimtime="00:01:57.73" />
                    <SPLIT distance="175" swimtime="00:02:19.95" />
                    <SPLIT distance="200" swimtime="00:02:42.46" />
                    <SPLIT distance="225" swimtime="00:03:06.86" />
                    <SPLIT distance="250" swimtime="00:03:31.90" />
                    <SPLIT distance="275" swimtime="00:03:56.61" />
                    <SPLIT distance="300" swimtime="00:04:21.40" />
                    <SPLIT distance="325" swimtime="00:04:40.99" />
                    <SPLIT distance="350" swimtime="00:04:59.93" />
                    <SPLIT distance="375" swimtime="00:05:18.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="421" reactiontime="+76" swimtime="00:01:07.20" resultid="2203" lane="4" heatid="7021" entrytime="00:01:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.55" />
                    <SPLIT distance="50" swimtime="00:00:31.39" />
                    <SPLIT distance="75" swimtime="00:00:49.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="409" reactiontime="+77" swimtime="00:00:30.91" resultid="2204" lane="5" heatid="7290" entrytime="00:00:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-07-17" firstname="Robert" gender="M" lastname="Rospondek" nation="POL" athleteid="2206">
              <RESULTS>
                <RESULT eventid="1764" points="220" reactiontime="+89" swimtime="00:00:35.25" resultid="2208" heatid="7343" entrytime="00:00:31.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="197" reactiontime="+102" swimtime="00:01:20.84" resultid="2207" lane="2" heatid="6839" entrytime="00:01:07.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.36" />
                    <SPLIT distance="50" swimtime="00:00:37.50" />
                    <SPLIT distance="75" swimtime="00:00:59.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-10-23" firstname="Wojciech" gender="M" lastname="Superson" nation="POL" athleteid="2209">
              <RESULTS>
                <RESULT eventid="1375" points="210" reactiontime="+112" swimtime="00:06:10.14" resultid="2211" heatid="6902" entrytime="00:06:28.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.43" />
                    <SPLIT distance="50" swimtime="00:00:43.25" />
                    <SPLIT distance="75" swimtime="00:01:06.17" />
                    <SPLIT distance="100" swimtime="00:02:16.07" />
                    <SPLIT distance="125" swimtime="00:01:52.55" />
                    <SPLIT distance="150" swimtime="00:03:50.39" />
                    <SPLIT distance="175" swimtime="00:03:26.24" />
                    <SPLIT distance="200" swimtime="00:04:36.67" />
                    <SPLIT distance="225" swimtime="00:04:13.35" />
                    <SPLIT distance="250" swimtime="00:05:23.41" />
                    <SPLIT distance="275" swimtime="00:04:59.65" />
                    <SPLIT distance="300" swimtime="00:06:10.14" />
                    <SPLIT distance="325" swimtime="00:05:46.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="209" reactiontime="+109" swimtime="00:02:53.43" resultid="2212" lane="2" heatid="7057" entrytime="00:02:57.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.16" />
                    <SPLIT distance="50" swimtime="00:00:40.56" />
                    <SPLIT distance="75" swimtime="00:01:02.51" />
                    <SPLIT distance="100" swimtime="00:01:24.66" />
                    <SPLIT distance="125" swimtime="00:01:47.80" />
                    <SPLIT distance="150" swimtime="00:02:09.97" />
                    <SPLIT distance="175" swimtime="00:02:32.68" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="przekroczony limit 24:30:00" eventid="1143" status="DSQ" swimtime="00:24:51.81" resultid="2210" lane="1" heatid="6750" entrytime="00:24:17.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-21" firstname="Wojciech" gender="M" lastname="Wolski" nation="POL" athleteid="2213">
              <RESULTS>
                <RESULT eventid="1109" points="256" reactiontime="+92" swimtime="00:01:20.51" resultid="2214" lane="7" heatid="6737" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.32" />
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                    <SPLIT distance="75" swimtime="00:01:01.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="193" reactiontime="+122" swimtime="00:00:47.01" resultid="2215" lane="1" heatid="6861" entrytime="00:00:37.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" status="DNS" swimtime="00:00:00.00" resultid="2220" heatid="7361" entrytime="00:06:50.00" entrycourse="SCM" />
                <RESULT eventid="1307" status="DNS" swimtime="00:00:00.00" resultid="2216" lane="8" heatid="6884" entrytime="00:03:20.00" entrycourse="SCM" />
                <RESULT eventid="1411" status="DNS" swimtime="00:00:00.00" resultid="2217" heatid="7009" entrytime="00:03:09.20" entrycourse="SCM" />
                <RESULT eventid="1598" status="DNS" swimtime="00:00:00.00" resultid="2218" lane="3" heatid="7071" />
                <RESULT eventid="1696" status="DNS" swimtime="00:00:00.00" resultid="2219" lane="1" heatid="7308" entrytime="00:01:25.25" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-07-17" firstname="Wojciech" gender="M" lastname="Liszkowski" nation="POL" athleteid="2221">
              <RESULTS>
                <RESULT eventid="1645" points="459" reactiontime="+73" swimtime="00:00:29.75" resultid="2226" lane="6" heatid="7291" entrytime="00:00:29.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="350" reactiontime="+83" swimtime="00:02:42.03" resultid="2225" lane="5" heatid="7078" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.17" />
                    <SPLIT distance="50" swimtime="00:00:31.28" />
                    <SPLIT distance="75" swimtime="00:00:52.43" />
                    <SPLIT distance="100" swimtime="00:01:12.92" />
                    <SPLIT distance="125" swimtime="00:01:36.96" />
                    <SPLIT distance="150" swimtime="00:02:01.24" />
                    <SPLIT distance="175" swimtime="00:02:22.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="406" reactiontime="+65" swimtime="00:00:33.03" resultid="2224" lane="2" heatid="7040" entrytime="00:00:33.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="437" reactiontime="+84" swimtime="00:00:35.80" resultid="2223" lane="6" heatid="6864" entrytime="00:00:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="351" reactiontime="+82" swimtime="00:01:12.51" resultid="2222" lane="7" heatid="6739" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.83" />
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                    <SPLIT distance="75" swimtime="00:00:54.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="2227" lane="5" heatid="7347" entrytime="00:00:28.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-03-21" firstname="Janusz" gender="M" lastname="Gołębiewski" nation="POL" athleteid="2228">
              <RESULTS>
                <RESULT eventid="1239" points="59" swimtime="00:01:09.72" resultid="2229" lane="6" heatid="6854" entrytime="00:01:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="30" swimtime="00:06:50.31" resultid="2230" lane="3" heatid="7002" entrytime="00:04:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:44.25" />
                    <SPLIT distance="50" swimtime="00:01:33.00" />
                    <SPLIT distance="75" swimtime="00:02:25.73" />
                    <SPLIT distance="100" swimtime="00:03:19.10" />
                    <SPLIT distance="125" swimtime="00:04:11.86" />
                    <SPLIT distance="150" swimtime="00:05:08.25" />
                    <SPLIT distance="175" swimtime="00:06:00.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" status="DNS" swimtime="00:00:00.00" resultid="2231" lane="1" heatid="7302" entrytime="00:02:15.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-27" firstname="Wacław" gender="M" lastname="Brożek" nation="POL" athleteid="2232">
              <RESULTS>
                <RESULT eventid="1598" points="153" reactiontime="+116" swimtime="00:03:33.53" resultid="2235" lane="4" heatid="7073" entrytime="00:03:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.14" />
                    <SPLIT distance="50" swimtime="00:00:40.48" />
                    <SPLIT distance="75" swimtime="00:01:10.49" />
                    <SPLIT distance="100" swimtime="00:01:41.25" />
                    <SPLIT distance="125" swimtime="00:02:13.53" />
                    <SPLIT distance="150" swimtime="00:02:47.20" />
                    <SPLIT distance="175" swimtime="00:03:10.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="178" reactiontime="+108" swimtime="00:06:31.05" resultid="2234" lane="3" heatid="6901" entrytime="00:06:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.66" />
                    <SPLIT distance="50" swimtime="00:00:38.24" />
                    <SPLIT distance="75" swimtime="00:01:00.16" />
                    <SPLIT distance="100" swimtime="00:01:23.21" />
                    <SPLIT distance="125" swimtime="00:01:47.00" />
                    <SPLIT distance="150" swimtime="00:02:11.69" />
                    <SPLIT distance="175" swimtime="00:02:36.34" />
                    <SPLIT distance="200" swimtime="00:03:01.91" />
                    <SPLIT distance="225" swimtime="00:03:27.74" />
                    <SPLIT distance="250" swimtime="00:03:53.74" />
                    <SPLIT distance="275" swimtime="00:04:20.03" />
                    <SPLIT distance="300" swimtime="00:04:46.05" />
                    <SPLIT distance="325" swimtime="00:05:12.57" />
                    <SPLIT distance="350" swimtime="00:05:38.73" />
                    <SPLIT distance="375" swimtime="00:06:04.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="220" reactiontime="+110" swimtime="00:00:35.20" resultid="2236" lane="2" heatid="7339" entrytime="00:00:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.94" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="przekroczony limit 13:30:00" eventid="1075" status="DSQ" swimtime="00:14:10.34" resultid="2233" lane="6" heatid="6718" entrytime="00:13:30.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-24" firstname="Robert" gender="M" lastname="Trzos" nation="POL" athleteid="2237">
              <RESULTS>
                <RESULT eventid="1411" points="350" reactiontime="+86" swimtime="00:03:00.82" resultid="2240" lane="5" heatid="7009" entrytime="00:03:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.24" />
                    <SPLIT distance="50" swimtime="00:00:41.68" />
                    <SPLIT distance="75" swimtime="00:01:04.26" />
                    <SPLIT distance="100" swimtime="00:01:27.38" />
                    <SPLIT distance="125" swimtime="00:01:50.47" />
                    <SPLIT distance="150" swimtime="00:02:13.75" />
                    <SPLIT distance="175" swimtime="00:02:37.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="347" reactiontime="+82" swimtime="00:01:23.81" resultid="2241" lane="2" heatid="7308" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.24" />
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                    <SPLIT distance="75" swimtime="00:01:00.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="286" reactiontime="+80" swimtime="00:01:17.58" resultid="2238" lane="3" heatid="6735" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.91" />
                    <SPLIT distance="50" swimtime="00:00:36.68" />
                    <SPLIT distance="75" swimtime="00:00:58.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="351" reactiontime="+80" swimtime="00:00:38.50" resultid="2239" lane="8" heatid="6863" entrytime="00:00:37.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" name="Masters Korona Kraków 1" number="1">
              <RESULTS>
                <RESULT eventid="1341" points="304" reactiontime="+79" swimtime="00:02:22.00" resultid="2255" lane="4" heatid="6986" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.74" />
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                    <SPLIT distance="75" swimtime="00:00:53.16" />
                    <SPLIT distance="100" swimtime="00:01:14.01" />
                    <SPLIT distance="125" swimtime="00:01:30.20" />
                    <SPLIT distance="150" swimtime="00:01:49.01" />
                    <SPLIT distance="175" swimtime="00:02:05.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2192" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="2237" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="2186" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="2184" number="4" reactiontime="+96" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" name="Masters Korona Kraków C" number="1">
              <RESULTS>
                <RESULT eventid="1177" points="457" reactiontime="+79" swimtime="00:01:52.62" resultid="2246" lane="4" heatid="6809" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.81" />
                    <SPLIT distance="50" swimtime="00:00:26.76" />
                    <SPLIT distance="75" swimtime="00:00:40.62" />
                    <SPLIT distance="100" swimtime="00:00:56.01" />
                    <SPLIT distance="125" swimtime="00:01:09.42" />
                    <SPLIT distance="150" swimtime="00:01:24.59" />
                    <SPLIT distance="175" swimtime="00:01:37.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2180" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="2200" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="2171" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="2221" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" name="Masters Korona Kraków 2" number="2">
              <RESULTS>
                <RESULT eventid="1341" points="437" swimtime="00:02:05.77" resultid="2256" lane="1" heatid="6988" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.28" />
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                    <SPLIT distance="75" swimtime="00:00:47.61" />
                    <SPLIT distance="100" swimtime="00:01:07.30" />
                    <SPLIT distance="125" swimtime="00:01:20.91" />
                    <SPLIT distance="150" swimtime="00:01:37.24" />
                    <SPLIT distance="175" swimtime="00:01:50.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2180" number="1" />
                    <RELAYPOSITION athleteid="2221" number="2" reactiontime="+28" />
                    <RELAYPOSITION athleteid="2171" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="2200" number="4" reactiontime="+51" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" name="Masters Korona Kraków C" number="2">
              <RESULTS>
                <RESULT eventid="1177" status="DNS" swimtime="00:00:00.00" resultid="2247" heatid="6809" entrytime="00:02:00.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2180" number="1" />
                    <RELAYPOSITION athleteid="2200" number="2" />
                    <RELAYPOSITION athleteid="2171" number="3" />
                    <RELAYPOSITION athleteid="2221" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" name="Masters Korona Kraków D" number="3">
              <RESULTS>
                <RESULT eventid="1177" points="128" swimtime="00:02:51.92" resultid="2248" heatid="6808" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.61" />
                    <SPLIT distance="50" swimtime="00:01:11.02" />
                    <SPLIT distance="75" swimtime="00:01:28.93" />
                    <SPLIT distance="100" swimtime="00:01:48.83" />
                    <SPLIT distance="125" swimtime="00:02:04.06" />
                    <SPLIT distance="150" swimtime="00:02:21.36" />
                    <SPLIT distance="175" swimtime="00:02:35.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2228" number="1" />
                    <RELAYPOSITION athleteid="2206" number="2" reactiontime="+97" />
                    <RELAYPOSITION athleteid="2213" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="2192" number="4" reactiontime="+75" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="F" name="Masters Korona Kraków B" number="1">
              <RESULTS>
                <RESULT eventid="1160" points="212" reactiontime="+86" swimtime="00:02:44.65" resultid="2257" lane="1" heatid="6813" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.93" />
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                    <SPLIT distance="75" swimtime="00:00:58.84" />
                    <SPLIT distance="100" swimtime="00:01:22.11" />
                    <SPLIT distance="125" swimtime="00:01:38.55" />
                    <SPLIT distance="150" swimtime="00:01:57.22" />
                    <SPLIT distance="175" swimtime="00:02:19.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2118" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="2131" number="2" reactiontime="+80" />
                    <RELAYPOSITION athleteid="2123" number="3" reactiontime="+18" />
                    <RELAYPOSITION athleteid="2137" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="F" name="Masters Korona Kraków C" number="1">
              <RESULTS>
                <RESULT eventid="1324" points="211" reactiontime="+74" swimtime="00:03:01.77" resultid="2254" lane="1" heatid="6979" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.27" />
                    <SPLIT distance="50" swimtime="00:00:52.19" />
                    <SPLIT distance="75" swimtime="00:01:11.40" />
                    <SPLIT distance="100" swimtime="00:01:34.39" />
                    <SPLIT distance="125" swimtime="00:01:52.72" />
                    <SPLIT distance="150" swimtime="00:02:16.50" />
                    <SPLIT distance="175" swimtime="00:02:39.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2137" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="2118" number="2" reactiontime="+4" />
                    <RELAYPOSITION athleteid="2123" number="3" reactiontime="+70" />
                    <RELAYPOSITION athleteid="2131" number="4" reactiontime="+66" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="F" name="Masters Korona Kraków D" number="2">
              <RESULTS>
                <RESULT eventid="1160" points="317" reactiontime="+77" swimtime="00:02:23.98" resultid="2244" lane="2" heatid="6813" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.99" />
                    <SPLIT distance="50" swimtime="00:00:31.03" />
                    <SPLIT distance="75" swimtime="00:00:46.86" />
                    <SPLIT distance="100" swimtime="00:01:04.70" />
                    <SPLIT distance="125" swimtime="00:01:25.54" />
                    <SPLIT distance="150" swimtime="00:01:50.39" />
                    <SPLIT distance="175" swimtime="00:02:06.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2105" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="2147" number="2" reactiontime="+25" />
                    <RELAYPOSITION athleteid="2113" number="3" reactiontime="+85" />
                    <RELAYPOSITION athleteid="2155" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1324" points="320" reactiontime="+60" swimtime="00:02:38.32" resultid="2245" lane="2" heatid="6979" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.25" />
                    <SPLIT distance="50" swimtime="00:00:36.91" />
                    <SPLIT distance="75" swimtime="00:00:55.92" />
                    <SPLIT distance="100" swimtime="00:01:18.02" />
                    <SPLIT distance="125" swimtime="00:01:33.85" />
                    <SPLIT distance="150" swimtime="00:01:52.32" />
                    <SPLIT distance="175" swimtime="00:02:13.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2105" number="1" reactiontime="+60" />
                    <RELAYPOSITION athleteid="2147" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="2155" number="3" reactiontime="+62" />
                    <RELAYPOSITION athleteid="2113" number="4" reactiontime="+86" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" name="Masters Korona Kraków B" number="1">
              <RESULTS>
                <RESULT eventid="1615" reactiontime="+112" swimtime="00:02:23.18" resultid="2243" lane="8" heatid="7442" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.01" />
                    <SPLIT distance="50" swimtime="00:00:44.35" />
                    <SPLIT distance="75" swimtime="00:00:59.79" />
                    <SPLIT distance="100" swimtime="00:01:16.13" />
                    <SPLIT distance="125" swimtime="00:01:34.26" />
                    <SPLIT distance="150" swimtime="00:01:53.75" />
                    <SPLIT distance="175" swimtime="00:02:07.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2131" number="1" reactiontime="+112" />
                    <RELAYPOSITION athleteid="2186" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="2118" number="3" reactiontime="+30" />
                    <RELAYPOSITION athleteid="2221" number="4" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" name="Masters Korona Kraków B" number="2">
              <RESULTS>
                <RESULT eventid="1815" reactiontime="+84" swimtime="00:02:22.61" resultid="2242" lane="4" heatid="7503" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.31" />
                    <SPLIT distance="50" swimtime="00:00:42.04" />
                    <SPLIT distance="75" swimtime="00:01:01.56" />
                    <SPLIT distance="125" swimtime="00:01:37.48" />
                    <SPLIT distance="150" swimtime="00:01:53.66" />
                    <SPLIT distance="175" swimtime="00:02:07.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2163" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="2118" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="2221" number="3" />
                    <RELAYPOSITION athleteid="2200" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" name="Masters Korona Kraków C" number="2">
              <RESULTS>
                <RESULT eventid="1815" reactiontime="+63" swimtime="00:02:13.29" resultid="2250" lane="1" heatid="7504" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.36" />
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                    <SPLIT distance="75" swimtime="00:00:48.82" />
                    <SPLIT distance="100" swimtime="00:01:09.76" />
                    <SPLIT distance="125" swimtime="00:01:23.34" />
                    <SPLIT distance="150" swimtime="00:01:39.53" />
                    <SPLIT distance="175" swimtime="00:01:55.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2180" number="1" reactiontime="+63" />
                    <RELAYPOSITION athleteid="2105" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="2171" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="2155" number="4" reactiontime="+62" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1615" reactiontime="+79" swimtime="00:02:01.26" resultid="2251" lane="7" heatid="7443" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.89" />
                    <SPLIT distance="50" swimtime="00:00:26.68" />
                    <SPLIT distance="75" swimtime="00:00:41.76" />
                    <SPLIT distance="100" swimtime="00:00:57.99" />
                    <SPLIT distance="125" swimtime="00:01:14.39" />
                    <SPLIT distance="150" swimtime="00:01:31.83" />
                    <SPLIT distance="175" swimtime="00:01:46.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2180" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="2105" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="2155" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="2171" number="4" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="X" name="Masters Korona Kraków D" number="3">
              <RESULTS>
                <RESULT eventid="1815" reactiontime="+67" swimtime="00:02:33.65" resultid="2252" lane="3" heatid="7503" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.12" />
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                    <SPLIT distance="75" swimtime="00:00:54.77" />
                    <SPLIT distance="100" swimtime="00:01:16.86" />
                    <SPLIT distance="125" swimtime="00:01:35.14" />
                    <SPLIT distance="150" swimtime="00:01:58.54" />
                    <SPLIT distance="175" swimtime="00:02:15.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2192" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="2147" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="2123" number="3" reactiontime="+70" />
                    <RELAYPOSITION athleteid="2206" number="4" reactiontime="+63" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1615" reactiontime="+96" swimtime="00:02:18.62" resultid="2253" lane="2" heatid="7442" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.57" />
                    <SPLIT distance="50" swimtime="00:00:36.78" />
                    <SPLIT distance="75" swimtime="00:00:53.03" />
                    <SPLIT distance="100" swimtime="00:01:11.01" />
                    <SPLIT distance="125" swimtime="00:01:28.72" />
                    <SPLIT distance="150" swimtime="00:01:47.85" />
                    <SPLIT distance="175" swimtime="00:02:02.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2206" number="1" reactiontime="+96" />
                    <RELAYPOSITION athleteid="2147" number="2" reactiontime="+47" />
                    <RELAYPOSITION athleteid="2123" number="3" reactiontime="+79" />
                    <RELAYPOSITION athleteid="2192" number="4" reactiontime="+71" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SMKRA" name="Straz Miejska Miasta Kraków" nation="POL" region="KR">
          <CONTACT city="Kraków" name="Jawień Krzysztof" phone="505593911" state="MAŁ" />
          <ATHLETES>
            <ATHLETE birthdate="1971-06-12" firstname="Krzysztof" gender="M" lastname="Jawień" nation="POL" athleteid="2292">
              <RESULTS>
                <RESULT eventid="1696" points="453" reactiontime="+79" swimtime="00:01:16.68" resultid="2298" lane="8" heatid="7304" entrytime="00:01:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.70" />
                    <SPLIT distance="50" swimtime="00:00:36.05" />
                    <SPLIT distance="75" swimtime="00:00:56.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="430" reactiontime="+82" swimtime="00:02:48.83" resultid="2296" lane="6" heatid="7004" entrytime="00:03:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.82" />
                    <SPLIT distance="50" swimtime="00:00:38.52" />
                    <SPLIT distance="75" swimtime="00:00:59.89" />
                    <SPLIT distance="100" swimtime="00:01:21.55" />
                    <SPLIT distance="125" swimtime="00:01:43.47" />
                    <SPLIT distance="150" swimtime="00:02:05.94" />
                    <SPLIT distance="175" swimtime="00:02:27.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="336" reactiontime="+80" swimtime="00:02:41.00" resultid="2295" lane="4" heatid="6873" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.88" />
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                    <SPLIT distance="75" swimtime="00:00:53.94" />
                    <SPLIT distance="100" swimtime="00:01:14.36" />
                    <SPLIT distance="125" swimtime="00:01:35.23" />
                    <SPLIT distance="150" swimtime="00:01:57.29" />
                    <SPLIT distance="175" swimtime="00:02:18.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="479" reactiontime="+83" swimtime="00:00:34.72" resultid="2294" lane="2" heatid="6855" entrytime="00:00:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="352" reactiontime="+86" swimtime="00:05:45.09" resultid="2299" lane="5" heatid="7363" entrytime="00:06:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.13" />
                    <SPLIT distance="50" swimtime="00:00:35.08" />
                    <SPLIT distance="75" swimtime="00:00:54.67" />
                    <SPLIT distance="100" swimtime="00:01:14.54" />
                    <SPLIT distance="125" swimtime="00:01:38.01" />
                    <SPLIT distance="150" swimtime="00:02:00.64" />
                    <SPLIT distance="175" swimtime="00:02:24.27" />
                    <SPLIT distance="200" swimtime="00:02:47.21" />
                    <SPLIT distance="225" swimtime="00:03:10.91" />
                    <SPLIT distance="250" swimtime="00:03:34.80" />
                    <SPLIT distance="275" swimtime="00:03:58.27" />
                    <SPLIT distance="300" swimtime="00:04:21.71" />
                    <SPLIT distance="325" swimtime="00:04:42.87" />
                    <SPLIT distance="350" swimtime="00:05:04.13" />
                    <SPLIT distance="375" swimtime="00:05:25.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="366" reactiontime="+81" swimtime="00:01:10.41" resultid="2297" lane="7" heatid="7021" entrytime="00:01:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.09" />
                    <SPLIT distance="50" swimtime="00:00:32.44" />
                    <SPLIT distance="75" swimtime="00:00:50.93" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="04" eventid="1075" status="DSQ" swimtime="00:00:00.00" resultid="2293" lane="6" heatid="6720" entrytime="00:12:00.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAGOR" name="Masters Gorzów" nation="POL" region="LBS">
          <CONTACT city="GORZOW WLKP." email="hohtor72@wp.pl" name="ŁOPACINSKI" state="LUBUS" street="DĘBOWA" zip="66-400" />
          <ATHLETES>
            <ATHLETE birthdate="1976-03-18" firstname="Beata" gender="F" lastname="Rojewska" nation="POL" athleteid="2301">
              <RESULTS>
                <RESULT eventid="1747" points="475" reactiontime="+86" swimtime="00:00:30.71" resultid="2304" lane="2" heatid="7334" entrytime="00:00:31.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="409" reactiontime="+82" swimtime="00:00:34.29" resultid="2303" lane="1" heatid="7280" entrytime="00:00:34.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="434" reactiontime="+68" swimtime="00:00:36.54" resultid="2302" heatid="7031" entrytime="00:00:36.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-05-08" firstname="Dawid" gender="M" lastname="Borus" nation="POL" athleteid="2305">
              <RESULTS>
                <RESULT eventid="1730" points="405" reactiontime="+66" swimtime="00:01:11.01" resultid="2308" lane="5" heatid="7324" entrytime="00:01:13.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.84" />
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                    <SPLIT distance="75" swimtime="00:00:52.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="400" reactiontime="+65" swimtime="00:00:33.20" resultid="2307" lane="3" heatid="7039" entrytime="00:00:34.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="433" reactiontime="+79" swimtime="00:00:28.11" resultid="2309" lane="8" heatid="7350" entrytime="00:00:27.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="399" reactiontime="+79" swimtime="00:01:03.89" resultid="2306" lane="2" heatid="6841" entrytime="00:01:03.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.35" />
                    <SPLIT distance="50" swimtime="00:00:30.55" />
                    <SPLIT distance="75" swimtime="00:00:46.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-06-11" firstname="Artur" gender="M" lastname="Łopaciński" nation="POL" athleteid="2310">
              <RESULTS>
                <RESULT eventid="1496" points="334" reactiontime="+58" swimtime="00:00:35.25" resultid="2311" lane="6" heatid="7039" entrytime="00:00:34.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="403" reactiontime="+51" swimtime="00:00:28.80" resultid="2314" lane="4" heatid="7346" entrytime="00:00:28.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="373" reactiontime="+62" swimtime="00:00:31.89" resultid="2313" lane="3" heatid="7287" entrytime="00:00:32.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" status="DNS" swimtime="00:00:00.00" resultid="2312" lane="1" heatid="7078" entrytime="00:02:45.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-09-21" firstname="Maciej" gender="M" lastname="Szypiórkowski" nation="POL" athleteid="2315">
              <RESULTS>
                <RESULT eventid="1696" points="306" reactiontime="+86" swimtime="00:01:27.39" resultid="2317" lane="1" heatid="7306" entrytime="00:01:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.69" />
                    <SPLIT distance="50" swimtime="00:00:41.07" />
                    <SPLIT distance="75" swimtime="00:01:03.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="163" reactiontime="+83" swimtime="00:01:32.14" resultid="2316" lane="3" heatid="7017" entrytime="00:01:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.95" />
                    <SPLIT distance="50" swimtime="00:00:42.09" />
                    <SPLIT distance="75" swimtime="00:01:07.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="281" reactiontime="+91" swimtime="00:00:32.48" resultid="2318" lane="8" heatid="7341" entrytime="00:00:32.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAOPO" name="Tp Masters Opole" nation="POL">
          <CONTACT city="OPOLE" email="krasnodebski@cb.com.pl" name="KRASNODĘBSKI" phone="694402057" />
          <ATHLETES>
            <ATHLETE birthdate="1931-01-01" firstname="Józef" gender="M" lastname="Kasperek" nation="POL" athleteid="2320">
              <RESULTS>
                <RESULT eventid="1564" points="20" reactiontime="+102" swimtime="00:06:16.58" resultid="2324" lane="6" heatid="7054" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:35.65" />
                    <SPLIT distance="50" swimtime="00:01:20.10" />
                    <SPLIT distance="75" swimtime="00:02:07.56" />
                    <SPLIT distance="100" swimtime="00:02:57.25" />
                    <SPLIT distance="125" swimtime="00:03:49.27" />
                    <SPLIT distance="150" swimtime="00:04:41.55" />
                    <SPLIT distance="175" swimtime="00:05:31.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="25" reactiontime="+80" swimtime="00:02:59.39" resultid="2325" lane="5" heatid="7318" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:41.08" />
                    <SPLIT distance="50" swimtime="00:01:26.18" />
                    <SPLIT distance="75" swimtime="00:02:12.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="22" reactiontime="+80" swimtime="00:01:26.12" resultid="2323" lane="3" heatid="7032" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:40.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="31" reactiontime="+112" swimtime="00:01:07.53" resultid="2326" lane="1" heatid="7336" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.00" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1205" points="24" reactiontime="+114" swimtime="00:02:41.89" resultid="2322" lane="7" heatid="6830" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.27" />
                    <SPLIT distance="50" swimtime="00:01:12.92" />
                    <SPLIT distance="75" swimtime="00:01:55.67" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="przekroczony limit 27:00:00" eventid="1075" status="DSQ" swimtime="00:27:45.91" resultid="2321" lane="5" heatid="6716" entrytime="00:25:23.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-01" firstname="Grzegorz" gender="M" lastname="Radomski" nation="POL" athleteid="2327">
              <RESULTS>
                <RESULT eventid="1730" points="612" reactiontime="+69" swimtime="00:01:01.86" resultid="2333" lane="5" heatid="7326" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.57" />
                    <SPLIT distance="50" swimtime="00:00:29.75" />
                    <SPLIT distance="75" swimtime="00:00:45.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="579" reactiontime="+77" swimtime="00:04:52.45" resultid="2334" lane="5" heatid="7364" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.03" />
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                    <SPLIT distance="75" swimtime="00:00:48.31" />
                    <SPLIT distance="100" swimtime="00:01:06.98" />
                    <SPLIT distance="125" swimtime="00:01:25.23" />
                    <SPLIT distance="150" swimtime="00:01:42.97" />
                    <SPLIT distance="175" swimtime="00:02:01.52" />
                    <SPLIT distance="200" swimtime="00:02:20.22" />
                    <SPLIT distance="225" swimtime="00:02:40.49" />
                    <SPLIT distance="250" swimtime="00:03:01.34" />
                    <SPLIT distance="275" swimtime="00:03:22.33" />
                    <SPLIT distance="300" swimtime="00:03:43.81" />
                    <SPLIT distance="325" swimtime="00:04:01.76" />
                    <SPLIT distance="350" swimtime="00:04:18.81" />
                    <SPLIT distance="375" swimtime="00:04:36.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="594" reactiontime="+75" swimtime="00:02:15.86" resultid="2332" lane="5" heatid="7080" entrytime="00:02:21.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.53" />
                    <SPLIT distance="50" swimtime="00:00:29.15" />
                    <SPLIT distance="75" swimtime="00:00:45.89" />
                    <SPLIT distance="100" swimtime="00:01:02.49" />
                    <SPLIT distance="125" swimtime="00:01:21.66" />
                    <SPLIT distance="150" swimtime="00:01:41.81" />
                    <SPLIT distance="175" swimtime="00:01:59.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="615" reactiontime="+72" swimtime="00:02:13.95" resultid="2329" lane="4" heatid="6887" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.83" />
                    <SPLIT distance="50" swimtime="00:00:30.40" />
                    <SPLIT distance="75" swimtime="00:00:46.78" />
                    <SPLIT distance="100" swimtime="00:01:03.67" />
                    <SPLIT distance="125" swimtime="00:01:20.83" />
                    <SPLIT distance="150" swimtime="00:01:38.39" />
                    <SPLIT distance="175" swimtime="00:01:56.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="507" swimtime="00:18:16.59" resultid="2328" lane="4" heatid="6752" entrytime="00:18:05.00" />
                <RESULT eventid="1375" points="557" reactiontime="+78" swimtime="00:04:27.38" resultid="2330" lane="5" heatid="6909" entrytime="00:04:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.37" />
                    <SPLIT distance="50" swimtime="00:00:28.77" />
                    <SPLIT distance="75" swimtime="00:00:44.72" />
                    <SPLIT distance="100" swimtime="00:01:01.05" />
                    <SPLIT distance="125" swimtime="00:01:17.45" />
                    <SPLIT distance="150" swimtime="00:01:34.14" />
                    <SPLIT distance="175" swimtime="00:01:50.88" />
                    <SPLIT distance="200" swimtime="00:02:08.01" />
                    <SPLIT distance="225" swimtime="00:02:25.05" />
                    <SPLIT distance="250" swimtime="00:02:42.51" />
                    <SPLIT distance="275" swimtime="00:02:59.67" />
                    <SPLIT distance="300" swimtime="00:03:17.27" />
                    <SPLIT distance="325" swimtime="00:03:34.68" />
                    <SPLIT distance="350" swimtime="00:03:52.39" />
                    <SPLIT distance="375" swimtime="00:04:10.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="406" reactiontime="+78" swimtime="00:02:19.03" resultid="2331" lane="3" heatid="7065" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.45" />
                    <SPLIT distance="50" swimtime="00:00:30.98" />
                    <SPLIT distance="75" swimtime="00:00:48.28" />
                    <SPLIT distance="100" swimtime="00:01:06.02" />
                    <SPLIT distance="125" swimtime="00:01:23.99" />
                    <SPLIT distance="150" swimtime="00:01:42.16" />
                    <SPLIT distance="175" swimtime="00:02:00.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Jerzy" gender="M" lastname="Minkiewicz" nation="POL" athleteid="2335">
              <RESULTS>
                <RESULT eventid="1462" points="198" reactiontime="+91" swimtime="00:01:26.36" resultid="2339" lane="3" heatid="7018" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.95" />
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                    <SPLIT distance="75" swimtime="00:01:01.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="141" reactiontime="+105" swimtime="00:03:35.04" resultid="2338" lane="4" heatid="6871" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.99" />
                    <SPLIT distance="50" swimtime="00:00:42.88" />
                    <SPLIT distance="75" swimtime="00:01:08.69" />
                    <SPLIT distance="100" swimtime="00:01:36.46" />
                    <SPLIT distance="125" swimtime="00:02:05.02" />
                    <SPLIT distance="150" swimtime="00:02:35.36" />
                    <SPLIT distance="175" swimtime="00:03:05.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="234" reactiontime="+91" swimtime="00:01:22.93" resultid="2336" lane="5" heatid="6735" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.33" />
                    <SPLIT distance="50" swimtime="00:00:38.83" />
                    <SPLIT distance="75" swimtime="00:01:04.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="309" reactiontime="+83" swimtime="00:01:09.52" resultid="2337" lane="5" heatid="6837" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.68" />
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                    <SPLIT distance="75" swimtime="00:00:51.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="268" reactiontime="+83" swimtime="00:00:35.58" resultid="2340" lane="4" heatid="7285" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="319" reactiontime="+88" swimtime="00:00:31.12" resultid="2341" lane="7" heatid="7343" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-01-01" firstname="Katarzyna" gender="F" lastname="Stolarczyk" nation="POL" athleteid="2342">
              <RESULTS>
                <RESULT eventid="1290" points="371" reactiontime="+75" swimtime="00:02:54.20" resultid="2344" heatid="6879" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.83" />
                    <SPLIT distance="50" swimtime="00:00:41.23" />
                    <SPLIT distance="75" swimtime="00:01:02.20" />
                    <SPLIT distance="100" swimtime="00:01:24.13" />
                    <SPLIT distance="125" swimtime="00:01:46.41" />
                    <SPLIT distance="150" swimtime="00:02:09.10" />
                    <SPLIT distance="175" swimtime="00:02:32.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="406" reactiontime="+73" swimtime="00:01:19.34" resultid="2346" heatid="7317" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.56" />
                    <SPLIT distance="50" swimtime="00:00:38.17" />
                    <SPLIT distance="75" swimtime="00:00:58.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="412" reactiontime="+75" swimtime="00:00:37.17" resultid="2345" lane="5" heatid="7030" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="345" reactiontime="+79" swimtime="00:01:23.81" resultid="2343" lane="8" heatid="6729" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.43" />
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                    <SPLIT distance="75" swimtime="00:01:03.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-01-01" firstname="Józef" gender="M" lastname="Ciupek" nation="POL" athleteid="2347">
              <RESULTS>
                <RESULT eventid="1645" points="198" reactiontime="+97" swimtime="00:00:39.39" resultid="2349" lane="2" heatid="7283" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="274" reactiontime="+93" swimtime="00:00:41.80" resultid="2348" lane="7" heatid="6858" entrytime="00:00:41.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Roman" gender="M" lastname="Birecki" nation="POL" athleteid="2350">
              <RESULTS>
                <RESULT eventid="1462" points="231" reactiontime="+102" swimtime="00:01:22.05" resultid="2354" lane="7" heatid="7019" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.90" />
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                    <SPLIT distance="75" swimtime="00:00:59.70" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1273" points="225" reactiontime="+102" swimtime="00:03:04.10" resultid="2352" lane="4" heatid="6872" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.06" />
                    <SPLIT distance="50" swimtime="00:00:40.06" />
                    <SPLIT distance="75" swimtime="00:01:02.96" />
                    <SPLIT distance="100" swimtime="00:01:26.81" />
                    <SPLIT distance="125" swimtime="00:01:51.05" />
                    <SPLIT distance="150" swimtime="00:02:15.40" />
                    <SPLIT distance="175" swimtime="00:02:39.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="244" swimtime="00:12:13.69" resultid="2351" lane="7" heatid="6719" entrytime="00:12:27.00" />
                <RESULT eventid="1564" points="274" reactiontime="+103" swimtime="00:02:38.39" resultid="2355" lane="2" heatid="7059" entrytime="00:02:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.80" />
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                    <SPLIT distance="75" swimtime="00:00:55.56" />
                    <SPLIT distance="100" swimtime="00:01:16.16" />
                    <SPLIT distance="125" swimtime="00:01:36.97" />
                    <SPLIT distance="150" swimtime="00:01:58.29" />
                    <SPLIT distance="175" swimtime="00:02:18.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="276" reactiontime="+97" swimtime="00:00:35.26" resultid="2356" lane="5" heatid="7286" entrytime="00:00:34.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="241" reactiontime="+111" swimtime="00:05:53.58" resultid="2353" lane="6" heatid="6904" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.07" />
                    <SPLIT distance="50" swimtime="00:00:38.42" />
                    <SPLIT distance="75" swimtime="00:00:59.21" />
                    <SPLIT distance="100" swimtime="00:01:20.88" />
                    <SPLIT distance="125" swimtime="00:01:43.45" />
                    <SPLIT distance="150" swimtime="00:02:06.08" />
                    <SPLIT distance="175" swimtime="00:02:28.65" />
                    <SPLIT distance="200" swimtime="00:02:51.38" />
                    <SPLIT distance="225" swimtime="00:03:13.55" />
                    <SPLIT distance="250" swimtime="00:03:36.53" />
                    <SPLIT distance="275" swimtime="00:03:59.45" />
                    <SPLIT distance="300" swimtime="00:04:22.94" />
                    <SPLIT distance="325" swimtime="00:04:45.51" />
                    <SPLIT distance="350" swimtime="00:05:08.68" />
                    <SPLIT distance="375" swimtime="00:05:31.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="311" reactiontime="+99" swimtime="00:00:31.38" resultid="2357" lane="3" heatid="7342" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Olgierd" gender="M" lastname="Mikosza" nation="POL" athleteid="2358">
              <RESULTS>
                <RESULT eventid="1307" points="209" reactiontime="+83" swimtime="00:03:11.78" resultid="2360" heatid="6884" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.55" />
                    <SPLIT distance="50" swimtime="00:00:42.84" />
                    <SPLIT distance="75" swimtime="00:01:06.01" />
                    <SPLIT distance="100" swimtime="00:01:30.70" />
                    <SPLIT distance="125" swimtime="00:01:56.56" />
                    <SPLIT distance="150" swimtime="00:02:22.20" />
                    <SPLIT distance="175" swimtime="00:02:47.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="173" reactiontime="+87" swimtime="00:01:30.28" resultid="2362" lane="7" heatid="7017" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.08" />
                    <SPLIT distance="50" swimtime="00:00:41.64" />
                    <SPLIT distance="75" swimtime="00:01:06.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="190" reactiontime="+98" swimtime="00:07:03.83" resultid="2365" lane="3" heatid="7360" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.25" />
                    <SPLIT distance="50" swimtime="00:00:45.58" />
                    <SPLIT distance="75" swimtime="00:01:12.58" />
                    <SPLIT distance="100" swimtime="00:01:40.18" />
                    <SPLIT distance="125" swimtime="00:02:08.81" />
                    <SPLIT distance="150" swimtime="00:02:36.19" />
                    <SPLIT distance="175" swimtime="00:03:03.53" />
                    <SPLIT distance="200" swimtime="00:03:29.59" />
                    <SPLIT distance="225" swimtime="00:04:00.46" />
                    <SPLIT distance="250" swimtime="00:04:30.75" />
                    <SPLIT distance="275" swimtime="00:05:00.53" />
                    <SPLIT distance="300" swimtime="00:05:31.41" />
                    <SPLIT distance="325" swimtime="00:05:56.44" />
                    <SPLIT distance="350" swimtime="00:06:19.66" />
                    <SPLIT distance="375" swimtime="00:06:42.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="226" swimtime="00:12:32.84" resultid="2359" lane="2" heatid="6718" entrytime="00:13:19.00" />
                <RESULT eventid="1375" points="216" reactiontime="+92" swimtime="00:06:06.64" resultid="2361" lane="7" heatid="6903" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.40" />
                    <SPLIT distance="50" swimtime="00:00:37.88" />
                    <SPLIT distance="75" swimtime="00:01:00.48" />
                    <SPLIT distance="100" swimtime="00:01:23.00" />
                    <SPLIT distance="125" swimtime="00:01:46.84" />
                    <SPLIT distance="150" swimtime="00:02:11.57" />
                    <SPLIT distance="175" swimtime="00:02:34.64" />
                    <SPLIT distance="200" swimtime="00:02:58.65" />
                    <SPLIT distance="225" swimtime="00:03:22.76" />
                    <SPLIT distance="250" swimtime="00:03:46.71" />
                    <SPLIT distance="275" swimtime="00:04:11.24" />
                    <SPLIT distance="300" swimtime="00:04:35.18" />
                    <SPLIT distance="325" swimtime="00:04:58.85" />
                    <SPLIT distance="350" swimtime="00:05:22.59" />
                    <SPLIT distance="375" swimtime="00:05:45.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="226" reactiontime="+89" swimtime="00:02:49.03" resultid="2363" lane="2" heatid="7058" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.37" />
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                    <SPLIT distance="75" swimtime="00:00:57.30" />
                    <SPLIT distance="100" swimtime="00:01:19.58" />
                    <SPLIT distance="125" swimtime="00:01:42.13" />
                    <SPLIT distance="150" swimtime="00:02:05.26" />
                    <SPLIT distance="175" swimtime="00:02:28.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="234" reactiontime="+76" swimtime="00:01:25.21" resultid="2364" lane="2" heatid="7322" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.25" />
                    <SPLIT distance="50" swimtime="00:00:40.64" />
                    <SPLIT distance="75" swimtime="00:01:03.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1937-01-01" firstname="Tadeusz" gender="M" lastname="Witkowski" nation="POL" athleteid="2366">
              <RESULTS>
                <RESULT eventid="1307" points="117" reactiontime="+89" swimtime="00:03:52.47" resultid="2369" lane="4" heatid="6881" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.61" />
                    <SPLIT distance="50" swimtime="00:00:54.58" />
                    <SPLIT distance="75" swimtime="00:01:23.43" />
                    <SPLIT distance="100" swimtime="00:01:53.49" />
                    <SPLIT distance="125" swimtime="00:02:23.68" />
                    <SPLIT distance="150" swimtime="00:02:54.28" />
                    <SPLIT distance="175" swimtime="00:03:24.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="162" reactiontime="+106" swimtime="00:01:26.23" resultid="2368" heatid="6832" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.12" />
                    <SPLIT distance="50" swimtime="00:00:39.24" />
                    <SPLIT distance="75" swimtime="00:01:02.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="120" reactiontime="+87" swimtime="00:00:49.60" resultid="2370" lane="7" heatid="7034" entrytime="00:00:50.00" />
                <RESULT eventid="1730" points="116" reactiontime="+85" swimtime="00:01:47.62" resultid="2372" lane="3" heatid="7319" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.91" />
                    <SPLIT distance="50" swimtime="00:00:52.68" />
                    <SPLIT distance="75" swimtime="00:01:21.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="227" reactiontime="+105" swimtime="00:00:34.88" resultid="2373" lane="5" heatid="7339" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="119" reactiontime="+101" swimtime="00:03:29.29" resultid="2371" lane="7" heatid="7055" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.41" />
                    <SPLIT distance="50" swimtime="00:00:46.13" />
                    <SPLIT distance="75" swimtime="00:01:13.95" />
                    <SPLIT distance="100" swimtime="00:01:40.92" />
                    <SPLIT distance="125" swimtime="00:02:08.13" />
                    <SPLIT distance="150" swimtime="00:02:35.18" />
                    <SPLIT distance="175" swimtime="00:03:04.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="107" reactiontime="+111" swimtime="00:01:47.44" resultid="2367" lane="7" heatid="6731" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.66" />
                    <SPLIT distance="50" swimtime="00:00:51.84" />
                    <SPLIT distance="75" swimtime="00:01:25.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="Janusz" gender="M" lastname="Szpala" nation="POL" athleteid="2374">
              <RESULTS>
                <RESULT eventid="1109" points="122" reactiontime="+100" swimtime="00:01:43.12" resultid="2375" lane="6" heatid="6731" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.90" />
                    <SPLIT distance="50" swimtime="00:00:48.76" />
                    <SPLIT distance="75" swimtime="00:01:19.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="186" reactiontime="+104" swimtime="00:00:37.22" resultid="2379" lane="7" heatid="7338" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="121" reactiontime="+97" swimtime="00:00:46.30" resultid="2378" heatid="7283" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1530" points="176" reactiontime="+102" swimtime="00:00:37.91" resultid="2376" lane="5" heatid="7047" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" status="DNS" swimtime="00:00:00.00" resultid="2377" lane="4" heatid="7072" entrytime="00:03:56.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1177" points="247" reactiontime="+78" swimtime="00:02:18.26" resultid="2380" lane="2" heatid="6808" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.62" />
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                    <SPLIT distance="75" swimtime="00:00:48.12" />
                    <SPLIT distance="100" swimtime="00:01:10.04" />
                    <SPLIT distance="125" swimtime="00:01:25.14" />
                    <SPLIT distance="150" swimtime="00:01:41.70" />
                    <SPLIT distance="175" swimtime="00:01:58.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2358" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="2366" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="2335" number="3" reactiontime="+78" />
                    <RELAYPOSITION athleteid="2347" number="4" reactiontime="+71" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1341" points="234" reactiontime="+76" swimtime="00:02:34.84" resultid="2381" lane="2" heatid="6986" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.47" />
                    <SPLIT distance="50" swimtime="00:00:41.27" />
                    <SPLIT distance="75" swimtime="00:00:59.84" />
                    <SPLIT distance="100" swimtime="00:01:22.75" />
                    <SPLIT distance="125" swimtime="00:01:39.45" />
                    <SPLIT distance="150" swimtime="00:01:58.72" />
                    <SPLIT distance="175" swimtime="00:02:16.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2358" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="2347" number="2" reactiontime="+40" />
                    <RELAYPOSITION athleteid="2350" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="2366" number="4" reactiontime="+76" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MAPOL" name="KS Masters Polkowice" nation="POL" region="DOL">
          <CONTACT city="Polkowice" email="bogdan.jawor@gmail.com" name="Jawor Bogdan" phone="519102742" state="DOL" street="Kollejowa 6/5" zip="59-100" />
          <ATHLETES>
            <ATHLETE birthdate="1952-05-30" firstname="Grażyna" gender="F" lastname="Grzegorzewska" nation="POL" athleteid="2390">
              <RESULTS>
                <RESULT eventid="1058" points="152" swimtime="00:15:25.29" resultid="2391" lane="1" heatid="6714" entrytime="00:14:49.00" entrycourse="SCM" />
                <RESULT eventid="1547" points="153" reactiontime="+96" swimtime="00:03:34.45" resultid="2395" heatid="7050" entrytime="00:03:33.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.92" />
                    <SPLIT distance="50" swimtime="00:00:48.40" />
                    <SPLIT distance="75" swimtime="00:01:16.01" />
                    <SPLIT distance="100" swimtime="00:01:44.15" />
                    <SPLIT distance="125" swimtime="00:02:13.33" />
                    <SPLIT distance="150" swimtime="00:02:42.10" />
                    <SPLIT distance="175" swimtime="00:03:09.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="172" reactiontime="+95" swimtime="00:01:34.99" resultid="2392" lane="7" heatid="6824" entrytime="00:01:34.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.65" />
                    <SPLIT distance="50" swimtime="00:00:45.38" />
                    <SPLIT distance="75" swimtime="00:01:10.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="103" reactiontime="+95" swimtime="00:00:54.23" resultid="2396" lane="7" heatid="7276" entrytime="00:00:52.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="199" reactiontime="+92" swimtime="00:00:41.01" resultid="2397" lane="6" heatid="7330" entrytime="00:00:40.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="130" reactiontime="+65" swimtime="00:00:54.51" resultid="2394" lane="5" heatid="7026" entrytime="00:00:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="145" reactiontime="+99" swimtime="00:07:39.74" resultid="2393" lane="5" heatid="6894" entrytime="00:07:53.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.51" />
                    <SPLIT distance="50" swimtime="00:00:48.53" />
                    <SPLIT distance="75" swimtime="00:01:16.71" />
                    <SPLIT distance="100" swimtime="00:01:45.80" />
                    <SPLIT distance="125" swimtime="00:02:16.27" />
                    <SPLIT distance="150" swimtime="00:02:46.62" />
                    <SPLIT distance="175" swimtime="00:03:16.89" />
                    <SPLIT distance="200" swimtime="00:03:46.48" />
                    <SPLIT distance="225" swimtime="00:04:16.20" />
                    <SPLIT distance="250" swimtime="00:04:46.41" />
                    <SPLIT distance="275" swimtime="00:05:16.67" />
                    <SPLIT distance="300" swimtime="00:05:46.36" />
                    <SPLIT distance="325" swimtime="00:06:16.33" />
                    <SPLIT distance="350" swimtime="00:06:45.92" />
                    <SPLIT distance="375" swimtime="00:07:14.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-06-21" firstname="Bogdan" gender="M" lastname="Puchalski" nation="POL" athleteid="2398">
              <RESULTS>
                <RESULT eventid="1143" points="180" swimtime="00:25:46.95" resultid="2399" lane="4" heatid="6749" entrytime="00:25:00.00" entrycourse="SCM" />
                <RESULT eventid="1411" points="223" reactiontime="+88" swimtime="00:03:30.14" resultid="2402" lane="7" heatid="7006" entrytime="00:03:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.87" />
                    <SPLIT distance="50" swimtime="00:00:47.29" />
                    <SPLIT distance="75" swimtime="00:01:13.14" />
                    <SPLIT distance="100" swimtime="00:01:40.73" />
                    <SPLIT distance="125" swimtime="00:02:08.54" />
                    <SPLIT distance="150" swimtime="00:02:36.05" />
                    <SPLIT distance="175" swimtime="00:03:03.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="158" reactiontime="+88" swimtime="00:07:30.11" resultid="2405" lane="5" heatid="7359" entrytime="00:07:31.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.52" />
                    <SPLIT distance="50" swimtime="00:00:49.60" />
                    <SPLIT distance="75" swimtime="00:01:17.75" />
                    <SPLIT distance="100" swimtime="00:01:46.39" />
                    <SPLIT distance="125" swimtime="00:02:20.55" />
                    <SPLIT distance="150" swimtime="00:02:52.25" />
                    <SPLIT distance="175" swimtime="00:03:24.65" />
                    <SPLIT distance="200" swimtime="00:03:56.48" />
                    <SPLIT distance="225" swimtime="00:04:24.65" />
                    <SPLIT distance="250" swimtime="00:04:52.46" />
                    <SPLIT distance="275" swimtime="00:05:20.73" />
                    <SPLIT distance="300" swimtime="00:05:49.78" />
                    <SPLIT distance="325" swimtime="00:06:15.39" />
                    <SPLIT distance="350" swimtime="00:06:41.01" />
                    <SPLIT distance="375" swimtime="00:07:06.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="223" reactiontime="+85" swimtime="00:01:37.03" resultid="2404" lane="6" heatid="7306" entrytime="00:01:33.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.50" />
                    <SPLIT distance="50" swimtime="00:00:45.90" />
                    <SPLIT distance="75" swimtime="00:01:10.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="244" reactiontime="+90" swimtime="00:00:43.49" resultid="2401" lane="4" heatid="6857" entrytime="00:00:42.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="120" reactiontime="+89" swimtime="00:01:42.05" resultid="2403" lane="5" heatid="7016" entrytime="00:01:41.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.07" />
                    <SPLIT distance="50" swimtime="00:00:45.75" />
                    <SPLIT distance="75" swimtime="00:01:12.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="256" reactiontime="+91" swimtime="00:01:14.05" resultid="2400" lane="6" heatid="6835" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.89" />
                    <SPLIT distance="50" swimtime="00:00:35.52" />
                    <SPLIT distance="75" swimtime="00:00:54.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-04-23" firstname="Bogdan" gender="M" lastname="Jawor" nation="POL" athleteid="2406">
              <RESULTS>
                <RESULT eventid="1143" points="105" swimtime="00:30:50.00" resultid="2407" heatid="6749" entrytime="00:30:00.00" entrycourse="SCM" />
                <RESULT eventid="1598" points="74" reactiontime="+87" swimtime="00:04:31.55" resultid="2411" lane="7" heatid="7072" entrytime="00:04:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.43" />
                    <SPLIT distance="50" swimtime="00:00:56.62" />
                    <SPLIT distance="75" swimtime="00:01:34.71" />
                    <SPLIT distance="100" swimtime="00:02:09.96" />
                    <SPLIT distance="125" swimtime="00:02:47.38" />
                    <SPLIT distance="150" swimtime="00:03:24.89" />
                    <SPLIT distance="175" swimtime="00:04:02.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="60" reactiontime="+83" swimtime="00:04:49.62" resultid="2409" lane="8" heatid="6881" entrytime="00:05:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:31.78" />
                    <SPLIT distance="50" swimtime="00:01:08.71" />
                    <SPLIT distance="75" swimtime="00:01:46.89" />
                    <SPLIT distance="100" swimtime="00:02:24.30" />
                    <SPLIT distance="125" swimtime="00:03:02.13" />
                    <SPLIT distance="150" swimtime="00:03:39.00" />
                    <SPLIT distance="175" swimtime="00:04:15.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="127" reactiontime="+95" swimtime="00:01:56.93" resultid="2413" lane="7" heatid="7303" entrytime="00:01:58.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.18" />
                    <SPLIT distance="50" swimtime="00:00:55.85" />
                    <SPLIT distance="75" swimtime="00:01:27.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="103" reactiontime="+93" swimtime="00:04:31.16" resultid="2410" lane="8" heatid="7003" entrytime="00:04:26.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.77" />
                    <SPLIT distance="50" swimtime="00:01:00.67" />
                    <SPLIT distance="75" swimtime="00:01:34.21" />
                    <SPLIT distance="100" swimtime="00:02:08.96" />
                    <SPLIT distance="125" swimtime="00:02:44.29" />
                    <SPLIT distance="150" swimtime="00:03:20.76" />
                    <SPLIT distance="175" swimtime="00:03:57.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="74" reactiontime="+101" swimtime="00:00:54.65" resultid="2412" lane="2" heatid="7281" entrytime="00:00:51.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.09" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K 11" eventid="1239" reactiontime="+93" status="DSQ" swimtime="00:00:51.23" resultid="2408" lane="7" heatid="6855" entrytime="00:00:51.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DECIE" name="MTP Delfin Cieszyn" nation="POL" region="SLA">
          <CONTACT name="Widzik" />
          <ATHLETES>
            <ATHLETE birthdate="1990-06-12" firstname="Katarzyna" gender="F" lastname="Widzik" nation="POL" athleteid="2415">
              <RESULTS>
                <RESULT eventid="1781" points="387" reactiontime="+94" swimtime="00:06:09.47" resultid="2422" lane="5" heatid="7356" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.97" />
                    <SPLIT distance="50" swimtime="00:00:40.49" />
                    <SPLIT distance="75" swimtime="00:01:04.10" />
                    <SPLIT distance="100" swimtime="00:01:28.78" />
                    <SPLIT distance="125" swimtime="00:01:51.88" />
                    <SPLIT distance="150" swimtime="00:02:14.39" />
                    <SPLIT distance="175" swimtime="00:02:36.91" />
                    <SPLIT distance="200" swimtime="00:02:58.93" />
                    <SPLIT distance="225" swimtime="00:03:25.07" />
                    <SPLIT distance="250" swimtime="00:03:51.84" />
                    <SPLIT distance="275" swimtime="00:04:19.26" />
                    <SPLIT distance="300" swimtime="00:04:45.92" />
                    <SPLIT distance="325" swimtime="00:05:07.57" />
                    <SPLIT distance="350" swimtime="00:05:28.32" />
                    <SPLIT distance="375" swimtime="00:05:49.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1126" points="357" swimtime="00:22:07.75" resultid="2416" lane="4" heatid="6747" entrytime="00:19:40.00" />
                <RESULT eventid="1290" points="456" reactiontime="+70" swimtime="00:02:42.68" resultid="2417" lane="4" heatid="6879" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.71" />
                    <SPLIT distance="50" swimtime="00:00:37.11" />
                    <SPLIT distance="75" swimtime="00:00:57.31" />
                    <SPLIT distance="100" swimtime="00:01:18.09" />
                    <SPLIT distance="125" swimtime="00:01:39.15" />
                    <SPLIT distance="150" swimtime="00:02:00.30" />
                    <SPLIT distance="175" swimtime="00:02:21.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="405" reactiontime="+93" swimtime="00:05:26.33" resultid="2418" heatid="6897" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.98" />
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                    <SPLIT distance="75" swimtime="00:00:56.70" />
                    <SPLIT distance="100" swimtime="00:01:17.03" />
                    <SPLIT distance="125" swimtime="00:01:37.67" />
                    <SPLIT distance="150" swimtime="00:01:58.57" />
                    <SPLIT distance="175" swimtime="00:02:19.58" />
                    <SPLIT distance="200" swimtime="00:02:40.53" />
                    <SPLIT distance="225" swimtime="00:03:01.14" />
                    <SPLIT distance="250" swimtime="00:03:22.38" />
                    <SPLIT distance="275" swimtime="00:03:43.29" />
                    <SPLIT distance="300" swimtime="00:04:04.44" />
                    <SPLIT distance="325" swimtime="00:04:25.30" />
                    <SPLIT distance="350" swimtime="00:04:46.28" />
                    <SPLIT distance="375" swimtime="00:05:06.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="478" reactiontime="+64" swimtime="00:00:35.37" resultid="2419" lane="2" heatid="7031" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="471" reactiontime="+60" swimtime="00:01:15.50" resultid="2421" lane="4" heatid="7317" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.44" />
                    <SPLIT distance="50" swimtime="00:00:36.33" />
                    <SPLIT distance="75" swimtime="00:00:56.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="406" reactiontime="+89" swimtime="00:02:35.04" resultid="2420" lane="6" heatid="7053" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.40" />
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                    <SPLIT distance="75" swimtime="00:00:54.27" />
                    <SPLIT distance="100" swimtime="00:01:14.02" />
                    <SPLIT distance="125" swimtime="00:01:34.33" />
                    <SPLIT distance="150" swimtime="00:01:54.82" />
                    <SPLIT distance="175" swimtime="00:02:15.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Łukasz" gender="M" lastname="Widzik" nation="POL" athleteid="2423">
              <RESULTS>
                <RESULT eventid="1075" points="420" swimtime="00:10:12.18" resultid="2424" lane="2" heatid="6722" entrytime="00:09:58.00" />
                <RESULT eventid="1307" points="456" reactiontime="+59" swimtime="00:02:28.01" resultid="2425" lane="1" heatid="6887" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.19" />
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                    <SPLIT distance="75" swimtime="00:00:52.17" />
                    <SPLIT distance="100" swimtime="00:01:10.82" />
                    <SPLIT distance="125" swimtime="00:01:29.59" />
                    <SPLIT distance="150" swimtime="00:01:49.09" />
                    <SPLIT distance="175" swimtime="00:02:08.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="451" reactiontime="+61" swimtime="00:01:08.47" resultid="2427" lane="8" heatid="7326" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.91" />
                    <SPLIT distance="50" swimtime="00:00:33.14" />
                    <SPLIT distance="75" swimtime="00:00:50.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="449" reactiontime="+65" swimtime="00:00:31.94" resultid="2426" lane="8" heatid="7043" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-09-07" firstname="Ryszard" gender="M" lastname="Jabłecki" nation="POL" athleteid="2428">
              <RESULTS>
                <RESULT eventid="1696" points="156" reactiontime="+126" swimtime="00:01:49.20" resultid="2431" lane="1" heatid="7304" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.42" />
                    <SPLIT distance="50" swimtime="00:00:49.46" />
                    <SPLIT distance="75" swimtime="00:01:18.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="128" reactiontime="+115" swimtime="00:00:42.15" resultid="2432" lane="8" heatid="7338" entrytime="00:00:37.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.29" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K  14" eventid="1411" reactiontime="+117" status="DSQ" swimtime="00:00:00.00" resultid="2430" lane="6" heatid="7003" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.59" />
                    <SPLIT distance="50" swimtime="00:00:52.63" />
                    <SPLIT distance="75" swimtime="00:01:23.39" />
                    <SPLIT distance="100" swimtime="00:01:55.01" />
                    <SPLIT distance="125" swimtime="00:02:26.83" />
                    <SPLIT distance="150" swimtime="00:02:58.43" />
                    <SPLIT distance="175" swimtime="00:03:28.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="2429" lane="5" heatid="6832" entrytime="00:01:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-09-13" firstname="Piotr" gender="M" lastname="Kopiec" nation="POL" athleteid="2433">
              <RESULTS>
                <RESULT eventid="1696" points="274" reactiontime="+71" swimtime="00:01:30.64" resultid="2436" lane="8" heatid="7307" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.91" />
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                    <SPLIT distance="75" swimtime="00:01:03.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="253" reactiontime="+89" swimtime="00:03:21.58" resultid="2435" lane="3" heatid="7005" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.56" />
                    <SPLIT distance="50" swimtime="00:00:41.57" />
                    <SPLIT distance="75" swimtime="00:01:05.70" />
                    <SPLIT distance="100" swimtime="00:01:31.45" />
                    <SPLIT distance="125" swimtime="00:01:58.46" />
                    <SPLIT distance="150" swimtime="00:02:26.33" />
                    <SPLIT distance="175" swimtime="00:02:54.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="353" reactiontime="+88" swimtime="00:00:38.43" resultid="2434" lane="2" heatid="6859" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MODAB" name="CSiR MOS Dąbrowa Górnicza" nation="POL" region="SLA">
          <CONTACT name="waliczek mariusz" phone="606448210" />
          <ATHLETES>
            <ATHLETE birthdate="1988-03-24" firstname="Kamil" gender="M" lastname="Samul" nation="POL" license="S02711200032" athleteid="2438">
              <RESULTS>
                <RESULT eventid="1375" points="632" reactiontime="+85" swimtime="00:04:16.36" resultid="2440" lane="4" heatid="6909" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.65" />
                    <SPLIT distance="50" swimtime="00:00:29.68" />
                    <SPLIT distance="75" swimtime="00:00:45.84" />
                    <SPLIT distance="100" swimtime="00:01:02.59" />
                    <SPLIT distance="125" swimtime="00:01:19.02" />
                    <SPLIT distance="150" swimtime="00:01:35.67" />
                    <SPLIT distance="175" swimtime="00:01:51.99" />
                    <SPLIT distance="200" swimtime="00:02:08.85" />
                    <SPLIT distance="225" swimtime="00:02:25.12" />
                    <SPLIT distance="250" swimtime="00:02:41.56" />
                    <SPLIT distance="275" swimtime="00:02:57.67" />
                    <SPLIT distance="300" swimtime="00:03:13.79" />
                    <SPLIT distance="325" swimtime="00:03:29.46" />
                    <SPLIT distance="350" swimtime="00:03:45.52" />
                    <SPLIT distance="375" swimtime="00:04:00.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="643" reactiontime="+83" swimtime="00:01:59.26" resultid="2441" lane="2" heatid="7066" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.88" />
                    <SPLIT distance="50" swimtime="00:00:27.49" />
                    <SPLIT distance="75" swimtime="00:00:42.55" />
                    <SPLIT distance="100" swimtime="00:00:58.01" />
                    <SPLIT distance="125" swimtime="00:01:13.19" />
                    <SPLIT distance="150" swimtime="00:01:28.92" />
                    <SPLIT distance="175" swimtime="00:01:44.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="609" reactiontime="+80" swimtime="00:00:55.48" resultid="2439" lane="1" heatid="6846" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.60" />
                    <SPLIT distance="50" swimtime="00:00:26.49" />
                    <SPLIT distance="75" swimtime="00:00:40.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="559" reactiontime="+79" swimtime="00:00:27.86" resultid="2442" lane="8" heatid="7294" entrytime="00:00:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="610" reactiontime="+71" swimtime="00:00:25.08" resultid="2443" lane="3" heatid="7353" entrytime="00:00:25.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TAKAS" name="Takas" nation="LTU">
          <CONTACT city="Kaunas" email="abicka@takas.lt" internet="www.klubastakas.lt" name="Romaldas Bickauskas" phone="+37068297778" street="Lentvario g. 19" zip="44439" />
          <ATHLETES>
            <ATHLETE birthdate="1927-04-21" firstname="Vladas" gender="M" lastname="VIMBARAS" nation="LTU" athleteid="2445">
              <RESULTS>
                <RESULT eventid="1496" points="33" reactiontime="+78" swimtime="00:01:15.67" resultid="2447" lane="8" heatid="7033" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="78" reactiontime="+104" swimtime="00:00:49.61" resultid="2448" lane="2" heatid="7336" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="43" reactiontime="+101" swimtime="00:02:14.22" resultid="2446" lane="2" heatid="6830" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.06" />
                    <SPLIT distance="50" swimtime="00:01:01.66" />
                    <SPLIT distance="75" swimtime="00:01:37.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-01-25" firstname="Dalicija" gender="F" lastname="FEDORAVICIENE" nation="LTU" athleteid="2449">
              <RESULTS>
                <RESULT eventid="1547" points="81" reactiontime="+115" swimtime="00:04:25.07" resultid="2451" heatid="7049" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.42" />
                    <SPLIT distance="50" swimtime="00:00:59.82" />
                    <SPLIT distance="75" swimtime="00:01:34.09" />
                    <SPLIT distance="100" swimtime="00:02:09.79" />
                    <SPLIT distance="125" swimtime="00:02:44.92" />
                    <SPLIT distance="150" swimtime="00:03:19.79" />
                    <SPLIT distance="175" swimtime="00:03:53.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="80" reactiontime="+117" swimtime="00:02:02.30" resultid="2450" lane="5" heatid="6822" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.89" />
                    <SPLIT distance="50" swimtime="00:00:57.91" />
                    <SPLIT distance="75" swimtime="00:01:30.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="96" reactiontime="+134" swimtime="00:00:52.21" resultid="2452" lane="8" heatid="7329" entrytime="00:00:54.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1945-09-25" firstname="Vytautas" gender="M" lastname="SVETIKAS" nation="LTU" athleteid="2453">
              <RESULTS>
                <RESULT eventid="1564" points="111" reactiontime="+102" swimtime="00:03:33.69" resultid="2455" lane="6" heatid="7055" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.70" />
                    <SPLIT distance="50" swimtime="00:00:45.02" />
                    <SPLIT distance="75" swimtime="00:01:11.27" />
                    <SPLIT distance="100" swimtime="00:01:39.14" />
                    <SPLIT distance="125" swimtime="00:02:08.17" />
                    <SPLIT distance="150" swimtime="00:02:37.16" />
                    <SPLIT distance="175" swimtime="00:03:06.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="210" reactiontime="+84" swimtime="00:00:35.77" resultid="2456" lane="6" heatid="7338" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="151" reactiontime="+112" swimtime="00:01:28.26" resultid="2454" lane="6" heatid="6832" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.07" />
                    <SPLIT distance="50" swimtime="00:00:40.12" />
                    <SPLIT distance="75" swimtime="00:01:03.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-11-16" firstname="Violeta" gender="F" lastname="POVILAITIENE" nation="LTU" athleteid="2457">
              <RESULTS>
                <RESULT eventid="1479" points="108" reactiontime="+87" swimtime="00:00:58.10" resultid="2459" lane="2" heatid="7026" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="134" reactiontime="+114" swimtime="00:00:59.15" resultid="2458" lane="2" heatid="6849" entrytime="00:00:53.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="101" reactiontime="+120" swimtime="00:00:51.42" resultid="2461" lane="1" heatid="7329" entrytime="00:00:49.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" status="DNS" swimtime="00:00:00.00" resultid="2460" lane="3" heatid="7275" entrytime="00:00:56.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-07-09" firstname="Antanas" gender="M" lastname="GUOGA" nation="LTU" athleteid="2462">
              <RESULTS>
                <RESULT eventid="1143" points="150" swimtime="00:27:22.55" resultid="2463" lane="2" heatid="6749" entrytime="00:28:00.00" />
                <RESULT eventid="1273" points="80" reactiontime="+112" swimtime="00:04:19.48" resultid="2464" lane="1" heatid="6870" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.63" />
                    <SPLIT distance="50" swimtime="00:00:57.54" />
                    <SPLIT distance="75" swimtime="00:01:28.45" />
                    <SPLIT distance="100" swimtime="00:02:01.03" />
                    <SPLIT distance="125" swimtime="00:02:33.87" />
                    <SPLIT distance="150" swimtime="00:03:09.15" />
                    <SPLIT distance="175" swimtime="00:03:43.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="110" reactiontime="+126" swimtime="00:03:58.13" resultid="2467" lane="5" heatid="7072" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.98" />
                    <SPLIT distance="50" swimtime="00:00:54.89" />
                    <SPLIT distance="75" swimtime="00:01:29.70" />
                    <SPLIT distance="100" swimtime="00:02:03.79" />
                    <SPLIT distance="125" swimtime="00:02:34.81" />
                    <SPLIT distance="150" swimtime="00:03:06.59" />
                    <SPLIT distance="175" swimtime="00:03:32.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="141" reactiontime="+107" swimtime="00:07:02.09" resultid="2465" lane="7" heatid="6900" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.98" />
                    <SPLIT distance="50" swimtime="00:00:43.81" />
                    <SPLIT distance="75" swimtime="00:01:08.92" />
                    <SPLIT distance="100" swimtime="00:01:34.67" />
                    <SPLIT distance="125" swimtime="00:02:01.27" />
                    <SPLIT distance="150" swimtime="00:02:28.36" />
                    <SPLIT distance="175" swimtime="00:02:55.80" />
                    <SPLIT distance="200" swimtime="00:03:23.09" />
                    <SPLIT distance="225" swimtime="00:03:50.48" />
                    <SPLIT distance="250" swimtime="00:04:18.14" />
                    <SPLIT distance="275" swimtime="00:04:46.24" />
                    <SPLIT distance="300" swimtime="00:05:13.69" />
                    <SPLIT distance="325" swimtime="00:05:41.99" />
                    <SPLIT distance="350" swimtime="00:06:09.49" />
                    <SPLIT distance="375" swimtime="00:06:36.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" status="DNS" swimtime="00:00:00.00" resultid="2468" lane="6" heatid="7303" entrytime="00:01:55.00" />
                <RESULT eventid="1411" status="DNS" swimtime="00:00:00.00" resultid="2466" lane="8" heatid="7004" entrytime="00:04:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-10-18" firstname="Ramune" gender="F" lastname="IVANAUSKAITE" nation="LTU" athleteid="2469">
              <RESULTS>
                <RESULT eventid="1058" points="306" swimtime="00:12:12.72" resultid="2470" heatid="6715" entrytime="00:12:10.00" />
                <RESULT eventid="1290" points="298" reactiontime="+85" swimtime="00:03:07.32" resultid="2471" lane="4" heatid="6878" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.56" />
                    <SPLIT distance="50" swimtime="00:00:43.90" />
                    <SPLIT distance="75" swimtime="00:01:06.91" />
                    <SPLIT distance="100" swimtime="00:01:30.80" />
                    <SPLIT distance="125" swimtime="00:01:54.77" />
                    <SPLIT distance="150" swimtime="00:02:19.24" />
                    <SPLIT distance="175" swimtime="00:02:43.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="312" reactiontime="+88" swimtime="00:05:55.79" resultid="2472" lane="7" heatid="6897" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.42" />
                    <SPLIT distance="50" swimtime="00:00:38.91" />
                    <SPLIT distance="75" swimtime="00:01:00.16" />
                    <SPLIT distance="100" swimtime="00:01:22.00" />
                    <SPLIT distance="125" swimtime="00:01:44.00" />
                    <SPLIT distance="150" swimtime="00:02:06.65" />
                    <SPLIT distance="175" swimtime="00:02:29.20" />
                    <SPLIT distance="200" swimtime="00:02:52.29" />
                    <SPLIT distance="225" swimtime="00:03:15.22" />
                    <SPLIT distance="250" swimtime="00:03:38.20" />
                    <SPLIT distance="275" swimtime="00:04:02.06" />
                    <SPLIT distance="300" swimtime="00:04:25.58" />
                    <SPLIT distance="325" swimtime="00:04:48.19" />
                    <SPLIT distance="350" swimtime="00:05:11.91" />
                    <SPLIT distance="375" swimtime="00:05:34.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="308" reactiontime="+79" swimtime="00:00:40.95" resultid="2473" lane="7" heatid="7030" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="309" swimtime="00:02:49.69" resultid="2474" lane="1" heatid="7052" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.96" />
                    <SPLIT distance="50" swimtime="00:00:38.39" />
                    <SPLIT distance="75" swimtime="00:00:59.42" />
                    <SPLIT distance="100" swimtime="00:01:21.05" />
                    <SPLIT distance="125" swimtime="00:01:43.30" />
                    <SPLIT distance="150" swimtime="00:02:05.68" />
                    <SPLIT distance="175" swimtime="00:02:28.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="306" reactiontime="+89" swimtime="00:01:27.18" resultid="2475" lane="1" heatid="7316" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.98" />
                    <SPLIT distance="50" swimtime="00:00:42.60" />
                    <SPLIT distance="75" swimtime="00:01:05.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-12-26" firstname="Arlandas" gender="M" lastname="JUODESKA" nation="LTU" athleteid="2476">
              <RESULTS>
                <RESULT eventid="1239" points="430" reactiontime="+82" swimtime="00:00:36.01" resultid="2478" lane="8" heatid="6862" entrytime="00:00:37.37">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="402" reactiontime="+76" swimtime="00:00:28.82" resultid="2481" lane="6" heatid="7345" entrytime="00:00:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="345" reactiontime="+67" swimtime="00:01:14.89" resultid="2480" lane="3" heatid="7323" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.25" />
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                    <SPLIT distance="75" swimtime="00:00:56.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="360" reactiontime="+70" swimtime="00:00:34.39" resultid="2479" lane="7" heatid="7040" entrytime="00:00:33.83">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="326" reactiontime="+83" swimtime="00:01:14.29" resultid="2477" lane="2" heatid="6740" entrytime="00:01:12.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.98" />
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                    <SPLIT distance="75" swimtime="00:00:55.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-08-03" firstname="Raimondas" gender="M" lastname="GARBATAVICIUS" nation="LTU" athleteid="2482">
              <RESULTS>
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="2483" lane="4" heatid="6740" entrytime="00:01:12.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-02-12" firstname="Irena" gender="F" lastname="JOKUBAITIENE" nation="LTU" athleteid="2485">
              <RESULTS>
                <RESULT eventid="1409" points="180" reactiontime="+104" swimtime="00:04:08.31" resultid="2487" lane="8" heatid="6999" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.39" />
                    <SPLIT distance="50" swimtime="00:00:55.41" />
                    <SPLIT distance="75" swimtime="00:01:26.05" />
                    <SPLIT distance="100" swimtime="00:01:58.18" />
                    <SPLIT distance="125" swimtime="00:02:30.62" />
                    <SPLIT distance="150" swimtime="00:03:03.03" />
                    <SPLIT distance="175" swimtime="00:03:35.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="183" reactiontime="+100" swimtime="00:01:54.54" resultid="2488" lane="7" heatid="7297" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.79" />
                    <SPLIT distance="50" swimtime="00:00:52.95" />
                    <SPLIT distance="75" swimtime="00:01:22.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="193" reactiontime="+103" swimtime="00:00:52.42" resultid="2486" lane="5" heatid="6849" entrytime="00:00:52.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-05-07" firstname="Jolanta" gender="F" lastname="Kozak" nation="LTU" athleteid="2489">
              <RESULTS>
                <RESULT eventid="1547" points="93" reactiontime="+106" swimtime="00:04:12.88" resultid="2493" lane="7" heatid="7049" entrytime="00:04:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.73" />
                    <SPLIT distance="50" swimtime="00:00:53.80" />
                    <SPLIT distance="75" swimtime="00:01:26.19" />
                    <SPLIT distance="100" swimtime="00:02:00.19" />
                    <SPLIT distance="125" swimtime="00:02:35.75" />
                    <SPLIT distance="150" swimtime="00:03:10.25" />
                    <SPLIT distance="175" swimtime="00:03:43.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="98" reactiontime="+79" swimtime="00:00:59.90" resultid="2492" lane="4" heatid="7025" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="104" reactiontime="+120" swimtime="00:01:52.21" resultid="2490" heatid="6823" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.86" />
                    <SPLIT distance="50" swimtime="00:00:53.05" />
                    <SPLIT distance="75" swimtime="00:01:24.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="103" reactiontime="+149" swimtime="00:00:50.99" resultid="2495" lane="7" heatid="7329" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.81" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="przekroczony limit 8:30:00" eventid="1358" reactiontime="+129" status="DSQ" swimtime="00:00:00.00" resultid="2491" lane="2" heatid="6894" entrytime="00:08:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.89" />
                    <SPLIT distance="50" swimtime="00:00:54.56" />
                    <SPLIT distance="75" swimtime="00:01:25.46" />
                    <SPLIT distance="100" swimtime="00:01:58.73" />
                    <SPLIT distance="125" swimtime="00:02:33.30" />
                    <SPLIT distance="150" swimtime="00:03:07.99" />
                    <SPLIT distance="175" swimtime="00:03:42.97" />
                    <SPLIT distance="200" swimtime="00:04:17.95" />
                    <SPLIT distance="225" swimtime="00:04:54.35" />
                    <SPLIT distance="250" swimtime="00:05:29.16" />
                    <SPLIT distance="275" swimtime="00:06:04.98" />
                    <SPLIT distance="300" swimtime="00:06:40.00" />
                    <SPLIT distance="325" swimtime="00:07:14.70" />
                    <SPLIT distance="350" swimtime="00:07:49.71" />
                    <SPLIT distance="375" swimtime="00:08:25.19" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G 8" eventid="1713" reactiontime="+129" status="DSQ" swimtime="00:00:00.00" resultid="2494" lane="5" heatid="7313" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:31.78" />
                    <SPLIT distance="50" swimtime="00:01:07.25" />
                    <SPLIT distance="75" swimtime="00:01:46.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1938-01-08" firstname="Pavelas" gender="M" lastname="Bezzubovas" nation="LTU" athleteid="2496">
              <RESULTS>
                <RESULT eventid="1645" points="204" reactiontime="+112" swimtime="00:00:38.98" resultid="2498" lane="1" heatid="7283" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="220" reactiontime="+106" swimtime="00:00:35.21" resultid="2499" lane="2" heatid="7338" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="142" reactiontime="+109" swimtime="00:01:37.95" resultid="2497" lane="5" heatid="6732" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.27" />
                    <SPLIT distance="50" swimtime="00:00:48.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-04-12" firstname="Aleksandra" gender="F" lastname="YLIENE" nation="LTU" athleteid="2500">
              <RESULTS>
                <RESULT eventid="1479" points="173" reactiontime="+84" swimtime="00:00:49.59" resultid="2503" lane="7" heatid="7027" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="137" reactiontime="+123" swimtime="00:07:48.25" resultid="2502" lane="3" heatid="6894" entrytime="00:07:52.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.51" />
                    <SPLIT distance="50" swimtime="00:00:49.14" />
                    <SPLIT distance="75" swimtime="00:01:17.69" />
                    <SPLIT distance="100" swimtime="00:01:46.97" />
                    <SPLIT distance="125" swimtime="00:02:16.95" />
                    <SPLIT distance="150" swimtime="00:02:46.53" />
                    <SPLIT distance="175" swimtime="00:03:16.75" />
                    <SPLIT distance="200" swimtime="00:03:46.70" />
                    <SPLIT distance="225" swimtime="00:04:16.41" />
                    <SPLIT distance="250" swimtime="00:04:47.28" />
                    <SPLIT distance="275" swimtime="00:05:17.61" />
                    <SPLIT distance="300" swimtime="00:05:47.65" />
                    <SPLIT distance="325" swimtime="00:06:17.94" />
                    <SPLIT distance="350" swimtime="00:06:48.07" />
                    <SPLIT distance="375" swimtime="00:07:17.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="127" reactiontime="+86" swimtime="00:04:08.59" resultid="2501" lane="5" heatid="6876" entrytime="00:04:24.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.40" />
                    <SPLIT distance="50" swimtime="00:00:55.52" />
                    <SPLIT distance="75" swimtime="00:01:27.20" />
                    <SPLIT distance="100" swimtime="00:01:59.47" />
                    <SPLIT distance="125" swimtime="00:02:32.67" />
                    <SPLIT distance="150" swimtime="00:03:06.06" />
                    <SPLIT distance="175" swimtime="00:03:38.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="132" reactiontime="+82" swimtime="00:01:55.36" resultid="2505" lane="6" heatid="7314" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.83" />
                    <SPLIT distance="50" swimtime="00:00:54.10" />
                    <SPLIT distance="75" swimtime="00:01:24.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" status="DNS" swimtime="00:00:00.00" resultid="2504" lane="2" heatid="7049" entrytime="00:03:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-06-14" firstname="Violeta" gender="F" lastname="KRAJAUSKIENE" nation="LTU" athleteid="2506">
              <RESULTS>
                <RESULT eventid="1581" points="114" reactiontime="+115" swimtime="00:04:24.80" resultid="2507" lane="4" heatid="7067" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.33" />
                    <SPLIT distance="50" swimtime="00:00:59.26" />
                    <SPLIT distance="75" swimtime="00:01:31.77" />
                    <SPLIT distance="100" swimtime="00:02:05.65" />
                    <SPLIT distance="125" swimtime="00:02:42.14" />
                    <SPLIT distance="150" swimtime="00:03:17.43" />
                    <SPLIT distance="175" swimtime="00:03:50.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="89" reactiontime="+99" swimtime="00:00:56.89" resultid="2508" lane="1" heatid="7276" entrytime="00:00:51.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1177" status="DNS" swimtime="00:00:00.00" resultid="6667" lane="1" heatid="6807">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2453" number="1" />
                    <RELAYPOSITION athleteid="2445" number="2" />
                    <RELAYPOSITION athleteid="2462" number="3" />
                    <RELAYPOSITION athleteid="2496" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="OROPO" name="ORS Opole" nation="POL" region="OPO">
          <CONTACT name="Waldemar Kania" phone="694299743" />
          <ATHLETES>
            <ATHLETE birthdate="1968-01-01" firstname="Grzegorz" gender="M" lastname="Stanek" nation="POL" athleteid="2510">
              <RESULTS>
                <RESULT comment="Rekord Polski " eventid="1205" points="559" reactiontime="+66" swimtime="00:00:57.10" resultid="2512" lane="3" heatid="6845" entrytime="00:00:57.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.98" />
                    <SPLIT distance="50" swimtime="00:00:27.43" />
                    <SPLIT distance="75" swimtime="00:00:42.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="511" reactiontime="+78" swimtime="00:02:08.77" resultid="2514" lane="5" heatid="7065" entrytime="00:02:08.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.97" />
                    <SPLIT distance="50" swimtime="00:00:30.24" />
                    <SPLIT distance="75" swimtime="00:00:46.86" />
                    <SPLIT distance="100" swimtime="00:01:03.56" />
                    <SPLIT distance="125" swimtime="00:01:20.24" />
                    <SPLIT distance="150" swimtime="00:01:36.88" />
                    <SPLIT distance="175" swimtime="00:01:53.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="477" reactiontime="+76" swimtime="00:01:05.44" resultid="2511" lane="5" heatid="6744" entrytime="00:01:04.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.31" />
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                    <SPLIT distance="75" swimtime="00:00:49.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" status="DNS" swimtime="00:00:00.00" resultid="2515" lane="2" heatid="7080" entrytime="00:02:21.60" />
                <RESULT eventid="1375" status="DNS" swimtime="00:00:00.00" resultid="2513" lane="1" heatid="6909" entrytime="00:04:33.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-01" firstname="Waldemar" gender="M" lastname="Kania" nation="POL" athleteid="2516">
              <RESULTS>
                <RESULT eventid="1375" points="307" reactiontime="+93" swimtime="00:05:26.12" resultid="2519" lane="5" heatid="6906" entrytime="00:05:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.20" />
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                    <SPLIT distance="75" swimtime="00:00:56.80" />
                    <SPLIT distance="100" swimtime="00:01:16.59" />
                    <SPLIT distance="125" swimtime="00:01:36.69" />
                    <SPLIT distance="150" swimtime="00:01:57.29" />
                    <SPLIT distance="175" swimtime="00:02:17.99" />
                    <SPLIT distance="200" swimtime="00:02:39.08" />
                    <SPLIT distance="225" swimtime="00:03:00.01" />
                    <SPLIT distance="250" swimtime="00:03:20.99" />
                    <SPLIT distance="275" swimtime="00:03:42.30" />
                    <SPLIT distance="300" swimtime="00:04:03.53" />
                    <SPLIT distance="325" swimtime="00:04:24.34" />
                    <SPLIT distance="350" swimtime="00:04:45.39" />
                    <SPLIT distance="375" swimtime="00:05:06.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="305" swimtime="00:21:38.99" resultid="2517" lane="4" heatid="6751" entrytime="00:21:30.00" />
                <RESULT eventid="1564" points="301" reactiontime="+93" swimtime="00:02:33.49" resultid="2520" lane="7" heatid="7062" entrytime="00:02:29.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.97" />
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                    <SPLIT distance="75" swimtime="00:00:53.29" />
                    <SPLIT distance="100" swimtime="00:01:12.95" />
                    <SPLIT distance="125" swimtime="00:01:33.21" />
                    <SPLIT distance="150" swimtime="00:01:53.82" />
                    <SPLIT distance="175" swimtime="00:02:14.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="314" reactiontime="+93" swimtime="00:01:09.20" resultid="2518" lane="6" heatid="6838" entrytime="00:01:08.35">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.70" />
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                    <SPLIT distance="75" swimtime="00:00:51.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Anna" gender="F" lastname="Dębińska" nation="POL" athleteid="2521">
              <RESULTS>
                <RESULT eventid="1222" points="444" reactiontime="+91" swimtime="00:00:39.72" resultid="2523" lane="1" heatid="6853" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1409" points="352" reactiontime="+90" swimtime="00:03:18.58" resultid="2525" lane="1" heatid="7001" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.19" />
                    <SPLIT distance="50" swimtime="00:00:41.66" />
                    <SPLIT distance="75" swimtime="00:01:06.21" />
                    <SPLIT distance="100" swimtime="00:01:31.45" />
                    <SPLIT distance="125" swimtime="00:01:57.25" />
                    <SPLIT distance="150" swimtime="00:02:24.27" />
                    <SPLIT distance="175" swimtime="00:02:51.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="371" reactiontime="+87" swimtime="00:01:21.76" resultid="2522" heatid="6729" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.10" />
                    <SPLIT distance="50" swimtime="00:00:38.19" />
                    <SPLIT distance="75" swimtime="00:01:01.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="361" reactiontime="+109" swimtime="00:00:38.83" resultid="2526" lane="8" heatid="7030" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="320" reactiontime="+106" swimtime="00:03:02.97" resultid="2524" lane="8" heatid="6878" entrytime="00:03:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.78" />
                    <SPLIT distance="50" swimtime="00:00:42.56" />
                    <SPLIT distance="75" swimtime="00:01:05.25" />
                    <SPLIT distance="100" swimtime="00:01:28.01" />
                    <SPLIT distance="125" swimtime="00:01:52.28" />
                    <SPLIT distance="150" swimtime="00:02:16.13" />
                    <SPLIT distance="175" swimtime="00:02:40.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WMWAR" name="Warsaw Masters Team" nation="POL" region="MAZ">
          <CONTACT city="Warszawa" email="jstobnic@gmail.com" internet="masters.waw.pl" name="Justyna Stobnicka" state="MAZ" street="¯ó³kiewskiego 40 m 11" zip="04-305" />
          <ATHLETES>
            <ATHLETE birthdate="1937-10-03" firstname="Ryszard" gender="M" lastname="Sielski" nation="POL" athleteid="2528">
              <RESULTS>
                <RESULT eventid="1075" points="79" swimtime="00:17:48.25" resultid="2529" lane="7" heatid="6717" entrytime="00:16:30.00" />
                <RESULT eventid="1798" points="81" reactiontime="+112" swimtime="00:09:21.29" resultid="2535" lane="8" heatid="7358" entrytime="00:08:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.53" />
                    <SPLIT distance="50" swimtime="00:01:08.04" />
                    <SPLIT distance="75" swimtime="00:01:45.93" />
                    <SPLIT distance="100" swimtime="00:02:26.56" />
                    <SPLIT distance="125" swimtime="00:03:04.08" />
                    <SPLIT distance="150" swimtime="00:03:40.90" />
                    <SPLIT distance="175" swimtime="00:04:16.49" />
                    <SPLIT distance="200" swimtime="00:04:51.55" />
                    <SPLIT distance="225" swimtime="00:05:27.30" />
                    <SPLIT distance="250" swimtime="00:06:01.92" />
                    <SPLIT distance="275" swimtime="00:06:38.52" />
                    <SPLIT distance="300" swimtime="00:07:13.89" />
                    <SPLIT distance="325" swimtime="00:07:43.99" />
                    <SPLIT distance="350" swimtime="00:08:16.61" />
                    <SPLIT distance="375" swimtime="00:08:48.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="81" reactiontime="+80" swimtime="00:04:22.39" resultid="2531" lane="5" heatid="6881" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.77" />
                    <SPLIT distance="50" swimtime="00:01:01.21" />
                    <SPLIT distance="75" swimtime="00:01:33.44" />
                    <SPLIT distance="100" swimtime="00:02:06.25" />
                    <SPLIT distance="125" swimtime="00:02:40.06" />
                    <SPLIT distance="150" swimtime="00:03:14.82" />
                    <SPLIT distance="175" swimtime="00:03:49.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="77" reactiontime="+110" swimtime="00:04:27.75" resultid="2533" heatid="7072" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.38" />
                    <SPLIT distance="50" swimtime="00:01:03.83" />
                    <SPLIT distance="75" swimtime="00:01:38.16" />
                    <SPLIT distance="100" swimtime="00:02:13.50" />
                    <SPLIT distance="125" swimtime="00:02:48.17" />
                    <SPLIT distance="150" swimtime="00:03:23.30" />
                    <SPLIT distance="175" swimtime="00:03:56.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="74" reactiontime="+77" swimtime="00:02:05.01" resultid="2534" lane="8" heatid="7319" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.74" />
                    <SPLIT distance="50" swimtime="00:01:01.12" />
                    <SPLIT distance="75" swimtime="00:01:33.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="45" reactiontime="+115" swimtime="00:05:14.39" resultid="2530" lane="6" heatid="6869" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.85" />
                    <SPLIT distance="50" swimtime="00:01:11.40" />
                    <SPLIT distance="75" swimtime="00:01:50.94" />
                    <SPLIT distance="100" swimtime="00:02:31.99" />
                    <SPLIT distance="125" swimtime="00:03:11.77" />
                    <SPLIT distance="150" swimtime="00:03:52.63" />
                    <SPLIT distance="175" swimtime="00:04:34.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="113" reactiontime="+114" swimtime="00:04:23.07" resultid="2532" lane="2" heatid="7003" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.30" />
                    <SPLIT distance="50" swimtime="00:00:59.96" />
                    <SPLIT distance="75" swimtime="00:01:33.78" />
                    <SPLIT distance="100" swimtime="00:02:07.14" />
                    <SPLIT distance="125" swimtime="00:02:41.93" />
                    <SPLIT distance="150" swimtime="00:03:16.25" />
                    <SPLIT distance="175" swimtime="00:03:50.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-05-14" firstname="Wojciech" gender="M" lastname="Kałużyński" nation="POL" athleteid="2536">
              <RESULTS>
                <RESULT eventid="1730" points="231" reactiontime="+83" swimtime="00:01:25.62" resultid="2541" lane="1" heatid="7322" entrytime="00:01:27.21">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.97" />
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                    <SPLIT distance="75" swimtime="00:01:03.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="270" reactiontime="+82" swimtime="00:02:39.20" resultid="2540" lane="2" heatid="7060" entrytime="00:02:38.44">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.27" />
                    <SPLIT distance="50" swimtime="00:00:34.91" />
                    <SPLIT distance="75" swimtime="00:00:54.39" />
                    <SPLIT distance="100" swimtime="00:01:14.88" />
                    <SPLIT distance="125" swimtime="00:01:35.79" />
                    <SPLIT distance="150" swimtime="00:01:57.71" />
                    <SPLIT distance="175" swimtime="00:02:18.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="246" reactiontime="+89" swimtime="00:05:51.16" resultid="2539" lane="4" heatid="6902" entrytime="00:06:00.59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.74" />
                    <SPLIT distance="50" swimtime="00:00:38.12" />
                    <SPLIT distance="75" swimtime="00:00:58.67" />
                    <SPLIT distance="100" swimtime="00:01:20.00" />
                    <SPLIT distance="125" swimtime="00:01:41.82" />
                    <SPLIT distance="150" swimtime="00:02:03.86" />
                    <SPLIT distance="175" swimtime="00:02:26.48" />
                    <SPLIT distance="200" swimtime="00:02:49.27" />
                    <SPLIT distance="225" swimtime="00:03:11.83" />
                    <SPLIT distance="250" swimtime="00:03:34.84" />
                    <SPLIT distance="275" swimtime="00:03:57.76" />
                    <SPLIT distance="300" swimtime="00:04:21.11" />
                    <SPLIT distance="325" swimtime="00:04:43.97" />
                    <SPLIT distance="350" swimtime="00:05:07.16" />
                    <SPLIT distance="375" swimtime="00:05:29.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="317" reactiontime="+90" swimtime="00:01:09.00" resultid="2538" lane="1" heatid="6838" entrytime="00:01:08.74">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.73" />
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                    <SPLIT distance="75" swimtime="00:00:49.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="226" reactiontime="+83" swimtime="00:01:23.94" resultid="2537" heatid="6736" entrytime="00:01:22.54">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.02" />
                    <SPLIT distance="50" swimtime="00:00:37.59" />
                    <SPLIT distance="75" swimtime="00:01:04.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="353" reactiontime="+83" swimtime="00:00:30.10" resultid="2542" lane="1" heatid="7343" entrytime="00:00:30.95">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-25" firstname="Marcin" gender="M" lastname="Kaczmarek" nation="POL" athleteid="2543">
              <RESULTS>
                <RESULT eventid="1496" points="643" reactiontime="+66" swimtime="00:00:28.34" resultid="2545" lane="3" heatid="7043" entrytime="00:00:27.27">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="646" reactiontime="+82" swimtime="00:00:58.28" resultid="2544" lane="2" heatid="7023" entrytime="00:00:58.58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.62" />
                    <SPLIT distance="50" swimtime="00:00:27.39" />
                    <SPLIT distance="75" swimtime="00:00:42.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="668" reactiontime="+80" swimtime="00:00:26.26" resultid="2546" lane="1" heatid="7294" entrytime="00:00:26.26">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="677" reactiontime="+65" swimtime="00:00:59.81" resultid="2547" lane="3" heatid="7326" entrytime="00:00:59.59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.33" />
                    <SPLIT distance="50" swimtime="00:00:29.71" />
                    <SPLIT distance="75" swimtime="00:00:45.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-10-02" firstname="Andrzej" gender="M" lastname="Wiszniewski" nation="POL" athleteid="2548">
              <RESULTS>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="2550" lane="6" heatid="6870" entrytime="00:03:58.30" />
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="2554" lane="6" heatid="7337" entrytime="00:00:39.65" />
                <RESULT eventid="1696" status="DNS" swimtime="00:00:00.00" resultid="2553" lane="7" heatid="7305" entrytime="00:01:38.90" />
                <RESULT eventid="1462" status="DNS" swimtime="00:00:00.00" resultid="2552" heatid="7016" entrytime="00:01:56.10" />
                <RESULT eventid="1411" status="DNS" swimtime="00:00:00.00" resultid="2551" lane="6" heatid="7005" entrytime="00:03:32.20" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="2549" lane="8" heatid="6856" entrytime="00:00:46.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-06-17" firstname="Leszek" gender="M" lastname="Madej" nation="POL" athleteid="2555">
              <RESULTS>
                <RESULT eventid="1205" points="540" reactiontime="+80" swimtime="00:00:57.75" resultid="2557" lane="6" heatid="6845" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.33" />
                    <SPLIT distance="50" swimtime="00:00:27.60" />
                    <SPLIT distance="75" swimtime="00:00:42.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="516" reactiontime="+78" swimtime="00:00:26.52" resultid="2559" lane="2" heatid="7350" entrytime="00:00:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="439" reactiontime="+80" swimtime="00:01:07.28" resultid="2556" lane="5" heatid="6743" entrytime="00:01:07.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.54" />
                    <SPLIT distance="50" swimtime="00:00:30.93" />
                    <SPLIT distance="75" swimtime="00:00:51.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="2558" lane="4" heatid="7064" entrytime="00:02:13.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-05" firstname="Rafał" gender="M" lastname="Skośkiewicz" nation="POL" athleteid="2560">
              <RESULTS>
                <RESULT eventid="1730" points="486" reactiontime="+73" swimtime="00:01:06.80" resultid="2566" heatid="7326" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.82" />
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                    <SPLIT distance="75" swimtime="00:00:49.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="433" reactiontime="+90" swimtime="00:01:07.56" resultid="2561" lane="7" heatid="6744" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.88" />
                    <SPLIT distance="50" swimtime="00:00:31.00" />
                    <SPLIT distance="75" swimtime="00:00:51.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="433" reactiontime="+70" swimtime="00:02:30.53" resultid="2563" lane="3" heatid="6886" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.29" />
                    <SPLIT distance="50" swimtime="00:00:34.12" />
                    <SPLIT distance="75" swimtime="00:00:53.25" />
                    <SPLIT distance="100" swimtime="00:01:12.67" />
                    <SPLIT distance="125" swimtime="00:01:32.12" />
                    <SPLIT distance="150" swimtime="00:01:51.89" />
                    <SPLIT distance="175" swimtime="00:02:11.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="397" reactiontime="+76" swimtime="00:00:33.27" resultid="2564" lane="2" heatid="7041" entrytime="00:00:31.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="410" reactiontime="+85" swimtime="00:00:36.57" resultid="2562" lane="1" heatid="6864" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="452" reactiontime="+83" swimtime="00:00:27.71" resultid="2567" lane="5" heatid="7346" entrytime="00:00:28.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" status="DNS" swimtime="00:00:00.00" resultid="2565" lane="8" heatid="7079" entrytime="00:02:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-09-25" firstname="Barbara" gender="F" lastname="Ropa" nation="POL" athleteid="2568">
              <RESULTS>
                <RESULT eventid="1126" points="270" swimtime="00:24:16.50" resultid="2569" lane="8" heatid="6747" entrytime="00:27:00.00" />
                <RESULT eventid="1781" points="244" reactiontime="+94" swimtime="00:07:10.82" resultid="2575" lane="1" heatid="7356" entrytime="00:07:08.03">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.53" />
                    <SPLIT distance="50" swimtime="00:00:45.78" />
                    <SPLIT distance="75" swimtime="00:01:13.31" />
                    <SPLIT distance="100" swimtime="00:01:41.13" />
                    <SPLIT distance="125" swimtime="00:02:13.19" />
                    <SPLIT distance="150" swimtime="00:02:42.93" />
                    <SPLIT distance="175" swimtime="00:03:12.10" />
                    <SPLIT distance="200" swimtime="00:03:41.29" />
                    <SPLIT distance="225" swimtime="00:04:09.95" />
                    <SPLIT distance="250" swimtime="00:04:38.15" />
                    <SPLIT distance="275" swimtime="00:05:06.72" />
                    <SPLIT distance="300" swimtime="00:05:35.39" />
                    <SPLIT distance="325" swimtime="00:06:00.98" />
                    <SPLIT distance="350" swimtime="00:06:25.96" />
                    <SPLIT distance="375" swimtime="00:06:49.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="276" reactiontime="+97" swimtime="00:06:10.58" resultid="2571" lane="4" heatid="6896" entrytime="00:06:05.15">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.15" />
                    <SPLIT distance="50" swimtime="00:00:42.37" />
                    <SPLIT distance="75" swimtime="00:01:05.55" />
                    <SPLIT distance="100" swimtime="00:01:28.92" />
                    <SPLIT distance="125" swimtime="00:01:52.60" />
                    <SPLIT distance="150" swimtime="00:02:16.24" />
                    <SPLIT distance="175" swimtime="00:02:40.22" />
                    <SPLIT distance="200" swimtime="00:03:03.94" />
                    <SPLIT distance="225" swimtime="00:03:27.80" />
                    <SPLIT distance="250" swimtime="00:03:51.75" />
                    <SPLIT distance="275" swimtime="00:04:15.54" />
                    <SPLIT distance="300" swimtime="00:04:39.21" />
                    <SPLIT distance="325" swimtime="00:05:02.86" />
                    <SPLIT distance="350" swimtime="00:05:26.70" />
                    <SPLIT distance="375" swimtime="00:05:49.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1409" points="292" reactiontime="+93" swimtime="00:03:31.13" resultid="2572" lane="5" heatid="7000" entrytime="00:03:24.18">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.47" />
                    <SPLIT distance="50" swimtime="00:00:46.88" />
                    <SPLIT distance="75" swimtime="00:01:13.21" />
                    <SPLIT distance="100" swimtime="00:01:39.98" />
                    <SPLIT distance="125" swimtime="00:02:07.77" />
                    <SPLIT distance="150" swimtime="00:02:35.73" />
                    <SPLIT distance="175" swimtime="00:03:03.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="294" reactiontime="+94" swimtime="00:01:37.88" resultid="2574" lane="3" heatid="7298" entrytime="00:01:41.08">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.82" />
                    <SPLIT distance="50" swimtime="00:00:46.71" />
                    <SPLIT distance="75" swimtime="00:01:12.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="310" reactiontime="+89" swimtime="00:00:44.75" resultid="2570" lane="6" heatid="6851" entrytime="00:00:45.06">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1581" status="DNS" swimtime="00:00:00.00" resultid="2573" lane="5" heatid="7069" entrytime="00:03:23.78" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-12-15" firstname="Jerzy" gender="M" lastname="Chrześcijański" nation="POL" athleteid="2576">
              <RESULTS>
                <RESULT eventid="1075" points="240" swimtime="00:12:17.68" resultid="2577" lane="4" heatid="6719" entrytime="00:12:13.00" />
                <RESULT eventid="1564" points="271" reactiontime="+80" swimtime="00:02:38.95" resultid="2580" lane="5" heatid="7059" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.63" />
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                    <SPLIT distance="75" swimtime="00:00:54.90" />
                    <SPLIT distance="100" swimtime="00:01:15.49" />
                    <SPLIT distance="125" swimtime="00:01:36.24" />
                    <SPLIT distance="150" swimtime="00:01:57.83" />
                    <SPLIT distance="175" swimtime="00:02:18.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="246" reactiontime="+72" swimtime="00:05:51.22" resultid="2579" lane="5" heatid="6904" entrytime="00:05:49.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.41" />
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                    <SPLIT distance="75" swimtime="00:01:01.88" />
                    <SPLIT distance="100" swimtime="00:01:24.04" />
                    <SPLIT distance="125" swimtime="00:01:46.76" />
                    <SPLIT distance="150" swimtime="00:02:09.46" />
                    <SPLIT distance="175" swimtime="00:02:31.73" />
                    <SPLIT distance="200" swimtime="00:02:54.71" />
                    <SPLIT distance="225" swimtime="00:03:17.58" />
                    <SPLIT distance="250" swimtime="00:03:40.01" />
                    <SPLIT distance="275" swimtime="00:04:02.64" />
                    <SPLIT distance="300" swimtime="00:04:25.23" />
                    <SPLIT distance="325" swimtime="00:04:47.50" />
                    <SPLIT distance="350" swimtime="00:05:09.50" />
                    <SPLIT distance="375" swimtime="00:05:31.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="261" reactiontime="+79" swimtime="00:01:13.60" resultid="2578" lane="5" heatid="6834" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.50" />
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                    <SPLIT distance="75" swimtime="00:00:54.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-02-29" firstname="Jan Maciej" gender="M" lastname="Boboli" nation="POL" athleteid="2581">
              <RESULTS>
                <RESULT eventid="1645" points="193" reactiontime="+85" swimtime="00:00:39.69" resultid="2586" lane="8" heatid="7284" entrytime="00:00:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="73" reactiontime="+92" swimtime="00:01:04.93" resultid="2584" lane="4" heatid="6854" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="208" reactiontime="+81" swimtime="00:00:35.86" resultid="2587" heatid="7340" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="160" reactiontime="+95" swimtime="00:01:26.52" resultid="2583" lane="7" heatid="6832" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.82" />
                    <SPLIT distance="50" swimtime="00:00:40.41" />
                    <SPLIT distance="75" swimtime="00:01:03.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="94" reactiontime="+69" swimtime="00:00:53.64" resultid="2585" heatid="7034" entrytime="00:00:53.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="68" reactiontime="+84" swimtime="00:02:05.20" resultid="2582" lane="2" heatid="6731" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.32" />
                    <SPLIT distance="50" swimtime="00:00:49.45" />
                    <SPLIT distance="75" swimtime="00:01:37.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-04-22" firstname="Karol" gender="M" lastname="Dzięcioł" nation="POL" athleteid="2588">
              <RESULTS>
                <RESULT eventid="1205" points="574" reactiontime="+74" swimtime="00:00:56.60" resultid="2589" lane="2" heatid="6845" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.91" />
                    <SPLIT distance="50" swimtime="00:00:27.46" />
                    <SPLIT distance="75" swimtime="00:00:41.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="515" reactiontime="+75" swimtime="00:02:08.39" resultid="2590" lane="7" heatid="7065" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.63" />
                    <SPLIT distance="50" swimtime="00:00:28.94" />
                    <SPLIT distance="75" swimtime="00:00:45.03" />
                    <SPLIT distance="100" swimtime="00:01:01.67" />
                    <SPLIT distance="125" swimtime="00:01:18.49" />
                    <SPLIT distance="150" swimtime="00:01:35.42" />
                    <SPLIT distance="175" swimtime="00:01:52.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="457" reactiontime="+75" swimtime="00:02:28.30" resultid="2591" lane="4" heatid="7078" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.84" />
                    <SPLIT distance="50" swimtime="00:00:30.50" />
                    <SPLIT distance="75" swimtime="00:00:50.69" />
                    <SPLIT distance="100" swimtime="00:01:09.85" />
                    <SPLIT distance="125" swimtime="00:01:32.21" />
                    <SPLIT distance="150" swimtime="00:01:54.39" />
                    <SPLIT distance="175" swimtime="00:02:12.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="556" reactiontime="+74" swimtime="00:00:25.87" resultid="2592" lane="1" heatid="7352" entrytime="00:00:26.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-02-17" firstname="Robert" gender="M" lastname="Nowicki" nation="POL" athleteid="2593">
              <RESULTS>
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="2597" lane="2" heatid="7337" entrytime="00:00:39.00" />
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="2596" lane="8" heatid="7056" entrytime="00:03:20.00" />
                <RESULT eventid="1375" status="DNS" swimtime="00:00:00.00" resultid="2595" lane="7" heatid="6901" entrytime="00:07:00.00" />
                <RESULT comment="przekroczony limit 14:15:00" eventid="1075" status="DSQ" swimtime="00:15:16.75" resultid="2594" lane="3" heatid="6717" entrytime="00:14:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-06-02" firstname="Wojciech" gender="M" lastname="Czupryn" nation="POL" athleteid="2598">
              <RESULTS>
                <RESULT eventid="1075" points="159" swimtime="00:14:04.99" resultid="2599" lane="4" heatid="6717" entrytime="00:14:09.65" />
                <RESULT eventid="1411" points="168" reactiontime="+107" swimtime="00:03:50.98" resultid="2602" lane="4" heatid="7004" entrytime="00:03:48.94">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.97" />
                    <SPLIT distance="50" swimtime="00:00:53.67" />
                    <SPLIT distance="75" swimtime="00:01:22.41" />
                    <SPLIT distance="100" swimtime="00:01:51.04" />
                    <SPLIT distance="125" swimtime="00:02:20.72" />
                    <SPLIT distance="150" swimtime="00:02:50.59" />
                    <SPLIT distance="175" swimtime="00:03:21.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="181" reactiontime="+89" swimtime="00:03:01.83" resultid="2603" lane="6" heatid="7057" entrytime="00:02:57.99">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.48" />
                    <SPLIT distance="50" swimtime="00:00:39.61" />
                    <SPLIT distance="75" swimtime="00:01:02.23" />
                    <SPLIT distance="100" swimtime="00:01:26.04" />
                    <SPLIT distance="125" swimtime="00:01:49.83" />
                    <SPLIT distance="150" swimtime="00:02:13.96" />
                    <SPLIT distance="175" swimtime="00:02:38.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="168" reactiontime="+87" swimtime="00:00:41.60" resultid="2604" lane="6" heatid="7282" entrytime="00:00:44.64">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="223" reactiontime="+87" swimtime="00:01:17.55" resultid="2600" lane="8" heatid="6834" entrytime="00:01:18.17">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.59" />
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                    <SPLIT distance="75" swimtime="00:00:57.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="250" reactiontime="+82" swimtime="00:00:33.74" resultid="2605" lane="4" heatid="7339" entrytime="00:00:34.08">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="177" reactiontime="+103" swimtime="00:06:31.91" resultid="2601" lane="8" heatid="6902" entrytime="00:06:28.18">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.06" />
                    <SPLIT distance="50" swimtime="00:00:43.13" />
                    <SPLIT distance="75" swimtime="00:01:06.21" />
                    <SPLIT distance="100" swimtime="00:01:30.75" />
                    <SPLIT distance="125" swimtime="00:01:55.49" />
                    <SPLIT distance="150" swimtime="00:02:20.48" />
                    <SPLIT distance="175" swimtime="00:02:45.59" />
                    <SPLIT distance="200" swimtime="00:03:10.84" />
                    <SPLIT distance="225" swimtime="00:03:36.17" />
                    <SPLIT distance="250" swimtime="00:04:01.99" />
                    <SPLIT distance="275" swimtime="00:04:27.25" />
                    <SPLIT distance="300" swimtime="00:04:52.88" />
                    <SPLIT distance="325" swimtime="00:05:18.24" />
                    <SPLIT distance="350" swimtime="00:05:43.61" />
                    <SPLIT distance="375" swimtime="00:06:08.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1935-06-16" firstname="Elżbieta" gender="F" lastname="Janik" nation="POL" athleteid="2606">
              <RESULTS>
                <RESULT eventid="1290" points="69" reactiontime="+72" swimtime="00:05:05.01" resultid="2607" lane="1" heatid="6876" entrytime="00:04:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.63" />
                    <SPLIT distance="50" swimtime="00:01:11.98" />
                    <SPLIT distance="75" swimtime="00:01:50.34" />
                    <SPLIT distance="100" swimtime="00:02:29.33" />
                    <SPLIT distance="125" swimtime="00:03:07.77" />
                    <SPLIT distance="150" swimtime="00:03:47.76" />
                    <SPLIT distance="175" swimtime="00:04:27.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="66" reactiontime="+99" swimtime="00:01:08.31" resultid="2608" lane="3" heatid="7025" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="61" reactiontime="+72" swimtime="00:02:28.96" resultid="2609" lane="2" heatid="7313" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.68" />
                    <SPLIT distance="50" swimtime="00:01:12.20" />
                    <SPLIT distance="75" swimtime="00:01:51.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1964-08-01" firstname="Edyta" gender="F" lastname="Olszewska" nation="POL" athleteid="2610">
              <RESULTS>
                <RESULT eventid="1409" points="365" reactiontime="+78" swimtime="00:03:16.07" resultid="2613" lane="3" heatid="7001" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.70" />
                    <SPLIT distance="50" swimtime="00:00:42.68" />
                    <SPLIT distance="75" swimtime="00:01:06.63" />
                    <SPLIT distance="100" swimtime="00:01:31.67" />
                    <SPLIT distance="125" swimtime="00:01:57.55" />
                    <SPLIT distance="150" swimtime="00:02:23.53" />
                    <SPLIT distance="175" swimtime="00:02:50.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="395" reactiontime="+79" swimtime="00:01:28.69" resultid="2614" lane="2" heatid="7300" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.39" />
                    <SPLIT distance="50" swimtime="00:00:40.60" />
                    <SPLIT distance="75" swimtime="00:01:03.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="438" reactiontime="+79" swimtime="00:00:39.90" resultid="2612" lane="7" heatid="6853" entrytime="00:00:39.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="348" reactiontime="+79" swimtime="00:01:23.58" resultid="2611" lane="8" heatid="6728" entrytime="00:01:24.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.78" />
                    <SPLIT distance="50" swimtime="00:00:39.02" />
                    <SPLIT distance="75" swimtime="00:01:02.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1969-04-17" firstname="Andrzej" gender="M" lastname="Skorykow" nation="POL" athleteid="2615">
              <RESULTS>
                <RESULT eventid="1075" points="542" swimtime="00:09:22.36" resultid="2616" lane="5" heatid="6722" entrytime="00:09:37.50" />
                <RESULT eventid="1307" points="528" reactiontime="+62" swimtime="00:02:20.92" resultid="2617" lane="6" heatid="6887" entrytime="00:02:23.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.50" />
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                    <SPLIT distance="75" swimtime="00:00:51.17" />
                    <SPLIT distance="100" swimtime="00:01:09.15" />
                    <SPLIT distance="125" swimtime="00:01:27.39" />
                    <SPLIT distance="150" swimtime="00:01:45.65" />
                    <SPLIT distance="175" swimtime="00:02:03.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="521" reactiontime="+72" swimtime="00:01:02.61" resultid="2618" lane="1" heatid="7023" entrytime="00:01:01.45">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.08" />
                    <SPLIT distance="50" swimtime="00:00:28.96" />
                    <SPLIT distance="75" swimtime="00:00:45.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="553" reactiontime="+62" swimtime="00:01:03.99" resultid="2621" lane="6" heatid="7326" entrytime="00:01:04.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.73" />
                    <SPLIT distance="50" swimtime="00:00:30.76" />
                    <SPLIT distance="75" swimtime="00:00:47.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="588" reactiontime="+71" swimtime="00:00:27.40" resultid="2620" lane="3" heatid="7293" entrytime="00:00:27.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.65" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Zawodnik został ukarany żółtą kartą za niesportowe zachowanie." eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="2619" heatid="7066" entrytime="00:02:04.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-30" firstname="Monika" gender="F" lastname="Jarecka" nation="POL" athleteid="2622">
              <RESULTS>
                <RESULT eventid="1222" points="494" reactiontime="+80" swimtime="00:00:38.32" resultid="2624" lane="5" heatid="6853" entrytime="00:00:37.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="464" reactiontime="+76" swimtime="00:01:24.06" resultid="2626" lane="5" heatid="7300" entrytime="00:01:25.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.38" />
                    <SPLIT distance="50" swimtime="00:00:39.41" />
                    <SPLIT distance="75" swimtime="00:01:01.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1409" points="451" reactiontime="+85" swimtime="00:03:02.79" resultid="2625" lane="5" heatid="7001" entrytime="00:03:06.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.03" />
                    <SPLIT distance="50" swimtime="00:00:41.61" />
                    <SPLIT distance="75" swimtime="00:01:04.55" />
                    <SPLIT distance="100" swimtime="00:01:27.19" />
                    <SPLIT distance="125" swimtime="00:01:50.53" />
                    <SPLIT distance="150" swimtime="00:02:14.01" />
                    <SPLIT distance="175" swimtime="00:02:37.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="398" reactiontime="+79" swimtime="00:01:19.88" resultid="2623" lane="7" heatid="6728" entrytime="00:01:22.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.76" />
                    <SPLIT distance="50" swimtime="00:00:37.88" />
                    <SPLIT distance="75" swimtime="00:01:00.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="427" reactiontime="+78" swimtime="00:00:31.82" resultid="2627" lane="6" heatid="7334" entrytime="00:00:31.57">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-05-10" firstname="Michał" gender="M" lastname="Rudziński" nation="POL" athleteid="2628">
              <RESULTS>
                <RESULT eventid="1496" points="76" reactiontime="+101" swimtime="00:00:57.72" resultid="2632" lane="2" heatid="7033" entrytime="00:00:55.33">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="191" reactiontime="+112" swimtime="00:03:41.19" resultid="2631" heatid="7004" entrytime="00:03:55.18">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.22" />
                    <SPLIT distance="50" swimtime="00:00:49.68" />
                    <SPLIT distance="75" swimtime="00:01:16.61" />
                    <SPLIT distance="100" swimtime="00:01:45.29" />
                    <SPLIT distance="125" swimtime="00:02:13.78" />
                    <SPLIT distance="150" swimtime="00:02:43.10" />
                    <SPLIT distance="175" swimtime="00:03:12.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="99" reactiontime="+116" swimtime="00:01:41.40" resultid="2629" lane="7" heatid="6831" entrytime="00:01:40.19">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.20" />
                    <SPLIT distance="50" swimtime="00:00:48.60" />
                    <SPLIT distance="75" swimtime="00:01:16.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="182" reactiontime="+124" swimtime="00:00:47.95" resultid="2630" lane="4" heatid="6855" entrytime="00:00:48.94">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-11-07" firstname="Andrzej" gender="M" lastname="Lewandowski" nation="POL" athleteid="2633">
              <RESULTS>
                <RESULT eventid="1239" points="398" reactiontime="+88" swimtime="00:00:36.93" resultid="2634" lane="2" heatid="6861" entrytime="00:00:37.65">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="326" reactiontime="+84" swimtime="00:01:25.56" resultid="2636" lane="6" heatid="7307" entrytime="00:01:28.37">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.48" />
                    <SPLIT distance="50" swimtime="00:00:40.15" />
                    <SPLIT distance="75" swimtime="00:01:02.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="291" reactiontime="+87" swimtime="00:03:12.37" resultid="2635" lane="6" heatid="7006" entrytime="00:03:29.87">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.17" />
                    <SPLIT distance="50" swimtime="00:00:42.05" />
                    <SPLIT distance="75" swimtime="00:01:06.50" />
                    <SPLIT distance="100" swimtime="00:01:31.77" />
                    <SPLIT distance="125" swimtime="00:01:57.90" />
                    <SPLIT distance="150" swimtime="00:02:23.58" />
                    <SPLIT distance="175" swimtime="00:02:49.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="316" reactiontime="+89" swimtime="00:00:31.21" resultid="2637" lane="6" heatid="7342" entrytime="00:00:31.24">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-28" firstname="Monika" gender="F" lastname="Figura" nation="POL" athleteid="2638">
              <RESULTS>
                <RESULT eventid="1547" points="309" reactiontime="+97" swimtime="00:02:49.76" resultid="2641" lane="6" heatid="7052" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.56" />
                    <SPLIT distance="50" swimtime="00:00:38.39" />
                    <SPLIT distance="75" swimtime="00:00:58.93" />
                    <SPLIT distance="100" swimtime="00:01:20.92" />
                    <SPLIT distance="125" swimtime="00:01:43.31" />
                    <SPLIT distance="150" swimtime="00:02:05.60" />
                    <SPLIT distance="175" swimtime="00:02:29.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="414" reactiontime="+89" swimtime="00:00:32.15" resultid="2642" lane="1" heatid="7332" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="414" reactiontime="+85" swimtime="00:00:37.12" resultid="2640" lane="2" heatid="7028" entrytime="00:00:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="379" reactiontime="+90" swimtime="00:01:13.05" resultid="2639" lane="1" heatid="6826" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.20" />
                    <SPLIT distance="50" swimtime="00:00:35.87" />
                    <SPLIT distance="75" swimtime="00:00:54.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-03-04" firstname="Stefan" gender="M" lastname="Borodziuk" nation="POL" athleteid="2643">
              <RESULTS>
                <RESULT eventid="1375" points="125" reactiontime="+99" swimtime="00:07:19.65" resultid="2646" lane="5" heatid="6900" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.31" />
                    <SPLIT distance="50" swimtime="00:00:44.36" />
                    <SPLIT distance="75" swimtime="00:01:10.74" />
                    <SPLIT distance="100" swimtime="00:01:38.08" />
                    <SPLIT distance="125" swimtime="00:02:07.07" />
                    <SPLIT distance="150" swimtime="00:02:35.91" />
                    <SPLIT distance="175" swimtime="00:03:04.44" />
                    <SPLIT distance="200" swimtime="00:03:32.52" />
                    <SPLIT distance="225" swimtime="00:04:01.04" />
                    <SPLIT distance="250" swimtime="00:04:29.68" />
                    <SPLIT distance="275" swimtime="00:04:58.12" />
                    <SPLIT distance="300" swimtime="00:05:26.89" />
                    <SPLIT distance="325" swimtime="00:05:54.73" />
                    <SPLIT distance="350" swimtime="00:06:24.04" />
                    <SPLIT distance="375" swimtime="00:06:52.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="123" swimtime="00:15:19.81" resultid="2644" lane="1" heatid="6717" entrytime="00:15:30.00" />
                <RESULT eventid="1564" points="152" reactiontime="+95" swimtime="00:03:12.88" resultid="2648" heatid="7056" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.61" />
                    <SPLIT distance="50" swimtime="00:00:41.69" />
                    <SPLIT distance="75" swimtime="00:01:05.57" />
                    <SPLIT distance="100" swimtime="00:01:31.59" />
                    <SPLIT distance="125" swimtime="00:01:57.39" />
                    <SPLIT distance="150" swimtime="00:02:23.57" />
                    <SPLIT distance="175" swimtime="00:02:48.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="114" reactiontime="+74" swimtime="00:01:48.32" resultid="2649" lane="7" heatid="7320" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.43" />
                    <SPLIT distance="50" swimtime="00:00:52.08" />
                    <SPLIT distance="75" swimtime="00:01:20.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="186" reactiontime="+94" swimtime="00:01:22.34" resultid="2645" lane="4" heatid="6832" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.81" />
                    <SPLIT distance="50" swimtime="00:00:37.79" />
                    <SPLIT distance="75" swimtime="00:01:00.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="208" reactiontime="+72" swimtime="00:00:35.90" resultid="2650" lane="3" heatid="7338" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" status="DNS" swimtime="00:00:00.00" resultid="2647" lane="4" heatid="7034" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-12-31" firstname="Paweł" gender="M" lastname="Witkowski" nation="POL" athleteid="2651">
              <RESULTS>
                <RESULT eventid="1239" points="571" reactiontime="+81" swimtime="00:00:32.76" resultid="2652" lane="3" heatid="6865" entrytime="00:00:32.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" status="DNS" swimtime="00:00:00.00" resultid="2653" lane="5" heatid="7010" entrytime="00:02:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-03-16" firstname="Ewa" gender="F" lastname="Kosmol" nation="POL" athleteid="2654">
              <RESULTS>
                <RESULT eventid="1747" points="196" reactiontime="+103" swimtime="00:00:41.22" resultid="2658" lane="8" heatid="7330" entrytime="00:00:42.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="151" reactiontime="+90" swimtime="00:03:35.49" resultid="2657" lane="4" heatid="7049" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.91" />
                    <SPLIT distance="50" swimtime="00:00:49.17" />
                    <SPLIT distance="75" swimtime="00:01:16.41" />
                    <SPLIT distance="100" swimtime="00:01:43.69" />
                    <SPLIT distance="125" swimtime="00:02:11.65" />
                    <SPLIT distance="150" swimtime="00:02:40.44" />
                    <SPLIT distance="175" swimtime="00:03:08.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="173" reactiontime="+83" swimtime="00:01:45.42" resultid="2655" lane="4" heatid="6724" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.45" />
                    <SPLIT distance="50" swimtime="00:00:48.62" />
                    <SPLIT distance="75" swimtime="00:01:20.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="162" reactiontime="+92" swimtime="00:01:36.83" resultid="2656" lane="8" heatid="6824" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.84" />
                    <SPLIT distance="50" swimtime="00:00:46.87" />
                    <SPLIT distance="75" swimtime="00:01:12.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-12-31" firstname="Marianna" gender="F" lastname="Michalczyk" nation="POL" athleteid="2659">
              <RESULTS>
                <RESULT eventid="1581" points="313" reactiontime="+80" swimtime="00:03:09.02" resultid="2663" lane="1" heatid="7070" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.07" />
                    <SPLIT distance="50" swimtime="00:00:37.86" />
                    <SPLIT distance="75" swimtime="00:01:03.69" />
                    <SPLIT distance="100" swimtime="00:01:27.84" />
                    <SPLIT distance="125" swimtime="00:01:55.91" />
                    <SPLIT distance="150" swimtime="00:02:24.06" />
                    <SPLIT distance="175" swimtime="00:02:48.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1409" points="308" reactiontime="+84" swimtime="00:03:27.57" resultid="2662" lane="4" heatid="7000" entrytime="00:03:19.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.22" />
                    <SPLIT distance="50" swimtime="00:00:46.42" />
                    <SPLIT distance="75" swimtime="00:01:12.32" />
                    <SPLIT distance="100" swimtime="00:01:38.96" />
                    <SPLIT distance="125" swimtime="00:02:05.98" />
                    <SPLIT distance="150" swimtime="00:02:33.45" />
                    <SPLIT distance="175" swimtime="00:03:00.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="321" reactiontime="+81" swimtime="00:01:35.04" resultid="2665" heatid="7300" entrytime="00:01:32.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.58" />
                    <SPLIT distance="50" swimtime="00:00:44.78" />
                    <SPLIT distance="75" swimtime="00:01:09.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="335" reactiontime="+80" swimtime="00:00:43.62" resultid="2661" heatid="6852" entrytime="00:00:43.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="352" reactiontime="+83" swimtime="00:01:14.86" resultid="2660" lane="5" heatid="6826" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.78" />
                    <SPLIT distance="50" swimtime="00:00:35.92" />
                    <SPLIT distance="75" swimtime="00:00:55.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="353" reactiontime="+79" swimtime="00:00:36.01" resultid="2664" lane="7" heatid="7279" entrytime="00:00:35.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-13" firstname="Stanisław" gender="M" lastname="Kozak" nation="POL" athleteid="2666">
              <RESULTS>
                <RESULT eventid="1696" points="545" reactiontime="+83" swimtime="00:01:12.10" resultid="2670" lane="2" heatid="7311" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.92" />
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                    <SPLIT distance="75" swimtime="00:00:52.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="510" reactiontime="+91" swimtime="00:02:39.58" resultid="2669" lane="7" heatid="7011" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.54" />
                    <SPLIT distance="50" swimtime="00:00:35.07" />
                    <SPLIT distance="75" swimtime="00:00:55.87" />
                    <SPLIT distance="100" swimtime="00:01:16.92" />
                    <SPLIT distance="125" swimtime="00:01:38.11" />
                    <SPLIT distance="150" swimtime="00:01:59.48" />
                    <SPLIT distance="175" swimtime="00:02:19.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="635" reactiontime="+87" swimtime="00:00:31.62" resultid="2668" lane="3" heatid="6866" entrytime="00:00:30.88">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="391" reactiontime="+89" swimtime="00:01:09.90" resultid="2667" heatid="6741" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.94" />
                    <SPLIT distance="50" swimtime="00:00:36.19" />
                    <SPLIT distance="75" swimtime="00:00:53.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="469" reactiontime="+87" swimtime="00:00:27.38" resultid="2671" lane="3" heatid="7350" entrytime="00:00:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-07-26" firstname="Anna" gender="F" lastname="Szemberg" nation="POL" athleteid="2672">
              <RESULTS>
                <RESULT eventid="1358" points="150" reactiontime="+93" swimtime="00:07:34.05" resultid="2675" lane="8" heatid="6895" entrytime="00:07:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.40" />
                    <SPLIT distance="50" swimtime="00:00:50.19" />
                    <SPLIT distance="75" swimtime="00:01:18.48" />
                    <SPLIT distance="100" swimtime="00:01:46.80" />
                    <SPLIT distance="125" swimtime="00:02:16.04" />
                    <SPLIT distance="150" swimtime="00:02:45.02" />
                    <SPLIT distance="175" swimtime="00:03:14.55" />
                    <SPLIT distance="200" swimtime="00:04:42.88" />
                    <SPLIT distance="225" swimtime="00:04:14.22" />
                    <SPLIT distance="250" swimtime="00:05:41.70" />
                    <SPLIT distance="275" swimtime="00:05:12.02" />
                    <SPLIT distance="300" swimtime="00:06:40.18" />
                    <SPLIT distance="325" swimtime="00:06:11.02" />
                    <SPLIT distance="375" swimtime="00:07:08.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1058" points="143" swimtime="00:15:44.34" resultid="2673" lane="8" heatid="6714" entrytime="00:15:45.00" />
                <RESULT eventid="1547" points="147" reactiontime="+91" swimtime="00:03:37.18" resultid="2676" lane="3" heatid="7049" entrytime="00:03:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.47" />
                    <SPLIT distance="50" swimtime="00:00:47.53" />
                    <SPLIT distance="75" swimtime="00:01:15.39" />
                    <SPLIT distance="100" swimtime="00:01:44.01" />
                    <SPLIT distance="125" swimtime="00:02:13.67" />
                    <SPLIT distance="150" swimtime="00:02:42.17" />
                    <SPLIT distance="175" swimtime="00:03:11.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="140" reactiontime="+95" swimtime="00:01:41.69" resultid="2674" lane="3" heatid="6823" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.80" />
                    <SPLIT distance="50" swimtime="00:00:47.37" />
                    <SPLIT distance="75" swimtime="00:01:14.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="168" reactiontime="+96" swimtime="00:00:43.40" resultid="2677" lane="5" heatid="7329" entrytime="00:00:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-05" firstname="Arkadiusz" gender="M" lastname="Dobrzyński" nation="POL" athleteid="2678">
              <RESULTS>
                <RESULT eventid="1730" points="433" reactiontime="+70" swimtime="00:01:09.43" resultid="2683" lane="2" heatid="7325" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.55" />
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                    <SPLIT distance="75" swimtime="00:00:51.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="501" reactiontime="+81" swimtime="00:00:26.79" resultid="2684" heatid="7352" entrytime="00:00:26.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="373" reactiontime="+73" swimtime="00:02:38.22" resultid="2681" lane="1" heatid="6886" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.40" />
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                    <SPLIT distance="75" swimtime="00:00:55.30" />
                    <SPLIT distance="100" swimtime="00:01:15.15" />
                    <SPLIT distance="125" swimtime="00:01:35.65" />
                    <SPLIT distance="150" swimtime="00:01:56.37" />
                    <SPLIT distance="175" swimtime="00:02:17.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="449" reactiontime="+92" swimtime="00:01:01.42" resultid="2680" lane="3" heatid="6842" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.97" />
                    <SPLIT distance="50" swimtime="00:00:29.57" />
                    <SPLIT distance="75" swimtime="00:00:45.34" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="05" eventid="1496" reactiontime="+84" status="DSQ" swimtime="00:00:00.00" resultid="2682" lane="5" heatid="7041" entrytime="00:00:31.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="2679" lane="7" heatid="6741" entrytime="00:01:11.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-12-31" firstname="Ewa" gender="F" lastname="Krzyżanowska" nation="POL" athleteid="2685">
              <RESULTS>
                <RESULT eventid="1547" points="250" reactiontime="+106" swimtime="00:03:02.11" resultid="2688" lane="3" heatid="7051" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.94" />
                    <SPLIT distance="50" swimtime="00:00:39.24" />
                    <SPLIT distance="75" swimtime="00:01:01.68" />
                    <SPLIT distance="100" swimtime="00:01:24.50" />
                    <SPLIT distance="125" swimtime="00:01:48.64" />
                    <SPLIT distance="150" swimtime="00:02:12.95" />
                    <SPLIT distance="175" swimtime="00:02:37.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="317" reactiontime="+78" swimtime="00:00:40.55" resultid="2687" lane="7" heatid="7028" entrytime="00:00:44.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="299" reactiontime="+110" swimtime="00:01:19.08" resultid="2686" lane="8" heatid="6827" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.95" />
                    <SPLIT distance="50" swimtime="00:00:36.52" />
                    <SPLIT distance="75" swimtime="00:00:57.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="365" reactiontime="+94" swimtime="00:00:33.53" resultid="2690" lane="7" heatid="7334" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SUWAL" name="Suwałki" nation="POL">
          <CONTACT name="Obukowicz" />
          <ATHLETES>
            <ATHLETE birthdate="1985-09-23" firstname="Marcin" gender="M" lastname="Obukowicz" nation="POL" athleteid="2692">
              <RESULTS>
                <RESULT eventid="1411" points="366" reactiontime="+78" swimtime="00:02:58.18" resultid="2695" lane="8" heatid="7011" entrytime="00:02:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.42" />
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                    <SPLIT distance="75" swimtime="00:01:00.37" />
                    <SPLIT distance="100" swimtime="00:01:23.12" />
                    <SPLIT distance="125" swimtime="00:01:47.01" />
                    <SPLIT distance="150" swimtime="00:02:11.17" />
                    <SPLIT distance="175" swimtime="00:02:35.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="507" reactiontime="+77" swimtime="00:00:34.07" resultid="2693" lane="2" heatid="6865" entrytime="00:00:33.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="225" reactiontime="+83" swimtime="00:03:04.10" resultid="2694" lane="1" heatid="6873" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.25" />
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="75" swimtime="00:00:59.72" />
                    <SPLIT distance="100" swimtime="00:01:24.21" />
                    <SPLIT distance="125" swimtime="00:01:49.21" />
                    <SPLIT distance="150" swimtime="00:02:13.82" />
                    <SPLIT distance="175" swimtime="00:02:39.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" status="DNS" swimtime="00:00:00.00" resultid="2696" heatid="7364" entrytime="00:05:50.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LUBLI" name="Lublin" nation="POL" region="WIE">
          <CONTACT city="Lublin" email="kazik_s@o2.pl" name="Sinicki Kazimierz" phone="663728678" />
          <ATHLETES>
            <ATHLETE birthdate="1955-02-18" firstname="Kazimierz" gender="M" lastname="Sinicki" nation="POL" athleteid="3584">
              <RESULTS>
                <RESULT eventid="1645" points="372" reactiontime="+79" swimtime="00:00:31.90" resultid="3587" heatid="7288" entrytime="00:00:32.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="360" reactiontime="+87" swimtime="00:01:06.11" resultid="3585" lane="8" heatid="6841" entrytime="00:01:04.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.82" />
                    <SPLIT distance="50" swimtime="00:00:31.73" />
                    <SPLIT distance="75" swimtime="00:00:49.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="322" reactiontime="+83" swimtime="00:02:30.18" resultid="3586" lane="3" heatid="7061" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.33" />
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                    <SPLIT distance="75" swimtime="00:00:51.18" />
                    <SPLIT distance="100" swimtime="00:01:10.46" />
                    <SPLIT distance="125" swimtime="00:01:30.12" />
                    <SPLIT distance="150" swimtime="00:01:50.48" />
                    <SPLIT distance="175" swimtime="00:02:10.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="424" reactiontime="+77" swimtime="00:00:28.32" resultid="3588" heatid="7346" entrytime="00:00:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="REWRO" name="Redeco Wrocław" nation="POL" region="DOL">
          <CONTACT city="Wrocław" name="Wolny Dariusz" phone="603630870" state="DOL" street="Rogowska 52a" zip="54-440" />
          <ATHLETES>
            <ATHLETE birthdate="1960-03-21" firstname="Dariusz" gender="M" lastname="Wolny" nation="POL" athleteid="2705">
              <RESULTS>
                <RESULT comment="Rekord Polski " eventid="1109" points="468" reactiontime="+79" swimtime="00:01:05.88" resultid="2706" lane="1" heatid="6744" entrytime="00:01:06.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.82" />
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                    <SPLIT distance="75" swimtime="00:00:50.01" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1307" points="500" reactiontime="+71" swimtime="00:02:23.54" resultid="2707" lane="2" heatid="6887" entrytime="00:02:22.22">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.15" />
                    <SPLIT distance="50" swimtime="00:00:33.14" />
                    <SPLIT distance="75" swimtime="00:00:50.65" />
                    <SPLIT distance="100" swimtime="00:01:08.70" />
                    <SPLIT distance="125" swimtime="00:01:26.93" />
                    <SPLIT distance="150" swimtime="00:01:45.77" />
                    <SPLIT distance="175" swimtime="00:02:05.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="496" reactiontime="+71" swimtime="00:00:30.90" resultid="2708" lane="8" heatid="7042" entrytime="00:00:30.99">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="446" reactiontime="+79" swimtime="00:00:30.04" resultid="2710" lane="5" heatid="7291" entrytime="00:00:29.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="488" reactiontime="+70" swimtime="00:01:06.73" resultid="2711" lane="1" heatid="7326" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.71" />
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                    <SPLIT distance="75" swimtime="00:00:49.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" status="DNS" swimtime="00:00:00.00" resultid="2709" lane="8" heatid="7080" entrytime="00:02:26.26" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-10-05" firstname="Zbigniew" gender="M" lastname="Gałgański" nation="POL" athleteid="2712">
              <RESULTS>
                <RESULT eventid="1273" points="128" reactiontime="+99" swimtime="00:03:42.16" resultid="2714" heatid="6871" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.64" />
                    <SPLIT distance="50" swimtime="00:00:49.18" />
                    <SPLIT distance="75" swimtime="00:01:17.91" />
                    <SPLIT distance="100" swimtime="00:01:46.05" />
                    <SPLIT distance="125" swimtime="00:02:14.46" />
                    <SPLIT distance="150" swimtime="00:02:44.19" />
                    <SPLIT distance="175" swimtime="00:03:13.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="228" reactiontime="+93" swimtime="00:03:28.44" resultid="2715" lane="3" heatid="7006" entrytime="00:03:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.69" />
                    <SPLIT distance="50" swimtime="00:00:47.44" />
                    <SPLIT distance="75" swimtime="00:01:14.62" />
                    <SPLIT distance="100" swimtime="00:01:41.76" />
                    <SPLIT distance="125" swimtime="00:02:08.40" />
                    <SPLIT distance="150" swimtime="00:02:36.06" />
                    <SPLIT distance="175" swimtime="00:03:03.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="168" reactiontime="+90" swimtime="00:01:32.67" resultid="2713" lane="7" heatid="6734" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.31" />
                    <SPLIT distance="50" swimtime="00:00:45.68" />
                    <SPLIT distance="75" swimtime="00:01:11.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="174" reactiontime="+96" swimtime="00:00:41.06" resultid="2716" lane="5" heatid="7283" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" status="DNS" swimtime="00:00:00.00" resultid="2717" heatid="7360" entrytime="00:07:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-01" firstname="Maciej" gender="M" lastname="Chojcan" nation="POL" athleteid="2718">
              <RESULTS>
                <RESULT eventid="1205" points="321" reactiontime="+82" swimtime="00:01:08.70" resultid="2719" lane="1" heatid="6839" entrytime="00:01:07.23">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.35" />
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                    <SPLIT distance="75" swimtime="00:00:50.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="271" reactiontime="+80" swimtime="00:00:35.46" resultid="2720" lane="4" heatid="7287" entrytime="00:00:32.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="338" reactiontime="+80" swimtime="00:00:30.53" resultid="2721" lane="8" heatid="7345" entrytime="00:00:29.71">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-02-02" firstname="Joanna" gender="F" lastname="Chojcan" nation="POL" athleteid="2722">
              <RESULTS>
                <RESULT eventid="1581" points="407" reactiontime="+82" swimtime="00:02:53.30" resultid="2727" lane="5" heatid="7070" entrytime="00:02:47.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.44" />
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                    <SPLIT distance="75" swimtime="00:00:58.91" />
                    <SPLIT distance="100" swimtime="00:01:21.35" />
                    <SPLIT distance="125" swimtime="00:01:46.94" />
                    <SPLIT distance="150" swimtime="00:02:12.93" />
                    <SPLIT distance="175" swimtime="00:02:33.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="381" reactiontime="+80" swimtime="00:05:32.97" resultid="2725" heatid="6898" entrytime="00:05:20.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.34" />
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                    <SPLIT distance="75" swimtime="00:00:54.78" />
                    <SPLIT distance="100" swimtime="00:01:14.73" />
                    <SPLIT distance="125" swimtime="00:01:35.01" />
                    <SPLIT distance="150" swimtime="00:01:55.69" />
                    <SPLIT distance="175" swimtime="00:02:16.95" />
                    <SPLIT distance="200" swimtime="00:02:38.28" />
                    <SPLIT distance="225" swimtime="00:02:59.59" />
                    <SPLIT distance="250" swimtime="00:03:20.97" />
                    <SPLIT distance="275" swimtime="00:03:42.81" />
                    <SPLIT distance="300" swimtime="00:04:04.77" />
                    <SPLIT distance="325" swimtime="00:04:26.96" />
                    <SPLIT distance="350" swimtime="00:04:49.37" />
                    <SPLIT distance="375" swimtime="00:05:11.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="394" reactiontime="+67" swimtime="00:02:50.73" resultid="2724" lane="2" heatid="6879" entrytime="00:02:45.55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.78" />
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                    <SPLIT distance="75" swimtime="00:00:58.98" />
                    <SPLIT distance="100" swimtime="00:01:20.48" />
                    <SPLIT distance="125" swimtime="00:01:42.76" />
                    <SPLIT distance="150" swimtime="00:02:05.30" />
                    <SPLIT distance="175" swimtime="00:02:28.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="414" reactiontime="+70" swimtime="00:01:18.82" resultid="2729" lane="1" heatid="7317" entrytime="00:01:17.43">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.54" />
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                    <SPLIT distance="75" swimtime="00:00:58.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="390" reactiontime="+79" swimtime="00:00:34.82" resultid="2728" lane="3" heatid="7279" entrytime="00:00:34.42">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="440" reactiontime="+66" swimtime="00:00:36.37" resultid="2726" lane="7" heatid="7031" entrytime="00:00:35.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="405" reactiontime="+81" swimtime="00:01:19.43" resultid="2723" lane="7" heatid="6729" entrytime="00:01:18.22">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.49" />
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                    <SPLIT distance="75" swimtime="00:01:00.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-03-03" firstname="Małgorzata" gender="F" lastname="Bogdan" nation="POL" athleteid="2730">
              <RESULTS>
                <RESULT eventid="1256" points="166" reactiontime="+100" swimtime="00:03:45.61" resultid="2732" lane="2" heatid="6868" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.38" />
                    <SPLIT distance="50" swimtime="00:00:46.80" />
                    <SPLIT distance="75" swimtime="00:01:13.84" />
                    <SPLIT distance="100" swimtime="00:01:42.36" />
                    <SPLIT distance="125" swimtime="00:02:11.27" />
                    <SPLIT distance="150" swimtime="00:02:41.66" />
                    <SPLIT distance="175" swimtime="00:03:13.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="293" reactiontime="+78" swimtime="00:03:08.49" resultid="2733" lane="3" heatid="6878" entrytime="00:03:11.24">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.08" />
                    <SPLIT distance="50" swimtime="00:00:43.83" />
                    <SPLIT distance="75" swimtime="00:01:06.95" />
                    <SPLIT distance="100" swimtime="00:01:31.49" />
                    <SPLIT distance="125" swimtime="00:01:55.57" />
                    <SPLIT distance="150" swimtime="00:02:20.69" />
                    <SPLIT distance="175" swimtime="00:02:44.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="301" swimtime="00:01:27.73" resultid="2731" lane="2" heatid="6726" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.56" />
                    <SPLIT distance="50" swimtime="00:00:40.66" />
                    <SPLIT distance="75" swimtime="00:01:06.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-02-02" firstname="Piotr" gender="M" lastname="Maroń" nation="POL" athleteid="2734">
              <RESULTS>
                <RESULT eventid="1411" status="DNS" swimtime="00:00:00.00" resultid="2737" heatid="7007" entrytime="00:03:25.25" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="2736" lane="8" heatid="6861" entrytime="00:00:38.00" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="2735" lane="1" heatid="6837" entrytime="00:01:09.09" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-01-01" firstname="Jakub" gender="M" lastname="Piątkowski" nation="POL" athleteid="2738">
              <RESULTS>
                <RESULT eventid="1496" points="561" reactiontime="+64" swimtime="00:00:29.66" resultid="2742" lane="1" heatid="7043" entrytime="00:00:29.11">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="572" reactiontime="+80" swimtime="00:00:32.74" resultid="2740" heatid="6866" entrytime="00:00:32.32">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="480" reactiontime="+71" swimtime="00:02:25.45" resultid="2741" lane="5" heatid="6887" entrytime="00:02:20.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.16" />
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                    <SPLIT distance="75" swimtime="00:00:53.10" />
                    <SPLIT distance="100" swimtime="00:01:12.05" />
                    <SPLIT distance="125" swimtime="00:01:30.07" />
                    <SPLIT distance="150" swimtime="00:01:48.43" />
                    <SPLIT distance="175" swimtime="00:02:07.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="475" reactiontime="+85" swimtime="00:01:05.55" resultid="2739" lane="3" heatid="6744" entrytime="00:01:04.44">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.12" />
                    <SPLIT distance="50" swimtime="00:00:29.16" />
                    <SPLIT distance="75" swimtime="00:00:49.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="2743" lane="8" heatid="7065" entrytime="00:02:12.22" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-01" firstname="Przemysław" gender="M" lastname="Matuszek" nation="POL" athleteid="2744">
              <RESULTS>
                <RESULT eventid="1462" points="332" reactiontime="+78" swimtime="00:01:12.72" resultid="2748" lane="3" heatid="7019" entrytime="00:01:18.45">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.59" />
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                    <SPLIT distance="75" swimtime="00:00:51.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="424" reactiontime="+77" swimtime="00:00:30.54" resultid="2750" lane="7" heatid="7290" entrytime="00:00:30.58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="409" reactiontime="+76" swimtime="00:01:03.37" resultid="2746" lane="7" heatid="6839" entrytime="00:01:07.56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.61" />
                    <SPLIT distance="50" swimtime="00:00:28.99" />
                    <SPLIT distance="75" swimtime="00:00:45.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="388" reactiontime="+79" swimtime="00:00:37.24" resultid="2747" heatid="6862" entrytime="00:00:37.35">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="311" reactiontime="+74" swimtime="00:01:15.46" resultid="2745" lane="3" heatid="6738" entrytime="00:01:15.45">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.66" />
                    <SPLIT distance="50" swimtime="00:00:34.22" />
                    <SPLIT distance="75" swimtime="00:00:56.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="456" reactiontime="+72" swimtime="00:00:27.63" resultid="2751" lane="2" heatid="7349" entrytime="00:00:27.58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" status="DNS" swimtime="00:00:00.00" resultid="2749" lane="8" heatid="7077" entrytime="00:02:55.55" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-09-23" firstname="Agnieszka" gender="F" lastname="Bystrzycka" nation="POL" athleteid="2752">
              <RESULTS>
                <RESULT eventid="1092" points="635" reactiontime="+80" swimtime="00:01:08.40" resultid="2753" lane="4" heatid="6729" entrytime="00:01:11.91">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.17" />
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="75" swimtime="00:00:51.51" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1222" points="734" reactiontime="+77" swimtime="00:00:33.60" resultid="2754" lane="4" heatid="6853" entrytime="00:00:34.65">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.62" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1409" points="678" reactiontime="+82" swimtime="00:02:39.59" resultid="2755" lane="4" heatid="7001" entrytime="00:02:43.62">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.44" />
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                    <SPLIT distance="75" swimtime="00:00:55.55" />
                    <SPLIT distance="100" swimtime="00:01:15.82" />
                    <SPLIT distance="125" swimtime="00:01:36.12" />
                    <SPLIT distance="150" swimtime="00:01:56.97" />
                    <SPLIT distance="175" swimtime="00:02:18.02" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1679" points="690" reactiontime="+76" swimtime="00:01:13.63" resultid="2756" lane="4" heatid="7300" entrytime="00:01:15.15">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.89" />
                    <SPLIT distance="50" swimtime="00:00:34.75" />
                    <SPLIT distance="75" swimtime="00:00:53.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" status="DNS" swimtime="00:00:00.00" resultid="2757" lane="3" heatid="7335" entrytime="00:00:28.66" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-04-27" firstname="Hanna" gender="F" lastname="Sikacz" nation="POL" athleteid="2758">
              <RESULTS>
                <RESULT eventid="1581" points="289" reactiontime="+76" swimtime="00:03:14.16" resultid="2763" lane="8" heatid="7070" entrytime="00:03:12.59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.25" />
                    <SPLIT distance="50" swimtime="00:00:45.13" />
                    <SPLIT distance="75" swimtime="00:01:11.04" />
                    <SPLIT distance="100" swimtime="00:01:35.08" />
                    <SPLIT distance="125" swimtime="00:02:02.41" />
                    <SPLIT distance="150" swimtime="00:02:29.82" />
                    <SPLIT distance="175" swimtime="00:02:53.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1781" points="284" reactiontime="+70" swimtime="00:06:49.92" resultid="2765" lane="6" heatid="7356" entrytime="00:06:56.77">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.01" />
                    <SPLIT distance="50" swimtime="00:00:45.10" />
                    <SPLIT distance="75" swimtime="00:01:11.85" />
                    <SPLIT distance="100" swimtime="00:01:39.68" />
                    <SPLIT distance="125" swimtime="00:02:07.31" />
                    <SPLIT distance="150" swimtime="00:02:33.55" />
                    <SPLIT distance="175" swimtime="00:02:59.15" />
                    <SPLIT distance="200" swimtime="00:03:25.97" />
                    <SPLIT distance="225" swimtime="00:03:53.95" />
                    <SPLIT distance="250" swimtime="00:04:22.68" />
                    <SPLIT distance="275" swimtime="00:04:51.63" />
                    <SPLIT distance="300" swimtime="00:05:20.31" />
                    <SPLIT distance="325" swimtime="00:05:43.28" />
                    <SPLIT distance="350" swimtime="00:06:06.10" />
                    <SPLIT distance="375" swimtime="00:06:29.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1058" points="317" swimtime="00:12:03.97" resultid="2759" lane="1" heatid="6715" entrytime="00:11:56.77" />
                <RESULT eventid="1358" points="322" reactiontime="+78" swimtime="00:05:52.33" resultid="2761" lane="2" heatid="6897" entrytime="00:05:46.05">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.68" />
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                    <SPLIT distance="75" swimtime="00:00:58.13" />
                    <SPLIT distance="100" swimtime="00:01:19.27" />
                    <SPLIT distance="125" swimtime="00:01:41.77" />
                    <SPLIT distance="150" swimtime="00:02:04.27" />
                    <SPLIT distance="175" swimtime="00:02:27.37" />
                    <SPLIT distance="200" swimtime="00:02:50.63" />
                    <SPLIT distance="225" swimtime="00:03:13.73" />
                    <SPLIT distance="250" swimtime="00:03:37.38" />
                    <SPLIT distance="275" swimtime="00:03:59.47" />
                    <SPLIT distance="300" swimtime="00:04:22.22" />
                    <SPLIT distance="325" swimtime="00:04:44.23" />
                    <SPLIT distance="350" swimtime="00:05:07.06" />
                    <SPLIT distance="375" swimtime="00:05:30.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" status="DNS" swimtime="00:00:00.00" resultid="2764" lane="5" heatid="7332" entrytime="00:00:35.41" />
                <RESULT eventid="1547" status="DNS" swimtime="00:00:00.00" resultid="2762" lane="4" heatid="7051" entrytime="00:02:48.20" />
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="2760" lane="8" heatid="6826" entrytime="00:01:17.72" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-05-10" firstname="Maciej" gender="M" lastname="Koszarek" nation="POL" athleteid="2766">
              <RESULTS>
                <RESULT eventid="1564" points="360" reactiontime="+93" swimtime="00:02:24.69" resultid="2771" lane="2" heatid="7061" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.20" />
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                    <SPLIT distance="75" swimtime="00:00:50.95" />
                    <SPLIT distance="100" swimtime="00:01:10.03" />
                    <SPLIT distance="125" swimtime="00:01:28.73" />
                    <SPLIT distance="150" swimtime="00:01:48.04" />
                    <SPLIT distance="175" swimtime="00:02:06.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="246" reactiontime="+92" swimtime="00:02:58.79" resultid="2768" lane="7" heatid="6873" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.84" />
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                    <SPLIT distance="75" swimtime="00:00:57.91" />
                    <SPLIT distance="100" swimtime="00:01:19.90" />
                    <SPLIT distance="125" swimtime="00:01:42.96" />
                    <SPLIT distance="150" swimtime="00:02:07.82" />
                    <SPLIT distance="175" swimtime="00:02:33.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="309" reactiontime="+89" swimtime="00:01:14.49" resultid="2770" lane="4" heatid="7019" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.43" />
                    <SPLIT distance="50" swimtime="00:00:34.00" />
                    <SPLIT distance="75" swimtime="00:00:53.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="393" reactiontime="+83" swimtime="00:00:29.05" resultid="2772" lane="3" heatid="7344" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.18" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="przekroczenie limitu 11:30:00" eventid="1075" status="DSQ" swimtime="00:11:36.60" resultid="2767" lane="8" heatid="6721" entrytime="00:11:30.00" />
                <RESULT eventid="1798" status="DNS" swimtime="00:00:00.00" resultid="2773" lane="8" heatid="7362" entrytime="00:06:30.00" />
                <RESULT eventid="1375" status="DNS" swimtime="00:00:00.00" resultid="2769" heatid="6907" entrytime="00:05:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Dariusz" gender="M" lastname="Patrzałek" nation="POL" athleteid="2774">
              <RESULTS>
                <RESULT eventid="1496" points="121" reactiontime="+74" swimtime="00:00:49.43" resultid="2776" lane="3" heatid="7033" entrytime="00:00:54.54">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="136" reactiontime="+85" swimtime="00:00:44.63" resultid="2777" lane="8" heatid="7282" entrytime="00:00:46.58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="151" reactiontime="+100" swimtime="00:01:50.40" resultid="2778" lane="3" heatid="7303" entrytime="00:01:50.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.38" />
                    <SPLIT distance="50" swimtime="00:00:51.55" />
                    <SPLIT distance="75" swimtime="00:01:20.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="104" reactiontime="+88" swimtime="00:01:48.75" resultid="2775" heatid="6731" entrytime="00:01:52.52">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.54" />
                    <SPLIT distance="50" swimtime="00:00:50.32" />
                    <SPLIT distance="75" swimtime="00:01:22.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-09-09" firstname="Marlena" gender="F" lastname="Jakubów" nation="POL" athleteid="2779">
              <RESULTS>
                <RESULT eventid="1547" points="219" reactiontime="+106" swimtime="00:03:10.45" resultid="2784" lane="4" heatid="7050" entrytime="00:03:09.83">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.97" />
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                    <SPLIT distance="75" swimtime="00:01:04.31" />
                    <SPLIT distance="100" swimtime="00:01:29.19" />
                    <SPLIT distance="125" swimtime="00:01:54.89" />
                    <SPLIT distance="150" swimtime="00:02:21.62" />
                    <SPLIT distance="175" swimtime="00:02:47.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="221" reactiontime="+108" swimtime="00:00:50.10" resultid="2782" lane="3" heatid="6851" entrytime="00:00:44.44">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="273" reactiontime="+100" swimtime="00:01:21.43" resultid="2781" lane="3" heatid="6824" entrytime="00:01:25.44">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.69" />
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                    <SPLIT distance="75" swimtime="00:01:00.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="226" reactiontime="+108" swimtime="00:01:36.46" resultid="2780" lane="1" heatid="6725" entrytime="00:01:42.42">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.84" />
                    <SPLIT distance="50" swimtime="00:00:46.76" />
                    <SPLIT distance="75" swimtime="00:01:15.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="313" reactiontime="+96" swimtime="00:00:35.28" resultid="2786" lane="2" heatid="7332" entrytime="00:00:35.72">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="207" reactiontime="+125" swimtime="00:01:49.89" resultid="2785" heatid="7298" entrytime="00:01:49.87">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.59" />
                    <SPLIT distance="50" swimtime="00:00:51.92" />
                    <SPLIT distance="75" swimtime="00:01:20.58" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K 8" eventid="1409" reactiontime="+105" status="DSQ" swimtime="00:00:00.00" resultid="2783" lane="1" heatid="6999" entrytime="00:03:56.56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.44" />
                    <SPLIT distance="50" swimtime="00:00:52.74" />
                    <SPLIT distance="75" swimtime="00:01:22.19" />
                    <SPLIT distance="100" swimtime="00:01:52.71" />
                    <SPLIT distance="125" swimtime="00:02:23.21" />
                    <SPLIT distance="150" swimtime="00:02:53.83" />
                    <SPLIT distance="175" swimtime="00:03:24.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1177" points="486" reactiontime="+71" swimtime="00:01:50.31" resultid="2791" lane="3" heatid="6808" entrytime="00:02:02.02">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.61" />
                    <SPLIT distance="50" swimtime="00:00:28.22" />
                    <SPLIT distance="75" swimtime="00:00:42.02" />
                    <SPLIT distance="100" swimtime="00:00:56.80" />
                    <SPLIT distance="125" swimtime="00:01:09.15" />
                    <SPLIT distance="150" swimtime="00:01:22.98" />
                    <SPLIT distance="175" swimtime="00:01:35.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2766" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="2738" number="2" reactiontime="+54" />
                    <RELAYPOSITION athleteid="2705" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="2744" number="4" reactiontime="+18" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1341" points="482" reactiontime="+64" swimtime="00:02:01.77" resultid="2793" lane="7" heatid="6988" entrytime="00:02:02.02">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.32" />
                    <SPLIT distance="50" swimtime="00:00:30.67" />
                    <SPLIT distance="75" swimtime="00:00:45.23" />
                    <SPLIT distance="100" swimtime="00:01:03.11" />
                    <SPLIT distance="125" swimtime="00:01:17.45" />
                    <SPLIT distance="150" swimtime="00:01:34.19" />
                    <SPLIT distance="175" swimtime="00:01:47.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2705" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="2738" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="2766" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="2744" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1160" points="437" reactiontime="+81" swimtime="00:02:09.37" resultid="2790" lane="3" heatid="6813" entrytime="00:02:08.56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.67" />
                    <SPLIT distance="50" swimtime="00:00:28.02" />
                    <SPLIT distance="75" swimtime="00:00:44.72" />
                    <SPLIT distance="100" swimtime="00:01:02.38" />
                    <SPLIT distance="125" swimtime="00:01:17.12" />
                    <SPLIT distance="150" swimtime="00:01:33.07" />
                    <SPLIT distance="175" swimtime="00:01:49.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2752" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="2758" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="2722" number="3" reactiontime="+62" />
                    <RELAYPOSITION athleteid="2730" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="F" number="4">
              <RESULTS>
                <RESULT eventid="1324" points="408" reactiontime="+74" swimtime="00:02:26.00" resultid="2792" lane="5" heatid="6979" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.64" />
                    <SPLIT distance="50" swimtime="00:00:43.43" />
                    <SPLIT distance="75" swimtime="00:00:58.90" />
                    <SPLIT distance="100" swimtime="00:01:17.03" />
                    <SPLIT distance="125" swimtime="00:01:32.64" />
                    <SPLIT distance="150" swimtime="00:01:51.11" />
                    <SPLIT distance="175" swimtime="00:02:08.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2758" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="2752" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="2722" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="2779" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="X" number="5">
              <RESULTS>
                <RESULT eventid="1615" reactiontime="+79" swimtime="00:01:55.51" resultid="2789" lane="6" heatid="7443" entrytime="00:01:56.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.75" />
                    <SPLIT distance="50" swimtime="00:00:28.26" />
                    <SPLIT distance="75" swimtime="00:00:42.19" />
                    <SPLIT distance="100" swimtime="00:00:57.34" />
                    <SPLIT distance="125" swimtime="00:01:11.93" />
                    <SPLIT distance="150" swimtime="00:01:28.03" />
                    <SPLIT distance="175" swimtime="00:01:40.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2752" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="2766" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="2722" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="2744" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="7">
              <RESULTS>
                <RESULT eventid="1815" status="DNS" swimtime="00:00:00.00" resultid="2788" lane="7" heatid="7504" entrytime="00:02:16.77">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2705" number="1" />
                    <RELAYPOSITION athleteid="2752" number="2" />
                    <RELAYPOSITION athleteid="2712" number="3" />
                    <RELAYPOSITION athleteid="2758" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="8">
              <RESULTS>
                <RESULT eventid="1615" reactiontime="+82" swimtime="00:02:14.32" resultid="2787" lane="6" heatid="7442" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.63" />
                    <SPLIT distance="50" swimtime="00:00:28.08" />
                    <SPLIT distance="75" swimtime="00:00:44.56" />
                    <SPLIT distance="100" swimtime="00:01:03.87" />
                    <SPLIT distance="125" swimtime="00:01:21.02" />
                    <SPLIT distance="150" swimtime="00:01:40.26" />
                    <SPLIT distance="175" swimtime="00:01:56.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2705" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="2712" number="2" reactiontime="+45" />
                    <RELAYPOSITION athleteid="2779" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="2758" number="4" reactiontime="+17" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" number="9">
              <RESULTS>
                <RESULT eventid="1815" status="DNS" swimtime="00:00:00.00" resultid="2794" heatid="7504" entrytime="00:02:17.99">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2766" number="1" />
                    <RELAYPOSITION athleteid="2744" number="2" />
                    <RELAYPOSITION athleteid="2722" number="3" />
                    <RELAYPOSITION athleteid="2779" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="STWRO" name="Steef Wrocław" nation="POL" region="DOL">
          <CONTACT city="Wrocław" email="ste1@wp.pl" fax="(71)3377810" name="Stefan Skrzypek" phone="500 388 374" street="Piaskowa 17" zip="50-158" />
          <ATHLETES>
            <ATHLETE birthdate="1956-09-02" firstname="Stefan" gender="M" lastname="Skrzypek" nation="POL" athleteid="2807">
              <RESULTS>
                <RESULT eventid="1143" points="243" swimtime="00:23:21.16" resultid="2808" heatid="6750" entrytime="00:24:30.00" />
                <RESULT eventid="1273" points="177" reactiontime="+99" swimtime="00:03:19.31" resultid="2809" lane="6" heatid="6871" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.01" />
                    <SPLIT distance="50" swimtime="00:00:44.72" />
                    <SPLIT distance="75" swimtime="00:01:10.07" />
                    <SPLIT distance="100" swimtime="00:01:35.65" />
                    <SPLIT distance="125" swimtime="00:02:02.55" />
                    <SPLIT distance="150" swimtime="00:02:29.16" />
                    <SPLIT distance="175" swimtime="00:02:54.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="201" reactiontime="+100" swimtime="00:06:55.93" resultid="2814" lane="5" heatid="7360" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.14" />
                    <SPLIT distance="50" swimtime="00:00:43.32" />
                    <SPLIT distance="75" swimtime="00:01:07.74" />
                    <SPLIT distance="100" swimtime="00:01:33.55" />
                    <SPLIT distance="125" swimtime="00:02:03.21" />
                    <SPLIT distance="150" swimtime="00:02:31.57" />
                    <SPLIT distance="175" swimtime="00:02:59.96" />
                    <SPLIT distance="200" swimtime="00:03:28.49" />
                    <SPLIT distance="225" swimtime="00:03:58.19" />
                    <SPLIT distance="250" swimtime="00:04:27.91" />
                    <SPLIT distance="275" swimtime="00:04:57.63" />
                    <SPLIT distance="300" swimtime="00:05:27.40" />
                    <SPLIT distance="325" swimtime="00:05:50.42" />
                    <SPLIT distance="350" swimtime="00:06:13.78" />
                    <SPLIT distance="375" swimtime="00:06:35.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="259" reactiontime="+96" swimtime="00:05:44.87" resultid="2810" lane="5" heatid="6903" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.07" />
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                    <SPLIT distance="75" swimtime="00:00:58.69" />
                    <SPLIT distance="100" swimtime="00:01:20.34" />
                    <SPLIT distance="125" swimtime="00:01:41.06" />
                    <SPLIT distance="150" swimtime="00:02:03.00" />
                    <SPLIT distance="175" swimtime="00:02:24.50" />
                    <SPLIT distance="200" swimtime="00:02:47.02" />
                    <SPLIT distance="225" swimtime="00:03:09.00" />
                    <SPLIT distance="250" swimtime="00:03:31.17" />
                    <SPLIT distance="275" swimtime="00:03:53.34" />
                    <SPLIT distance="300" swimtime="00:04:16.08" />
                    <SPLIT distance="325" swimtime="00:04:37.99" />
                    <SPLIT distance="350" swimtime="00:05:00.84" />
                    <SPLIT distance="375" swimtime="00:05:22.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="211" reactiontime="+94" swimtime="00:03:11.69" resultid="2812" lane="5" heatid="7075" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.34" />
                    <SPLIT distance="50" swimtime="00:00:40.08" />
                    <SPLIT distance="75" swimtime="00:01:06.06" />
                    <SPLIT distance="100" swimtime="00:01:31.80" />
                    <SPLIT distance="125" swimtime="00:02:00.33" />
                    <SPLIT distance="150" swimtime="00:02:28.46" />
                    <SPLIT distance="175" swimtime="00:02:50.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="198" reactiontime="+97" swimtime="00:01:26.42" resultid="2811" heatid="7018" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.53" />
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                    <SPLIT distance="75" swimtime="00:01:02.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="2813" lane="4" heatid="7284" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WEZAB" name="Weteran  Zabrze" nation="POL">
          <CONTACT city="ZABRZE" name="BOSOWSKI  WŁODZIMIERZ" street="ŚW.JANA  4A/4" zip="41803" />
          <ATHLETES>
            <ATHLETE birthdate="1950-01-01" firstname="Barbara" gender="F" lastname="Brendler" nation="POL" athleteid="2816">
              <RESULTS>
                <RESULT eventid="1641" points="80" reactiontime="+99" swimtime="00:00:58.88" resultid="2821" heatid="7276" entrytime="00:00:53.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="195" reactiontime="+87" swimtime="00:00:41.27" resultid="2822" lane="7" heatid="7330" entrytime="00:00:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="165" reactiontime="+96" swimtime="00:01:36.36" resultid="2818" lane="5" heatid="6823" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.06" />
                    <SPLIT distance="50" swimtime="00:00:45.32" />
                    <SPLIT distance="75" swimtime="00:01:10.41" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K 8" eventid="1092" reactiontime="+90" status="DSQ" swimtime="00:00:00.00" resultid="2817" lane="5" heatid="6724" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.00" />
                    <SPLIT distance="50" swimtime="00:00:58.99" />
                    <SPLIT distance="75" swimtime="00:01:35.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" status="DNS" swimtime="00:00:00.00" resultid="2820" lane="5" heatid="7049" entrytime="00:03:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-01-01" firstname="Alfred" gender="M" lastname="Zabrzański" nation="POL" athleteid="2823">
              <RESULTS>
                <RESULT eventid="1205" points="338" reactiontime="+78" swimtime="00:01:07.51" resultid="2825" lane="2" heatid="6837" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.98" />
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                    <SPLIT distance="75" swimtime="00:00:49.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="226" swimtime="00:23:54.06" resultid="2824" lane="2" heatid="6750" entrytime="00:23:45.00" />
                <RESULT eventid="1764" points="340" reactiontime="+84" swimtime="00:00:30.46" resultid="2829" lane="4" heatid="7343" entrytime="00:00:30.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="256" reactiontime="+85" swimtime="00:05:46.34" resultid="2826" lane="1" heatid="6903" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.51" />
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                    <SPLIT distance="75" swimtime="00:00:57.19" />
                    <SPLIT distance="100" swimtime="00:01:18.25" />
                    <SPLIT distance="125" swimtime="00:01:40.25" />
                    <SPLIT distance="150" swimtime="00:02:02.25" />
                    <SPLIT distance="175" swimtime="00:02:24.89" />
                    <SPLIT distance="200" swimtime="00:02:47.11" />
                    <SPLIT distance="225" swimtime="00:03:09.49" />
                    <SPLIT distance="250" swimtime="00:03:31.70" />
                    <SPLIT distance="275" swimtime="00:03:54.61" />
                    <SPLIT distance="300" swimtime="00:04:17.43" />
                    <SPLIT distance="325" swimtime="00:04:39.64" />
                    <SPLIT distance="350" swimtime="00:05:02.50" />
                    <SPLIT distance="375" swimtime="00:05:25.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="270" reactiontime="+84" swimtime="00:02:39.20" resultid="2828" lane="6" heatid="7059" entrytime="00:02:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.27" />
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                    <SPLIT distance="75" swimtime="00:00:54.58" />
                    <SPLIT distance="100" swimtime="00:01:14.93" />
                    <SPLIT distance="125" swimtime="00:01:36.02" />
                    <SPLIT distance="150" swimtime="00:01:57.28" />
                    <SPLIT distance="175" swimtime="00:02:18.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="243" reactiontime="+73" swimtime="00:00:39.20" resultid="2827" lane="8" heatid="7037" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-01-01" firstname="Bernard" gender="M" lastname="Poloczek" nation="POL" athleteid="2830">
              <RESULTS>
                <RESULT eventid="1307" points="134" swimtime="00:03:42.37" resultid="2831" heatid="6883" entrytime="00:03:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.35" />
                    <SPLIT distance="50" swimtime="00:00:49.60" />
                    <SPLIT distance="75" swimtime="00:01:16.07" />
                    <SPLIT distance="100" swimtime="00:01:45.21" />
                    <SPLIT distance="125" swimtime="00:02:14.78" />
                    <SPLIT distance="150" swimtime="00:02:43.97" />
                    <SPLIT distance="175" swimtime="00:03:14.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="190" reactiontime="+64" swimtime="00:00:42.55" resultid="2832" lane="2" heatid="7036" entrytime="00:00:41.58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="166" reactiontime="+64" swimtime="00:01:35.41" resultid="2833" lane="2" heatid="7321" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.74" />
                    <SPLIT distance="50" swimtime="00:00:44.63" />
                    <SPLIT distance="75" swimtime="00:01:09.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-01" firstname="Beata" gender="F" lastname="Sulewska" nation="POL" athleteid="2834">
              <RESULTS>
                <RESULT eventid="1409" points="481" reactiontime="+85" swimtime="00:02:58.84" resultid="2838" lane="6" heatid="7001" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.73" />
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                    <SPLIT distance="75" swimtime="00:01:02.91" />
                    <SPLIT distance="100" swimtime="00:01:25.68" />
                    <SPLIT distance="125" swimtime="00:01:49.11" />
                    <SPLIT distance="150" swimtime="00:02:12.58" />
                    <SPLIT distance="175" swimtime="00:02:35.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="447" reactiontime="+87" swimtime="00:01:16.90" resultid="2835" lane="6" heatid="6729" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.28" />
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                    <SPLIT distance="75" swimtime="00:00:58.65" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1358" points="513" reactiontime="+83" swimtime="00:05:01.58" resultid="2837" lane="6" heatid="6898" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.38" />
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                    <SPLIT distance="75" swimtime="00:00:53.11" />
                    <SPLIT distance="100" swimtime="00:01:12.14" />
                    <SPLIT distance="125" swimtime="00:01:30.98" />
                    <SPLIT distance="150" swimtime="00:01:50.18" />
                    <SPLIT distance="175" swimtime="00:02:09.14" />
                    <SPLIT distance="200" swimtime="00:02:28.46" />
                    <SPLIT distance="225" swimtime="00:02:47.76" />
                    <SPLIT distance="250" swimtime="00:03:07.02" />
                    <SPLIT distance="275" swimtime="00:03:26.33" />
                    <SPLIT distance="300" swimtime="00:03:45.83" />
                    <SPLIT distance="325" swimtime="00:04:04.95" />
                    <SPLIT distance="350" swimtime="00:04:24.32" />
                    <SPLIT distance="375" swimtime="00:04:43.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="502" reactiontime="+87" swimtime="00:02:24.46" resultid="2839" lane="5" heatid="7053" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.15" />
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                    <SPLIT distance="75" swimtime="00:00:51.08" />
                    <SPLIT distance="100" swimtime="00:01:09.24" />
                    <SPLIT distance="125" swimtime="00:01:27.90" />
                    <SPLIT distance="150" swimtime="00:01:47.08" />
                    <SPLIT distance="175" swimtime="00:02:06.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="476" reactiontime="+83" swimtime="00:01:07.68" resultid="2836" lane="1" heatid="6828" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.83" />
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                    <SPLIT distance="75" swimtime="00:00:50.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="470" reactiontime="+87" swimtime="00:01:23.66" resultid="2840" lane="3" heatid="7300" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.91" />
                    <SPLIT distance="50" swimtime="00:00:39.95" />
                    <SPLIT distance="75" swimtime="00:01:01.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-01-01" firstname="Daniel" gender="M" lastname="Fecica" nation="POL" athleteid="2841">
              <RESULTS>
                <RESULT eventid="1239" points="244" reactiontime="+89" swimtime="00:00:43.47" resultid="2842" lane="1" heatid="6857" entrytime="00:00:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="221" reactiontime="+93" swimtime="00:03:30.65" resultid="2843" lane="4" heatid="7006" entrytime="00:03:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.54" />
                    <SPLIT distance="50" swimtime="00:00:46.70" />
                    <SPLIT distance="75" swimtime="00:01:12.91" />
                    <SPLIT distance="100" swimtime="00:01:39.70" />
                    <SPLIT distance="125" swimtime="00:02:07.19" />
                    <SPLIT distance="150" swimtime="00:02:34.78" />
                    <SPLIT distance="175" swimtime="00:03:02.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="226" reactiontime="+93" swimtime="00:01:36.71" resultid="2844" lane="4" heatid="7305" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.03" />
                    <SPLIT distance="50" swimtime="00:00:45.19" />
                    <SPLIT distance="75" swimtime="00:01:10.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-01-01" firstname="Krystyna" gender="F" lastname="Fecica" nation="POL" athleteid="2845">
              <RESULTS>
                <RESULT eventid="1445" points="124" swimtime="00:01:53.26" resultid="2849" lane="8" heatid="7013" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.83" />
                    <SPLIT distance="50" swimtime="00:00:54.27" />
                    <SPLIT distance="75" swimtime="00:01:24.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="118" swimtime="00:00:51.81" resultid="2850" lane="6" heatid="7276" entrytime="00:00:51.00" />
                <RESULT comment="Rekord Polski " eventid="1126" points="123" swimtime="00:31:31.00" resultid="2846" lane="5" heatid="6746" entrytime="00:33:00.00" />
                <RESULT eventid="1256" points="133" swimtime="00:04:02.81" resultid="2847" lane="4" heatid="6867" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.53" />
                    <SPLIT distance="50" swimtime="00:00:56.24" />
                    <SPLIT distance="75" swimtime="00:01:27.16" />
                    <SPLIT distance="100" swimtime="00:01:58.45" />
                    <SPLIT distance="125" swimtime="00:02:30.02" />
                    <SPLIT distance="150" swimtime="00:03:01.30" />
                    <SPLIT distance="175" swimtime="00:03:33.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1409" points="194" swimtime="00:04:02.11" resultid="2848" heatid="6999" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.70" />
                    <SPLIT distance="50" swimtime="00:00:58.06" />
                    <SPLIT distance="75" swimtime="00:01:28.19" />
                    <SPLIT distance="100" swimtime="00:01:59.22" />
                    <SPLIT distance="125" swimtime="00:02:29.84" />
                    <SPLIT distance="150" swimtime="00:03:01.19" />
                    <SPLIT distance="175" swimtime="00:03:32.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="190" swimtime="00:01:53.09" resultid="2851" lane="8" heatid="7297" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.37" />
                    <SPLIT distance="50" swimtime="00:00:55.69" />
                    <SPLIT distance="75" swimtime="00:01:24.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Grażyna" gender="F" lastname="Kiszczak" nation="POL" athleteid="2852">
              <RESULTS>
                <RESULT comment="Rekord Polski " eventid="1290" points="282" reactiontime="+76" swimtime="00:03:10.98" resultid="2854" lane="2" heatid="6878" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.82" />
                    <SPLIT distance="50" swimtime="00:00:45.25" />
                    <SPLIT distance="75" swimtime="00:01:09.15" />
                    <SPLIT distance="100" swimtime="00:01:33.93" />
                    <SPLIT distance="125" swimtime="00:01:58.51" />
                    <SPLIT distance="150" swimtime="00:02:22.98" />
                    <SPLIT distance="175" swimtime="00:02:48.03" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1479" points="344" reactiontime="+75" swimtime="00:00:39.47" resultid="2855" lane="8" heatid="7029" entrytime="00:00:40.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="311" reactiontime="+71" swimtime="00:01:26.73" resultid="2857" heatid="7316" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.64" />
                    <SPLIT distance="50" swimtime="00:00:42.65" />
                    <SPLIT distance="75" swimtime="00:01:04.97" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1092" points="292" reactiontime="+78" swimtime="00:01:28.56" resultid="2853" lane="4" heatid="6726" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.23" />
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                    <SPLIT distance="75" swimtime="00:01:06.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1581" status="DNS" swimtime="00:00:00.00" resultid="2856" lane="1" heatid="7069" entrytime="00:03:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="Stanisław" gender="M" lastname="Kiszczak" nation="POL" athleteid="2858">
              <RESULTS>
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="2860" heatid="7341" entrytime="00:00:32.50" />
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="2859" lane="7" heatid="6733" entrytime="00:01:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-01-01" firstname="Maria" gender="F" lastname="Buczkowska" nation="POL" athleteid="2861">
              <RESULTS>
                <RESULT eventid="1222" points="247" reactiontime="+111" swimtime="00:00:48.29" resultid="2862" lane="8" heatid="6850" entrytime="00:00:52.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="225" reactiontime="+114" swimtime="00:01:46.92" resultid="2864" lane="2" heatid="7297" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.40" />
                    <SPLIT distance="50" swimtime="00:00:52.75" />
                    <SPLIT distance="75" swimtime="00:01:20.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="144" reactiontime="+72" swimtime="00:00:52.74" resultid="2863" lane="3" heatid="7026" entrytime="00:00:54.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1942-01-01" firstname="Władysław" gender="M" lastname="Buczkowski" nation="POL" athleteid="2865">
              <RESULTS>
                <RESULT eventid="1564" points="196" reactiontime="+100" swimtime="00:02:57.19" resultid="2870" lane="7" heatid="7057" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.06" />
                    <SPLIT distance="50" swimtime="00:00:40.96" />
                    <SPLIT distance="75" swimtime="00:01:03.27" />
                    <SPLIT distance="100" swimtime="00:01:25.92" />
                    <SPLIT distance="125" swimtime="00:01:49.20" />
                    <SPLIT distance="150" swimtime="00:02:12.68" />
                    <SPLIT distance="175" swimtime="00:02:36.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="188" reactiontime="+73" swimtime="00:00:42.69" resultid="2869" heatid="7036" entrytime="00:00:44.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="255" reactiontime="+98" swimtime="00:01:32.81" resultid="2871" lane="2" heatid="7306" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.47" />
                    <SPLIT distance="50" swimtime="00:00:42.19" />
                    <SPLIT distance="75" swimtime="00:01:06.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="326" reactiontime="+93" swimtime="00:00:39.47" resultid="2868" lane="7" heatid="6859" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="266" reactiontime="+83" swimtime="00:00:33.06" resultid="2872" lane="8" heatid="7340" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="261" reactiontime="+95" swimtime="00:01:13.62" resultid="2867" lane="3" heatid="6834" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.69" />
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="75" swimtime="00:00:53.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="2866" lane="1" heatid="6735" entrytime="00:01:26.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1943-01-01" firstname="Renata" gender="F" lastname="Bastek" nation="POL" athleteid="2873">
              <RESULTS>
                <RESULT eventid="1092" points="236" reactiontime="+87" swimtime="00:01:35.09" resultid="2874" lane="7" heatid="6726" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.27" />
                    <SPLIT distance="50" swimtime="00:00:43.62" />
                    <SPLIT distance="75" swimtime="00:01:13.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="280" reactiontime="+84" swimtime="00:01:20.76" resultid="2875" lane="6" heatid="6825" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.81" />
                    <SPLIT distance="50" swimtime="00:00:38.09" />
                    <SPLIT distance="75" swimtime="00:00:59.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="270" reactiontime="+72" swimtime="00:00:42.77" resultid="2876" heatid="7028" entrytime="00:00:44.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="318" reactiontime="+85" swimtime="00:00:35.10" resultid="2878" lane="8" heatid="7332" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" status="DNS" swimtime="00:00:00.00" resultid="2877" lane="6" heatid="7277" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-01-01" firstname="Janina" gender="F" lastname="Bosowska" nation="POL" athleteid="2879">
              <RESULTS>
                <RESULT eventid="1679" points="198" reactiontime="+84" swimtime="00:01:51.50" resultid="2881" lane="4" heatid="7296" entrytime="00:01:58.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.94" />
                    <SPLIT distance="50" swimtime="00:00:52.01" />
                    <SPLIT distance="75" swimtime="00:01:20.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="237" reactiontime="+96" swimtime="00:00:48.97" resultid="2880" lane="6" heatid="6849" entrytime="00:00:53.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="175" reactiontime="+85" swimtime="00:00:42.78" resultid="2882" lane="4" heatid="7329" entrytime="00:00:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="Włodzimierz" gender="M" lastname="Bosowski" nation="POL" athleteid="2883">
              <RESULTS>
                <RESULT eventid="1764" points="188" reactiontime="+83" swimtime="00:00:37.09" resultid="2886" lane="4" heatid="7338" entrytime="00:00:35.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="167" reactiontime="+101" swimtime="00:00:41.65" resultid="2885" lane="3" heatid="7283" entrytime="00:00:38.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="100" reactiontime="+100" swimtime="00:00:52.60" resultid="2884" lane="8" heatid="7034" entrytime="00:00:53.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-01" firstname="Wiesław" gender="M" lastname="Kornicki" nation="POL" athleteid="2887">
              <RESULTS>
                <RESULT eventid="1764" points="320" reactiontime="+82" swimtime="00:00:31.09" resultid="2892" lane="4" heatid="7342" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="292" reactiontime="+87" swimtime="00:00:34.59" resultid="2891" lane="1" heatid="7286" entrytime="00:00:34.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="189" reactiontime="+75" swimtime="00:01:29.05" resultid="2888" lane="1" heatid="6734" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.92" />
                    <SPLIT distance="50" swimtime="00:00:41.02" />
                    <SPLIT distance="75" swimtime="00:01:08.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="264" reactiontime="+77" swimtime="00:01:13.33" resultid="2889" lane="6" heatid="6836" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.84" />
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                    <SPLIT distance="75" swimtime="00:00:53.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" status="DNS" swimtime="00:00:00.00" resultid="2890" lane="2" heatid="7035" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1615" reactiontime="+82" swimtime="00:02:14.52" resultid="2900" lane="4" heatid="7441" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.94" />
                    <SPLIT distance="50" swimtime="00:00:35.21" />
                    <SPLIT distance="75" swimtime="00:00:50.62" />
                    <SPLIT distance="100" swimtime="00:01:07.60" />
                    <SPLIT distance="125" swimtime="00:01:24.95" />
                    <SPLIT distance="150" swimtime="00:01:43.63" />
                    <SPLIT distance="175" swimtime="00:01:58.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2873" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="2865" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="2852" number="3" reactiontime="+54" />
                    <RELAYPOSITION athleteid="2823" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="PWWRO" name="Wrocławski Park Wodny S.A." nation="POL" region="DOL">
          <CONTACT city="Wrocław" name="Kujat Szymon" street="Borowska 99" zip="50-558" />
          <ATHLETES>
            <ATHLETE birthdate="1984-11-17" firstname="Michał" gender="M" lastname="Stasiaczek" nation="POL" athleteid="2902">
              <RESULTS>
                <RESULT eventid="1239" points="719" reactiontime="+69" swimtime="00:00:30.33" resultid="2904" lane="4" heatid="6866" entrytime="00:00:30.09">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="630" reactiontime="+68" swimtime="00:02:28.70" resultid="2905" lane="3" heatid="7011" entrytime="00:02:26.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.84" />
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                    <SPLIT distance="75" swimtime="00:00:51.45" />
                    <SPLIT distance="100" swimtime="00:01:11.15" />
                    <SPLIT distance="125" swimtime="00:01:30.51" />
                    <SPLIT distance="150" swimtime="00:01:49.79" />
                    <SPLIT distance="175" swimtime="00:02:09.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="720" reactiontime="+69" swimtime="00:01:05.70" resultid="2907" lane="4" heatid="7311" entrytime="00:01:06.99">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.14" />
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                    <SPLIT distance="75" swimtime="00:00:47.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="589" reactiontime="+74" swimtime="00:02:16.20" resultid="2906" lane="4" heatid="7080" entrytime="00:02:19.99">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.27" />
                    <SPLIT distance="50" swimtime="00:00:29.65" />
                    <SPLIT distance="75" swimtime="00:00:48.07" />
                    <SPLIT distance="100" swimtime="00:01:06.10" />
                    <SPLIT distance="125" swimtime="00:01:25.30" />
                    <SPLIT distance="150" swimtime="00:01:44.92" />
                    <SPLIT distance="175" swimtime="00:02:01.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="600" swimtime="00:01:00.64" resultid="2903" lane="5" heatid="6745" entrytime="00:01:00.50" />
                <RESULT eventid="1764" points="641" reactiontime="+69" swimtime="00:00:24.68" resultid="2908" lane="6" heatid="7354" entrytime="00:00:24.49">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-10-01" firstname="Tomasz" gender="M" lastname="Cimicki" nation="POL" athleteid="2909">
              <RESULTS>
                <RESULT eventid="1696" points="541" reactiontime="+82" swimtime="00:01:12.29" resultid="2913" lane="6" heatid="7311" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.83" />
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                    <SPLIT distance="75" swimtime="00:00:52.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="466" reactiontime="+84" swimtime="00:02:44.46" resultid="2912" lane="2" heatid="7011" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.38" />
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                    <SPLIT distance="75" swimtime="00:00:55.08" />
                    <SPLIT distance="100" swimtime="00:01:15.52" />
                    <SPLIT distance="125" swimtime="00:01:36.40" />
                    <SPLIT distance="150" swimtime="00:01:58.22" />
                    <SPLIT distance="175" swimtime="00:02:20.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="354" reactiontime="+93" swimtime="00:05:44.64" resultid="2914" heatid="7362" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.84" />
                    <SPLIT distance="50" swimtime="00:00:34.83" />
                    <SPLIT distance="75" swimtime="00:00:54.80" />
                    <SPLIT distance="100" swimtime="00:01:15.33" />
                    <SPLIT distance="125" swimtime="00:01:39.06" />
                    <SPLIT distance="150" swimtime="00:02:01.62" />
                    <SPLIT distance="175" swimtime="00:02:24.28" />
                    <SPLIT distance="200" swimtime="00:02:47.01" />
                    <SPLIT distance="225" swimtime="00:03:09.26" />
                    <SPLIT distance="250" swimtime="00:03:32.68" />
                    <SPLIT distance="275" swimtime="00:03:56.03" />
                    <SPLIT distance="300" swimtime="00:04:20.11" />
                    <SPLIT distance="325" swimtime="00:04:43.14" />
                    <SPLIT distance="350" swimtime="00:05:05.26" />
                    <SPLIT distance="375" swimtime="00:05:25.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="565" reactiontime="+82" swimtime="00:00:32.87" resultid="2911" lane="7" heatid="6866" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="416" reactiontime="+84" swimtime="00:01:08.49" resultid="2910" lane="8" heatid="6744" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.29" />
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                    <SPLIT distance="75" swimtime="00:00:51.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-04-08" firstname="Joanna" gender="F" lastname="Barabasz" nation="POL" athleteid="2915">
              <RESULTS>
                <RESULT comment="Rekord Polski " eventid="1290" points="490" reactiontime="+67" swimtime="00:02:38.81" resultid="2917" lane="6" heatid="6879" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.12" />
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                    <SPLIT distance="75" swimtime="00:00:57.03" />
                    <SPLIT distance="100" swimtime="00:01:17.54" />
                    <SPLIT distance="125" swimtime="00:01:38.34" />
                    <SPLIT distance="150" swimtime="00:01:59.24" />
                    <SPLIT distance="175" swimtime="00:02:20.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="513" reactiontime="+65" swimtime="00:01:13.37" resultid="2919" lane="2" heatid="7317" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.38" />
                    <SPLIT distance="50" swimtime="00:00:35.53" />
                    <SPLIT distance="75" swimtime="00:00:54.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="539" reactiontime="+65" swimtime="00:00:33.98" resultid="2918" lane="1" heatid="7031" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="487" reactiontime="+71" swimtime="00:01:14.73" resultid="2916" lane="5" heatid="6728" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.80" />
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                    <SPLIT distance="75" swimtime="00:00:56.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-07-28" firstname="Sylwia" gender="F" lastname="Madej" nation="POL" athleteid="2920">
              <RESULTS>
                <RESULT eventid="1547" points="465" reactiontime="+80" swimtime="00:02:28.14" resultid="2923" lane="4" heatid="7052" entrytime="00:02:35.33">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.93" />
                    <SPLIT distance="50" swimtime="00:00:33.59" />
                    <SPLIT distance="75" swimtime="00:00:51.90" />
                    <SPLIT distance="100" swimtime="00:01:10.90" />
                    <SPLIT distance="125" swimtime="00:01:30.04" />
                    <SPLIT distance="150" swimtime="00:01:49.78" />
                    <SPLIT distance="175" swimtime="00:02:09.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="501" reactiontime="+74" swimtime="00:01:06.56" resultid="2922" lane="6" heatid="6828" entrytime="00:01:06.83">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.21" />
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                    <SPLIT distance="75" swimtime="00:00:49.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="489" reactiontime="+85" swimtime="00:00:30.41" resultid="2925" lane="4" heatid="7334" entrytime="00:00:30.67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="417" reactiontime="+74" swimtime="00:01:18.68" resultid="2921" lane="3" heatid="6728" entrytime="00:01:20.11">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.73" />
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                    <SPLIT distance="75" swimtime="00:01:00.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" status="DNS" swimtime="00:00:00.00" resultid="2924" lane="5" heatid="7279" entrytime="00:00:34.71" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-04-20" firstname="Robert" gender="M" lastname="Kazimirów" nation="POL" athleteid="2926">
              <RESULTS>
                <RESULT eventid="1462" points="467" reactiontime="+86" swimtime="00:01:04.95" resultid="2928" lane="1" heatid="7022" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.83" />
                    <SPLIT distance="50" swimtime="00:00:30.04" />
                    <SPLIT distance="75" swimtime="00:00:47.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="505" reactiontime="+82" swimtime="00:00:59.05" resultid="2927" lane="4" heatid="6845" entrytime="00:00:57.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.63" />
                    <SPLIT distance="50" swimtime="00:00:28.56" />
                    <SPLIT distance="75" swimtime="00:00:43.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="522" reactiontime="+85" swimtime="00:00:26.42" resultid="2930" lane="4" heatid="7352" entrytime="00:00:26.25">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="501" reactiontime="+87" swimtime="00:00:28.89" resultid="2929" lane="5" heatid="7292" entrytime="00:00:28.48">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-09" firstname="Michał" gender="M" lastname="Witkowski" nation="POL" athleteid="2931">
              <RESULTS>
                <RESULT eventid="1496" points="563" reactiontime="+76" swimtime="00:00:29.62" resultid="2934" lane="5" heatid="7043" entrytime="00:00:27.81">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="623" reactiontime="+77" swimtime="00:00:55.08" resultid="2933" lane="4" heatid="6846" entrytime="00:00:52.93">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.43" />
                    <SPLIT distance="50" swimtime="00:00:26.20" />
                    <SPLIT distance="75" swimtime="00:00:40.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="667" reactiontime="+75" swimtime="00:00:24.35" resultid="2937" lane="4" heatid="7354" entrytime="00:00:23.27">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="542" swimtime="00:01:02.73" resultid="2932" lane="3" heatid="6745" entrytime="00:00:59.91" />
                <RESULT eventid="1564" points="509" reactiontime="+79" swimtime="00:02:08.95" resultid="2935" lane="3" heatid="7066" entrytime="00:01:55.54">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.82" />
                    <SPLIT distance="50" swimtime="00:00:27.35" />
                    <SPLIT distance="75" swimtime="00:00:42.67" />
                    <SPLIT distance="100" swimtime="00:00:58.50" />
                    <SPLIT distance="125" swimtime="00:01:15.11" />
                    <SPLIT distance="150" swimtime="00:01:32.65" />
                    <SPLIT distance="175" swimtime="00:01:50.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="538" reactiontime="+74" swimtime="00:00:28.23" resultid="2936" lane="2" heatid="7294" entrytime="00:00:25.88">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-08-06" firstname="Jakub" gender="M" lastname="Balcerzak" nation="POL" athleteid="2938">
              <RESULTS>
                <RESULT eventid="1730" points="448" reactiontime="+61" swimtime="00:01:08.66" resultid="2943" lane="5" heatid="7325" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.47" />
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                    <SPLIT distance="75" swimtime="00:00:50.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="356" reactiontime="+60" swimtime="00:02:40.71" resultid="2940" lane="6" heatid="6885" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.92" />
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                    <SPLIT distance="75" swimtime="00:00:57.12" />
                    <SPLIT distance="100" swimtime="00:01:18.21" />
                    <SPLIT distance="125" swimtime="00:01:37.95" />
                    <SPLIT distance="150" swimtime="00:01:58.67" />
                    <SPLIT distance="175" swimtime="00:02:20.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="385" reactiontime="+74" swimtime="00:01:10.26" resultid="2939" heatid="6742" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.33" />
                    <SPLIT distance="50" swimtime="00:00:29.79" />
                    <SPLIT distance="75" swimtime="00:00:51.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="2942" lane="7" heatid="7292" entrytime="00:00:29.00" />
                <RESULT comment="04" eventid="1496" status="DSQ" swimtime="00:00:00.00" resultid="2941" lane="7" heatid="7042" entrytime="00:00:30.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-04-26" firstname="Łukasz" gender="M" lastname="Mazurkiewicz" nation="POL" athleteid="2944">
              <RESULTS>
                <RESULT eventid="1598" points="290" reactiontime="+95" swimtime="00:02:52.52" resultid="2946" lane="2" heatid="7078" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.56" />
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                    <SPLIT distance="75" swimtime="00:00:54.34" />
                    <SPLIT distance="100" swimtime="00:01:15.95" />
                    <SPLIT distance="125" swimtime="00:01:39.41" />
                    <SPLIT distance="150" swimtime="00:02:04.64" />
                    <SPLIT distance="175" swimtime="00:02:28.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="499" reactiontime="+79" swimtime="00:00:26.82" resultid="2948" lane="8" heatid="7349" entrytime="00:00:27.77">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="440" reactiontime="+78" swimtime="00:00:30.17" resultid="2947" heatid="7289" entrytime="00:00:31.52">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.83" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Z 2" eventid="1109" reactiontime="+87" status="DSQ" swimtime="00:01:13.31" resultid="2945" lane="6" heatid="6740" entrytime="00:01:12.99">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.75" />
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                    <SPLIT distance="75" swimtime="00:00:55.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-07-05" firstname="Sebastian" gender="M" lastname="Figarski" nation="POL" athleteid="2949">
              <RESULTS>
                <RESULT eventid="1496" points="575" reactiontime="+68" swimtime="00:00:29.42" resultid="2952" lane="7" heatid="7043" entrytime="00:00:29.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="588" reactiontime="+74" swimtime="00:02:15.97" resultid="2951" lane="3" heatid="6887" entrytime="00:02:19.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.23" />
                    <SPLIT distance="50" swimtime="00:00:31.07" />
                    <SPLIT distance="75" swimtime="00:00:47.47" />
                    <SPLIT distance="100" swimtime="00:01:04.50" />
                    <SPLIT distance="125" swimtime="00:01:21.77" />
                    <SPLIT distance="150" swimtime="00:01:39.51" />
                    <SPLIT distance="175" swimtime="00:01:57.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="598" reactiontime="+65" swimtime="00:01:02.33" resultid="2954" lane="2" heatid="7326" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.87" />
                    <SPLIT distance="50" swimtime="00:00:30.31" />
                    <SPLIT distance="75" swimtime="00:00:46.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="554" reactiontime="+87" swimtime="00:02:19.05" resultid="2953" lane="7" heatid="7080" entrytime="00:02:25.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.43" />
                    <SPLIT distance="50" swimtime="00:00:29.05" />
                    <SPLIT distance="75" swimtime="00:00:47.13" />
                    <SPLIT distance="100" swimtime="00:01:04.46" />
                    <SPLIT distance="125" swimtime="00:01:24.75" />
                    <SPLIT distance="150" swimtime="00:01:45.55" />
                    <SPLIT distance="175" swimtime="00:02:02.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="530" reactiontime="+79" swimtime="00:01:03.20" resultid="2950" lane="2" heatid="6744" entrytime="00:01:05.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.25" />
                    <SPLIT distance="50" swimtime="00:00:28.82" />
                    <SPLIT distance="75" swimtime="00:00:47.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1985-02-27" firstname="Patrycja" gender="F" lastname="Skibińska" nation="POL" athleteid="2955">
              <RESULTS>
                <RESULT eventid="1092" points="503" reactiontime="+82" swimtime="00:01:13.93" resultid="2956" lane="1" heatid="6728" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.21" />
                    <SPLIT distance="50" swimtime="00:00:34.49" />
                    <SPLIT distance="75" swimtime="00:00:55.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1445" points="452" reactiontime="+84" swimtime="00:01:13.76" resultid="2957" heatid="7014" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.76" />
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                    <SPLIT distance="75" swimtime="00:00:53.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="469" reactiontime="+83" swimtime="00:00:32.76" resultid="2958" lane="6" heatid="7279" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" status="DNS" swimtime="00:00:00.00" resultid="2959" lane="3" heatid="7333" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-29" firstname="Karolina" gender="F" lastname="Kubatek" nation="POL" athleteid="2960">
              <RESULTS>
                <RESULT eventid="1445" points="295" reactiontime="+87" swimtime="00:01:25.03" resultid="2962" lane="1" heatid="7012">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.91" />
                    <SPLIT distance="50" swimtime="00:00:38.01" />
                    <SPLIT distance="75" swimtime="00:01:00.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="382" swimtime="00:01:20.99" resultid="2961" lane="2" heatid="6723">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.99" />
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                    <SPLIT distance="75" swimtime="00:01:01.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="346" reactiontime="+90" swimtime="00:00:36.24" resultid="2963" lane="1" heatid="7275">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" status="DNS" swimtime="00:00:00.00" resultid="2964" lane="3" heatid="7327" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-07-21" firstname="Mateusz" gender="M" lastname="Dudek" nation="POL" athleteid="2965">
              <RESULTS>
                <RESULT eventid="1411" points="579" reactiontime="+77" swimtime="00:02:32.94" resultid="2967" lane="4" heatid="7011" entrytime="00:02:15.54">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.30" />
                    <SPLIT distance="50" swimtime="00:00:33.64" />
                    <SPLIT distance="75" swimtime="00:00:52.56" />
                    <SPLIT distance="100" swimtime="00:01:12.09" />
                    <SPLIT distance="125" swimtime="00:01:31.58" />
                    <SPLIT distance="150" swimtime="00:01:51.44" />
                    <SPLIT distance="175" swimtime="00:02:11.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="612" reactiontime="+72" swimtime="00:01:09.38" resultid="2968" lane="5" heatid="7311" entrytime="00:01:09.82">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.75" />
                    <SPLIT distance="50" swimtime="00:00:32.16" />
                    <SPLIT distance="75" swimtime="00:00:50.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="655" reactiontime="+74" swimtime="00:00:31.29" resultid="2966" lane="2" heatid="6866" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1177" points="662" reactiontime="+77" swimtime="00:01:39.54" resultid="2973" lane="4" heatid="6810" entrytime="00:01:39.99">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.66" />
                    <SPLIT distance="50" swimtime="00:00:49.66" />
                    <SPLIT distance="75" swimtime="00:01:01.97" />
                    <SPLIT distance="100" swimtime="00:01:15.38" />
                    <SPLIT distance="125" swimtime="00:01:27.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2949" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="2926" number="2" reactiontime="+64" />
                    <RELAYPOSITION athleteid="2902" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="2931" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1341" points="645" reactiontime="+65" swimtime="00:01:50.54" resultid="2974" lane="4" heatid="6988" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.67" />
                    <SPLIT distance="50" swimtime="00:00:29.47" />
                    <SPLIT distance="75" swimtime="00:00:42.95" />
                    <SPLIT distance="100" swimtime="00:00:59.13" />
                    <SPLIT distance="125" swimtime="00:01:10.84" />
                    <SPLIT distance="150" swimtime="00:01:25.33" />
                    <SPLIT distance="175" swimtime="00:01:37.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2949" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="2902" number="2" reactiontime="+42" />
                    <RELAYPOSITION athleteid="2931" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="2926" number="4" reactiontime="+9" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1324" points="498" reactiontime="+65" swimtime="00:02:16.58" resultid="2971" lane="4" heatid="6979" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.09" />
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                    <SPLIT distance="75" swimtime="00:00:51.91" />
                    <SPLIT distance="100" swimtime="00:01:12.35" />
                    <SPLIT distance="125" swimtime="00:01:28.06" />
                    <SPLIT distance="150" swimtime="00:01:47.12" />
                    <SPLIT distance="175" swimtime="00:02:01.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2915" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="2955" number="2" reactiontime="+72" />
                    <RELAYPOSITION athleteid="2960" number="3" reactiontime="+71" />
                    <RELAYPOSITION athleteid="2920" number="4" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1160" points="495" reactiontime="+81" swimtime="00:02:04.09" resultid="2972" lane="4" heatid="6813" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.19" />
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                    <SPLIT distance="75" swimtime="00:00:46.90" />
                    <SPLIT distance="100" swimtime="00:01:03.46" />
                    <SPLIT distance="125" swimtime="00:01:18.46" />
                    <SPLIT distance="150" swimtime="00:01:34.27" />
                    <SPLIT distance="175" swimtime="00:01:48.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2955" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="2960" number="2" reactiontime="+81" />
                    <RELAYPOSITION athleteid="2915" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="2920" number="4" reactiontime="+64" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1615" reactiontime="+84" swimtime="00:01:52.30" resultid="2975" lane="5" heatid="7443" entrytime="00:01:51.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.93" />
                    <SPLIT distance="50" swimtime="00:00:26.39" />
                    <SPLIT distance="75" swimtime="00:00:41.76" />
                    <SPLIT distance="100" swimtime="00:00:57.99" />
                    <SPLIT distance="125" swimtime="00:01:12.40" />
                    <SPLIT distance="150" swimtime="00:01:27.95" />
                    <SPLIT distance="175" swimtime="00:01:39.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2926" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="2915" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="2920" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="2931" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1815" reactiontime="+64" swimtime="00:02:02.82" resultid="2976" lane="4" heatid="7504" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.19" />
                    <SPLIT distance="50" swimtime="00:00:34.80" />
                    <SPLIT distance="75" swimtime="00:00:48.91" />
                    <SPLIT distance="100" swimtime="00:01:05.30" />
                    <SPLIT distance="125" swimtime="00:01:17.41" />
                    <SPLIT distance="150" swimtime="00:01:32.42" />
                    <SPLIT distance="175" swimtime="00:01:46.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2915" number="1" reactiontime="+64" />
                    <RELAYPOSITION athleteid="2902" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="2931" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="2920" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1815" reactiontime="+72" swimtime="00:02:06.29" resultid="2969" lane="5" heatid="7504" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.85" />
                    <SPLIT distance="50" swimtime="00:00:29.70" />
                    <SPLIT distance="75" swimtime="00:00:44.59" />
                    <SPLIT distance="100" swimtime="00:01:02.24" />
                    <SPLIT distance="125" swimtime="00:01:16.95" />
                    <SPLIT distance="150" swimtime="00:01:34.76" />
                    <SPLIT distance="175" swimtime="00:01:49.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2949" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="2909" number="2" reactiontime="+68" />
                    <RELAYPOSITION athleteid="2955" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="2960" number="4" reactiontime="+67" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1615" status="DNS" swimtime="00:00:00.00" resultid="2970" lane="1" heatid="7443" entrytime="00:01:58.00" />
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MASOP" name="Sopot Masters" nation="POL" region="POM">
          <CONTACT city="SOPOT" email="sopotmasters@o2.pl" internet="www.sopotmasters.pl" name="Gorbaczow Mirosław" phone="696 258 185" state="POMOR" street="ul. Haffnera 57" zip="81-715" />
          <ATHLETES>
            <ATHLETE birthdate="1964-08-04" firstname="Joanna" gender="F" lastname="Puchalska" nation="POL" athleteid="2989">
              <RESULTS>
                <RESULT comment="Rekord Polski " eventid="1581" points="481" reactiontime="+80" swimtime="00:02:43.90" resultid="2993" lane="2" heatid="7070" entrytime="00:02:52.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.88" />
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                    <SPLIT distance="75" swimtime="00:00:57.15" />
                    <SPLIT distance="100" swimtime="00:01:20.42" />
                    <SPLIT distance="125" swimtime="00:01:42.98" />
                    <SPLIT distance="150" swimtime="00:02:06.96" />
                    <SPLIT distance="175" swimtime="00:02:26.20" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1445" points="489" reactiontime="+79" swimtime="00:01:11.83" resultid="2992" lane="6" heatid="7014" entrytime="00:01:17.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.70" />
                    <SPLIT distance="50" swimtime="00:00:33.87" />
                    <SPLIT distance="75" swimtime="00:00:52.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="465" reactiontime="+69" swimtime="00:00:32.86" resultid="2994" lane="2" heatid="7279" entrytime="00:00:34.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.33" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1256" points="475" reactiontime="+85" swimtime="00:02:39.07" resultid="2990" lane="4" heatid="6868" entrytime="00:02:52.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.18" />
                    <SPLIT distance="50" swimtime="00:00:35.84" />
                    <SPLIT distance="75" swimtime="00:00:55.56" />
                    <SPLIT distance="100" swimtime="00:01:15.75" />
                    <SPLIT distance="125" swimtime="00:01:36.04" />
                    <SPLIT distance="150" swimtime="00:01:57.00" />
                    <SPLIT distance="175" swimtime="00:02:17.98" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1781" points="476" reactiontime="+81" swimtime="00:05:44.99" resultid="2995" lane="4" heatid="7356" entrytime="00:05:59.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.22" />
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                    <SPLIT distance="75" swimtime="00:00:57.11" />
                    <SPLIT distance="100" swimtime="00:01:17.68" />
                    <SPLIT distance="125" swimtime="00:01:41.92" />
                    <SPLIT distance="150" swimtime="00:02:04.46" />
                    <SPLIT distance="175" swimtime="00:02:27.32" />
                    <SPLIT distance="200" swimtime="00:02:49.80" />
                    <SPLIT distance="225" swimtime="00:03:14.27" />
                    <SPLIT distance="250" swimtime="00:03:38.63" />
                    <SPLIT distance="275" swimtime="00:04:02.75" />
                    <SPLIT distance="300" swimtime="00:04:27.26" />
                    <SPLIT distance="325" swimtime="00:04:47.50" />
                    <SPLIT distance="350" swimtime="00:05:07.19" />
                    <SPLIT distance="375" swimtime="00:05:26.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="480" reactiontime="+81" swimtime="00:05:08.29" resultid="2991" lane="5" heatid="6898" entrytime="00:05:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.62" />
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                    <SPLIT distance="75" swimtime="00:00:54.92" />
                    <SPLIT distance="100" swimtime="00:01:14.38" />
                    <SPLIT distance="125" swimtime="00:01:34.14" />
                    <SPLIT distance="150" swimtime="00:01:54.27" />
                    <SPLIT distance="175" swimtime="00:02:13.57" />
                    <SPLIT distance="200" swimtime="00:02:33.30" />
                    <SPLIT distance="225" swimtime="00:02:53.06" />
                    <SPLIT distance="250" swimtime="00:03:12.67" />
                    <SPLIT distance="275" swimtime="00:03:32.39" />
                    <SPLIT distance="300" swimtime="00:03:51.87" />
                    <SPLIT distance="325" swimtime="00:04:11.25" />
                    <SPLIT distance="350" swimtime="00:04:31.15" />
                    <SPLIT distance="375" swimtime="00:04:49.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-04-08" firstname="Jerzy" gender="M" lastname="Bendig" nation="POL" athleteid="2996">
              <RESULTS>
                <RESULT eventid="1564" points="236" reactiontime="+114" swimtime="00:02:46.54" resultid="3000" lane="7" heatid="7060" entrytime="00:02:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.68" />
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                    <SPLIT distance="75" swimtime="00:00:57.91" />
                    <SPLIT distance="100" swimtime="00:01:19.42" />
                    <SPLIT distance="125" swimtime="00:01:41.07" />
                    <SPLIT distance="150" swimtime="00:02:02.82" />
                    <SPLIT distance="175" swimtime="00:02:24.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="240" swimtime="00:23:26.66" resultid="2997" lane="4" heatid="6750" entrytime="00:23:17.00" entrycourse="SCM" />
                <RESULT eventid="1205" points="244" reactiontime="+98" swimtime="00:01:15.27" resultid="2998" heatid="6837" entrytime="00:01:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.88" />
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                    <SPLIT distance="75" swimtime="00:00:55.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="258" reactiontime="+109" swimtime="00:05:45.37" resultid="2999" lane="5" heatid="6905" entrytime="00:05:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.27" />
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                    <SPLIT distance="75" swimtime="00:00:59.74" />
                    <SPLIT distance="100" swimtime="00:01:21.00" />
                    <SPLIT distance="125" swimtime="00:01:42.52" />
                    <SPLIT distance="150" swimtime="00:02:05.14" />
                    <SPLIT distance="175" swimtime="00:02:27.18" />
                    <SPLIT distance="200" swimtime="00:02:49.57" />
                    <SPLIT distance="225" swimtime="00:03:11.50" />
                    <SPLIT distance="250" swimtime="00:03:34.20" />
                    <SPLIT distance="275" swimtime="00:03:56.07" />
                    <SPLIT distance="300" swimtime="00:04:18.27" />
                    <SPLIT distance="325" swimtime="00:04:40.36" />
                    <SPLIT distance="350" swimtime="00:05:02.71" />
                    <SPLIT distance="375" swimtime="00:05:23.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="210" reactiontime="+99" swimtime="00:00:38.62" resultid="3001" lane="7" heatid="7285" entrytime="00:00:36.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="210" reactiontime="+113" swimtime="00:06:50.01" resultid="3002" lane="2" heatid="7361" entrytime="00:06:40.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.46" />
                    <SPLIT distance="50" swimtime="00:00:46.61" />
                    <SPLIT distance="75" swimtime="00:01:13.88" />
                    <SPLIT distance="100" swimtime="00:01:42.76" />
                    <SPLIT distance="125" swimtime="00:02:10.62" />
                    <SPLIT distance="150" swimtime="00:02:37.81" />
                    <SPLIT distance="175" swimtime="00:03:04.57" />
                    <SPLIT distance="200" swimtime="00:03:30.75" />
                    <SPLIT distance="225" swimtime="00:03:59.32" />
                    <SPLIT distance="250" swimtime="00:04:27.78" />
                    <SPLIT distance="275" swimtime="00:04:56.00" />
                    <SPLIT distance="300" swimtime="00:05:24.17" />
                    <SPLIT distance="325" swimtime="00:05:47.12" />
                    <SPLIT distance="350" swimtime="00:06:08.68" />
                    <SPLIT distance="375" swimtime="00:06:30.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-10-13" firstname="Mirosław" gender="M" lastname="Gorbaczow" nation="POL" athleteid="3003">
              <RESULTS>
                <RESULT eventid="1496" points="153" reactiontime="+106" swimtime="00:00:45.67" resultid="3008" lane="4" heatid="7035" entrytime="00:00:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="114" reactiontime="+89" swimtime="00:01:48.21" resultid="3009" lane="5" heatid="7320" entrytime="00:01:45.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.61" />
                    <SPLIT distance="50" swimtime="00:00:50.78" />
                    <SPLIT distance="75" swimtime="00:01:19.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="118" reactiontime="+82" swimtime="00:03:51.91" resultid="3006" lane="6" heatid="6882" entrytime="00:03:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.70" />
                    <SPLIT distance="50" swimtime="00:00:50.09" />
                    <SPLIT distance="75" swimtime="00:01:18.17" />
                    <SPLIT distance="100" swimtime="00:01:48.81" />
                    <SPLIT distance="125" swimtime="00:02:21.24" />
                    <SPLIT distance="150" swimtime="00:02:53.89" />
                    <SPLIT distance="175" swimtime="00:03:24.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="169" reactiontime="+102" swimtime="00:03:50.48" resultid="3007" lane="7" heatid="7004" entrytime="00:03:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.19" />
                    <SPLIT distance="50" swimtime="00:00:53.85" />
                    <SPLIT distance="75" swimtime="00:01:23.27" />
                    <SPLIT distance="100" swimtime="00:01:53.26" />
                    <SPLIT distance="125" swimtime="00:02:24.42" />
                    <SPLIT distance="150" swimtime="00:02:55.99" />
                    <SPLIT distance="175" swimtime="00:03:24.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="94" reactiontime="+117" swimtime="00:08:55.87" resultid="3010" heatid="7358" entrytime="00:08:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.13" />
                    <SPLIT distance="50" swimtime="00:01:00.67" />
                    <SPLIT distance="75" swimtime="00:01:35.36" />
                    <SPLIT distance="100" swimtime="00:02:11.28" />
                    <SPLIT distance="125" swimtime="00:02:48.28" />
                    <SPLIT distance="150" swimtime="00:03:27.05" />
                    <SPLIT distance="175" swimtime="00:04:02.72" />
                    <SPLIT distance="200" swimtime="00:04:39.41" />
                    <SPLIT distance="225" swimtime="00:05:16.07" />
                    <SPLIT distance="250" swimtime="00:05:52.33" />
                    <SPLIT distance="275" swimtime="00:06:27.67" />
                    <SPLIT distance="300" swimtime="00:07:02.72" />
                    <SPLIT distance="325" swimtime="00:07:33.82" />
                    <SPLIT distance="350" swimtime="00:08:06.47" />
                    <SPLIT distance="375" swimtime="00:08:35.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="151" reactiontime="+103" swimtime="00:01:36.04" resultid="3004" lane="3" heatid="6732" entrytime="00:01:36.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.30" />
                    <SPLIT distance="50" swimtime="00:00:45.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="185" reactiontime="+101" swimtime="00:01:22.43" resultid="3005" lane="8" heatid="6833" entrytime="00:01:24.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.93" />
                    <SPLIT distance="50" swimtime="00:00:40.68" />
                    <SPLIT distance="75" swimtime="00:01:01.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-02-08" firstname="Anna" gender="F" lastname="Maciejowska" nation="POL" athleteid="3011">
              <RESULTS>
                <RESULT comment="Rekord Polski " eventid="1126" points="268" swimtime="00:24:21.06" resultid="3012" lane="6" heatid="6747" entrytime="00:24:30.00" entrycourse="SCM" />
                <RESULT eventid="1187" points="328" reactiontime="+84" swimtime="00:01:16.63" resultid="3013" lane="7" heatid="6826" entrytime="00:01:16.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.94" />
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                    <SPLIT distance="75" swimtime="00:00:57.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="353" reactiontime="+77" swimtime="00:00:39.13" resultid="3014" lane="4" heatid="7028" entrytime="00:00:41.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.23" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1547" points="316" reactiontime="+81" swimtime="00:02:48.52" resultid="3015" lane="2" heatid="7051" entrytime="00:02:54.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.10" />
                    <SPLIT distance="50" swimtime="00:00:37.59" />
                    <SPLIT distance="75" swimtime="00:00:59.01" />
                    <SPLIT distance="100" swimtime="00:01:21.59" />
                    <SPLIT distance="125" swimtime="00:01:43.75" />
                    <SPLIT distance="150" swimtime="00:02:06.02" />
                    <SPLIT distance="175" swimtime="00:02:28.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="292" reactiontime="+82" swimtime="00:00:38.36" resultid="3016" lane="5" heatid="7278" entrytime="00:00:39.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="370" reactiontime="+81" swimtime="00:00:33.37" resultid="3017" lane="8" heatid="7333" entrytime="00:00:34.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-04-20" firstname="Piotr" gender="M" lastname="Suwara" nation="POL" athleteid="3018">
              <RESULTS>
                <RESULT eventid="1375" points="417" reactiontime="+92" swimtime="00:04:54.41" resultid="3021" lane="4" heatid="6907" entrytime="00:05:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.79" />
                    <SPLIT distance="50" swimtime="00:00:32.42" />
                    <SPLIT distance="75" swimtime="00:00:50.06" />
                    <SPLIT distance="100" swimtime="00:01:08.38" />
                    <SPLIT distance="125" swimtime="00:01:27.09" />
                    <SPLIT distance="150" swimtime="00:01:46.05" />
                    <SPLIT distance="175" swimtime="00:02:05.10" />
                    <SPLIT distance="200" swimtime="00:02:24.49" />
                    <SPLIT distance="225" swimtime="00:02:43.60" />
                    <SPLIT distance="250" swimtime="00:03:02.86" />
                    <SPLIT distance="275" swimtime="00:03:22.28" />
                    <SPLIT distance="300" swimtime="00:03:41.58" />
                    <SPLIT distance="325" swimtime="00:04:00.50" />
                    <SPLIT distance="350" swimtime="00:04:19.40" />
                    <SPLIT distance="375" swimtime="00:04:37.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="405" swimtime="00:10:19.53" resultid="3019" lane="4" heatid="6721" entrytime="00:10:45.00" entrycourse="SCM" />
                <RESULT eventid="1564" points="438" reactiontime="+85" swimtime="00:02:15.56" resultid="3023" lane="7" heatid="7063" entrytime="00:02:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.16" />
                    <SPLIT distance="50" swimtime="00:00:30.05" />
                    <SPLIT distance="75" swimtime="00:00:46.79" />
                    <SPLIT distance="100" swimtime="00:01:04.13" />
                    <SPLIT distance="125" swimtime="00:01:21.82" />
                    <SPLIT distance="150" swimtime="00:01:40.11" />
                    <SPLIT distance="175" swimtime="00:01:58.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="504" reactiontime="+85" swimtime="00:00:59.09" resultid="3020" lane="2" heatid="6842" entrytime="00:01:01.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.41" />
                    <SPLIT distance="50" swimtime="00:00:28.26" />
                    <SPLIT distance="75" swimtime="00:00:43.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="436" reactiontime="+84" swimtime="00:00:30.27" resultid="3024" lane="5" heatid="7288" entrytime="00:00:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="474" reactiontime="+85" swimtime="00:00:27.29" resultid="3025" heatid="7347" entrytime="00:00:28.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" status="DNS" swimtime="00:00:00.00" resultid="3022" lane="4" heatid="7036" entrytime="00:00:40.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-06-03" firstname="Leszek" gender="M" lastname="Wilkowski" nation="POL" athleteid="3026">
              <RESULTS>
                <RESULT eventid="1143" points="260" swimtime="00:22:50.13" resultid="3027" lane="3" heatid="6751" entrytime="00:21:40.00" entrycourse="SCM" />
                <RESULT eventid="1307" points="240" reactiontime="+95" swimtime="00:03:03.13" resultid="3029" lane="6" heatid="6884" entrytime="00:03:01.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.14" />
                    <SPLIT distance="50" swimtime="00:00:41.29" />
                    <SPLIT distance="75" swimtime="00:01:03.48" />
                    <SPLIT distance="100" swimtime="00:01:26.53" />
                    <SPLIT distance="125" swimtime="00:01:49.66" />
                    <SPLIT distance="150" swimtime="00:02:14.52" />
                    <SPLIT distance="175" swimtime="00:02:39.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="268" reactiontime="+92" swimtime="00:06:17.92" resultid="3033" lane="1" heatid="7362" entrytime="00:06:28.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.24" />
                    <SPLIT distance="50" swimtime="00:00:41.25" />
                    <SPLIT distance="75" swimtime="00:01:05.34" />
                    <SPLIT distance="100" swimtime="00:01:31.62" />
                    <SPLIT distance="125" swimtime="00:01:57.36" />
                    <SPLIT distance="150" swimtime="00:02:20.78" />
                    <SPLIT distance="175" swimtime="00:02:43.84" />
                    <SPLIT distance="200" swimtime="00:03:07.50" />
                    <SPLIT distance="225" swimtime="00:03:33.98" />
                    <SPLIT distance="250" swimtime="00:04:01.23" />
                    <SPLIT distance="275" swimtime="00:04:27.88" />
                    <SPLIT distance="300" swimtime="00:04:55.58" />
                    <SPLIT distance="325" swimtime="00:05:17.51" />
                    <SPLIT distance="350" swimtime="00:05:38.79" />
                    <SPLIT distance="375" swimtime="00:05:59.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="400" reactiontime="+97" swimtime="00:00:28.87" resultid="3032" lane="8" heatid="7348" entrytime="00:00:28.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="253" reactiontime="+97" swimtime="00:03:21.44" resultid="3030" lane="4" heatid="7005" entrytime="00:03:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.51" />
                    <SPLIT distance="50" swimtime="00:00:41.73" />
                    <SPLIT distance="75" swimtime="00:01:06.34" />
                    <SPLIT distance="100" swimtime="00:01:32.69" />
                    <SPLIT distance="125" swimtime="00:01:59.28" />
                    <SPLIT distance="150" swimtime="00:02:26.93" />
                    <SPLIT distance="175" swimtime="00:02:54.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="374" reactiontime="+110" swimtime="00:01:05.30" resultid="3028" lane="3" heatid="6840" entrytime="00:01:05.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.31" />
                    <SPLIT distance="50" swimtime="00:00:30.04" />
                    <SPLIT distance="75" swimtime="00:00:47.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" status="DNS" swimtime="00:00:00.00" resultid="3031" lane="5" heatid="7077" entrytime="00:02:53.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-03-28" firstname="Krzysztof" gender="M" lastname="Tarasek" nation="POL" athleteid="3034">
              <RESULTS>
                <RESULT eventid="1375" points="398" reactiontime="+79" swimtime="00:04:59.15" resultid="3037" heatid="6906" entrytime="00:05:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.77" />
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                    <SPLIT distance="75" swimtime="00:00:52.27" />
                    <SPLIT distance="100" swimtime="00:01:11.07" />
                    <SPLIT distance="125" swimtime="00:01:29.67" />
                    <SPLIT distance="150" swimtime="00:01:48.67" />
                    <SPLIT distance="175" swimtime="00:02:07.78" />
                    <SPLIT distance="200" swimtime="00:02:26.84" />
                    <SPLIT distance="225" swimtime="00:02:45.95" />
                    <SPLIT distance="250" swimtime="00:03:05.49" />
                    <SPLIT distance="275" swimtime="00:03:24.92" />
                    <SPLIT distance="300" swimtime="00:03:44.17" />
                    <SPLIT distance="325" swimtime="00:04:03.41" />
                    <SPLIT distance="350" swimtime="00:04:22.72" />
                    <SPLIT distance="375" swimtime="00:04:41.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="426" reactiontime="+61" swimtime="00:00:32.51" resultid="3038" lane="7" heatid="7038" entrytime="00:00:36.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="407" reactiontime="+69" swimtime="00:01:10.85" resultid="3041" lane="2" heatid="7323" entrytime="00:01:18.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.79" />
                    <SPLIT distance="50" swimtime="00:00:34.41" />
                    <SPLIT distance="75" swimtime="00:00:52.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="387" reactiontime="+79" swimtime="00:00:31.50" resultid="3040" lane="8" heatid="7287" entrytime="00:00:34.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="364" reactiontime="+82" swimtime="00:01:11.63" resultid="3035" lane="8" heatid="6738" entrytime="00:01:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.46" />
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                    <SPLIT distance="75" swimtime="00:00:54.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="3039" lane="1" heatid="7062" entrytime="00:02:28.00" entrycourse="SCM" />
                <RESULT eventid="1307" status="DNS" swimtime="00:00:00.00" resultid="3036" lane="8" heatid="6885" entrytime="00:02:57.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1177" status="DNS" swimtime="00:00:00.00" resultid="3043" lane="1" heatid="6809" entrytime="00:01:56.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3026" number="1" />
                    <RELAYPOSITION athleteid="2996" number="2" />
                    <RELAYPOSITION athleteid="3034" number="3" />
                    <RELAYPOSITION athleteid="3018" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1341" status="DNS" swimtime="00:00:00.00" resultid="3042" lane="8" heatid="6987" entrytime="00:02:16.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3034" number="1" />
                    <RELAYPOSITION athleteid="3026" number="2" />
                    <RELAYPOSITION athleteid="2996" number="3" />
                    <RELAYPOSITION athleteid="3018" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1615" status="DNS" swimtime="00:00:00.00" resultid="3044" lane="7" heatid="7442" entrytime="00:02:16.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3011" number="1" />
                    <RELAYPOSITION athleteid="3003" number="2" />
                    <RELAYPOSITION athleteid="2989" number="3" />
                    <RELAYPOSITION athleteid="2996" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="1815" status="DNS" swimtime="00:00:00.00" resultid="3045" lane="8" heatid="7504" entrytime="00:02:19.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3034" number="1" />
                    <RELAYPOSITION athleteid="3011" number="2" />
                    <RELAYPOSITION athleteid="2989" number="3" />
                    <RELAYPOSITION athleteid="3018" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MABIA" name="Masters Białystok" nation="POL">
          <CONTACT email="wzmasters@wp.pl" name="Żmiejko" phone="797309140" />
          <ATHLETES>
            <ATHLETE birthdate="1979-01-01" firstname="Dominika" gender="F" lastname="Michalik" nation="POL" athleteid="3052">
              <RESULTS>
                <RESULT eventid="1187" points="472" reactiontime="+78" swimtime="00:01:07.90" resultid="3053" lane="7" heatid="6828" entrytime="00:01:08.09">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.05" />
                    <SPLIT distance="50" swimtime="00:00:33.16" />
                    <SPLIT distance="75" swimtime="00:00:50.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="419" reactiontime="+81" swimtime="00:05:22.60" resultid="3054" lane="3" heatid="6898" entrytime="00:05:17.63">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.99" />
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                    <SPLIT distance="75" swimtime="00:00:54.78" />
                    <SPLIT distance="100" swimtime="00:01:14.42" />
                    <SPLIT distance="125" swimtime="00:01:34.21" />
                    <SPLIT distance="150" swimtime="00:01:54.44" />
                    <SPLIT distance="175" swimtime="00:02:14.53" />
                    <SPLIT distance="200" swimtime="00:02:34.79" />
                    <SPLIT distance="225" swimtime="00:02:55.10" />
                    <SPLIT distance="250" swimtime="00:03:15.67" />
                    <SPLIT distance="275" swimtime="00:03:36.16" />
                    <SPLIT distance="300" swimtime="00:03:57.17" />
                    <SPLIT distance="325" swimtime="00:04:17.94" />
                    <SPLIT distance="350" swimtime="00:04:38.97" />
                    <SPLIT distance="375" swimtime="00:05:01.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="458" reactiontime="+83" swimtime="00:02:28.95" resultid="3055" lane="7" heatid="7053" entrytime="00:02:30.73">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.39" />
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                    <SPLIT distance="75" swimtime="00:00:52.25" />
                    <SPLIT distance="100" swimtime="00:01:10.61" />
                    <SPLIT distance="125" swimtime="00:01:29.79" />
                    <SPLIT distance="150" swimtime="00:01:49.32" />
                    <SPLIT distance="175" swimtime="00:02:09.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="364" reactiontime="+80" swimtime="00:00:35.65" resultid="3056" lane="1" heatid="7279" entrytime="00:00:35.21">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="338" reactiontime="+65" swimtime="00:01:24.29" resultid="3057" lane="6" heatid="7316" entrytime="00:01:26.88">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.55" />
                    <SPLIT distance="50" swimtime="00:00:42.17" />
                    <SPLIT distance="75" swimtime="00:01:03.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Mirosław" gender="M" lastname="Matusik" nation="POL" athleteid="3058">
              <RESULTS>
                <RESULT eventid="1411" points="336" reactiontime="+84" swimtime="00:03:03.41" resultid="3061" lane="4" heatid="7009" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.52" />
                    <SPLIT distance="50" swimtime="00:00:41.01" />
                    <SPLIT distance="75" swimtime="00:01:03.91" />
                    <SPLIT distance="100" swimtime="00:01:27.62" />
                    <SPLIT distance="125" swimtime="00:01:51.95" />
                    <SPLIT distance="150" swimtime="00:02:16.60" />
                    <SPLIT distance="175" swimtime="00:02:40.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="413" reactiontime="+93" swimtime="00:01:19.05" resultid="3063" lane="6" heatid="7309" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.84" />
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                    <SPLIT distance="75" swimtime="00:00:57.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="447" reactiontime="+84" swimtime="00:00:35.53" resultid="3060" lane="4" heatid="6863" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="279" reactiontime="+84" swimtime="00:01:18.26" resultid="3059" lane="1" heatid="6738" entrytime="00:01:17.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.27" />
                    <SPLIT distance="50" swimtime="00:00:36.88" />
                    <SPLIT distance="75" swimtime="00:00:59.31" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="04" eventid="1645" reactiontime="+48" status="DSQ" swimtime="00:00:00.00" resultid="3062" lane="5" heatid="7282" entrytime="00:00:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Joanna" gender="F" lastname="Wasilewicz" nation="POL" athleteid="3064">
              <RESULTS>
                <RESULT eventid="1547" points="205" reactiontime="+95" swimtime="00:03:14.58" resultid="3067" lane="5" heatid="7050" entrytime="00:03:12.32">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.82" />
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                    <SPLIT distance="75" swimtime="00:01:04.50" />
                    <SPLIT distance="100" swimtime="00:01:29.93" />
                    <SPLIT distance="125" swimtime="00:01:55.49" />
                    <SPLIT distance="150" swimtime="00:02:22.48" />
                    <SPLIT distance="175" swimtime="00:02:49.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="199" reactiontime="+90" swimtime="00:06:53.33" resultid="3066" lane="5" heatid="6895" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.17" />
                    <SPLIT distance="50" swimtime="00:00:43.77" />
                    <SPLIT distance="75" swimtime="00:01:08.67" />
                    <SPLIT distance="100" swimtime="00:01:34.07" />
                    <SPLIT distance="125" swimtime="00:01:59.97" />
                    <SPLIT distance="150" swimtime="00:02:26.94" />
                    <SPLIT distance="175" swimtime="00:02:53.94" />
                    <SPLIT distance="200" swimtime="00:03:20.05" />
                    <SPLIT distance="225" swimtime="00:03:47.70" />
                    <SPLIT distance="250" swimtime="00:04:14.11" />
                    <SPLIT distance="275" swimtime="00:04:41.50" />
                    <SPLIT distance="300" swimtime="00:05:07.88" />
                    <SPLIT distance="325" swimtime="00:05:36.09" />
                    <SPLIT distance="350" swimtime="00:06:02.32" />
                    <SPLIT distance="375" swimtime="00:06:29.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="247" reactiontime="+83" swimtime="00:01:24.22" resultid="3065" lane="7" heatid="6825" entrytime="00:01:22.77">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.15" />
                    <SPLIT distance="50" swimtime="00:00:39.36" />
                    <SPLIT distance="75" swimtime="00:01:02.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="276" reactiontime="+85" swimtime="00:00:36.78" resultid="3068" lane="6" heatid="7332" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-01" firstname="Maciej" gender="M" lastname="Daszuta" nation="POL" athleteid="3069">
              <RESULTS>
                <RESULT eventid="1496" points="468" reactiontime="+63" swimtime="00:00:31.51" resultid="3073" lane="4" heatid="7041" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="379" reactiontime="+65" swimtime="00:01:12.55" resultid="3075" lane="2" heatid="7324" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.51" />
                    <SPLIT distance="50" swimtime="00:00:34.71" />
                    <SPLIT distance="75" swimtime="00:00:53.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="487" reactiontime="+88" swimtime="00:00:29.18" resultid="3074" lane="1" heatid="7291" entrytime="00:00:29.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="530" reactiontime="+79" swimtime="00:00:33.57" resultid="3071" lane="6" heatid="6865" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="407" reactiontime="+93" swimtime="00:01:08.99" resultid="3070" lane="7" heatid="6742" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.59" />
                    <SPLIT distance="50" swimtime="00:00:31.26" />
                    <SPLIT distance="75" swimtime="00:00:51.88" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K 11" eventid="1411" reactiontime="+81" status="DSQ" swimtime="00:00:00.00" resultid="3072" lane="5" heatid="7008" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.91" />
                    <SPLIT distance="50" swimtime="00:00:40.20" />
                    <SPLIT distance="75" swimtime="00:01:03.49" />
                    <SPLIT distance="100" swimtime="00:01:27.09" />
                    <SPLIT distance="125" swimtime="00:01:51.64" />
                    <SPLIT distance="150" swimtime="00:02:15.39" />
                    <SPLIT distance="175" swimtime="00:02:38.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Elżbieta" gender="F" lastname="Piwowarczyk" nation="POL" athleteid="3076">
              <RESULTS>
                <RESULT eventid="1290" points="297" reactiontime="+66" swimtime="00:03:07.52" resultid="3079" lane="5" heatid="6878" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.82" />
                    <SPLIT distance="50" swimtime="00:00:43.13" />
                    <SPLIT distance="75" swimtime="00:01:06.42" />
                    <SPLIT distance="100" swimtime="00:01:30.54" />
                    <SPLIT distance="125" swimtime="00:01:54.70" />
                    <SPLIT distance="150" swimtime="00:02:19.53" />
                    <SPLIT distance="175" swimtime="00:02:44.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1581" points="309" reactiontime="+77" swimtime="00:03:09.95" resultid="3081" heatid="7070" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.88" />
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                    <SPLIT distance="75" swimtime="00:01:04.92" />
                    <SPLIT distance="100" swimtime="00:01:29.43" />
                    <SPLIT distance="125" swimtime="00:01:57.59" />
                    <SPLIT distance="150" swimtime="00:02:26.18" />
                    <SPLIT distance="175" swimtime="00:02:48.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="321" reactiontime="+67" swimtime="00:01:25.82" resultid="3083" lane="7" heatid="7316" entrytime="00:01:27.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.29" />
                    <SPLIT distance="50" swimtime="00:00:41.93" />
                    <SPLIT distance="75" swimtime="00:01:04.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="300" reactiontime="+75" swimtime="00:00:38.02" resultid="3082" lane="6" heatid="7278" entrytime="00:00:39.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="342" reactiontime="+69" swimtime="00:00:39.54" resultid="3080" lane="5" heatid="7029" entrytime="00:00:39.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="370" reactiontime="+77" swimtime="00:01:13.64" resultid="3078" lane="3" heatid="6826" entrytime="00:01:14.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.17" />
                    <SPLIT distance="50" swimtime="00:00:36.05" />
                    <SPLIT distance="75" swimtime="00:00:55.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="329" reactiontime="+73" swimtime="00:01:25.09" resultid="3077" lane="1" heatid="6727" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.76" />
                    <SPLIT distance="50" swimtime="00:00:38.86" />
                    <SPLIT distance="75" swimtime="00:01:04.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-01" firstname="Wojciech" gender="M" lastname="Żmiejko" nation="POL" athleteid="3084">
              <RESULTS>
                <RESULT eventid="1462" points="408" reactiontime="+77" swimtime="00:01:07.95" resultid="3087" lane="8" heatid="7022" entrytime="00:01:07.95">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.77" />
                    <SPLIT distance="50" swimtime="00:00:31.55" />
                    <SPLIT distance="75" swimtime="00:00:49.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="404" reactiontime="+82" swimtime="00:02:34.41" resultid="3088" lane="7" heatid="7079" entrytime="00:02:33.95">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.74" />
                    <SPLIT distance="50" swimtime="00:00:32.38" />
                    <SPLIT distance="75" swimtime="00:00:52.25" />
                    <SPLIT distance="100" swimtime="00:01:11.70" />
                    <SPLIT distance="125" swimtime="00:01:34.25" />
                    <SPLIT distance="150" swimtime="00:01:57.74" />
                    <SPLIT distance="175" swimtime="00:02:16.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="456" reactiontime="+77" swimtime="00:00:29.82" resultid="3089" lane="6" heatid="7290" entrytime="00:00:30.25">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="418" reactiontime="+79" swimtime="00:01:08.36" resultid="3085" lane="5" heatid="6742" entrytime="00:01:09.35">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.82" />
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                    <SPLIT distance="75" swimtime="00:00:51.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="476" reactiontime="+79" swimtime="00:00:27.25" resultid="3090" lane="7" heatid="7349" entrytime="00:00:27.75">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="477" reactiontime="+78" swimtime="00:01:00.21" resultid="3086" lane="8" heatid="6843" entrytime="00:01:00.95">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.10" />
                    <SPLIT distance="50" swimtime="00:00:29.22" />
                    <SPLIT distance="75" swimtime="00:00:44.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ASBYD" name="Astoria Bydgoszcz" nation="POL">
          <CONTACT email="sikoreczka7@o2.pl" name="Sikorska Małgorzata" />
          <ATHLETES>
            <ATHLETE birthdate="1957-01-01" firstname="Krzysztof" gender="M" lastname="Kawecki" nation="POL" athleteid="3094">
              <RESULTS>
                <RESULT eventid="1598" points="290" reactiontime="+84" swimtime="00:02:52.44" resultid="3099" lane="3" heatid="7077" entrytime="00:02:52.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.82" />
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                    <SPLIT distance="75" swimtime="00:01:00.81" />
                    <SPLIT distance="100" swimtime="00:01:23.35" />
                    <SPLIT distance="125" swimtime="00:01:47.99" />
                    <SPLIT distance="150" swimtime="00:02:12.54" />
                    <SPLIT distance="175" swimtime="00:02:33.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="281" reactiontime="+67" swimtime="00:02:53.81" resultid="3097" lane="5" heatid="6885" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.85" />
                    <SPLIT distance="50" swimtime="00:00:40.77" />
                    <SPLIT distance="75" swimtime="00:01:02.69" />
                    <SPLIT distance="100" swimtime="00:01:24.65" />
                    <SPLIT distance="125" swimtime="00:01:46.99" />
                    <SPLIT distance="150" swimtime="00:02:09.61" />
                    <SPLIT distance="175" swimtime="00:02:32.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="307" reactiontime="+82" swimtime="00:03:08.94" resultid="3098" lane="6" heatid="7009" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.78" />
                    <SPLIT distance="50" swimtime="00:00:42.89" />
                    <SPLIT distance="75" swimtime="00:01:06.61" />
                    <SPLIT distance="100" swimtime="00:01:30.31" />
                    <SPLIT distance="125" swimtime="00:01:55.09" />
                    <SPLIT distance="150" swimtime="00:02:19.96" />
                    <SPLIT distance="175" swimtime="00:02:45.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="276" reactiontime="+83" swimtime="00:06:14.32" resultid="3101" lane="1" heatid="7363" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.18" />
                    <SPLIT distance="50" swimtime="00:00:40.94" />
                    <SPLIT distance="75" swimtime="00:01:05.37" />
                    <SPLIT distance="100" swimtime="00:01:30.83" />
                    <SPLIT distance="125" swimtime="00:01:55.10" />
                    <SPLIT distance="150" swimtime="00:02:18.40" />
                    <SPLIT distance="175" swimtime="00:02:42.10" />
                    <SPLIT distance="200" swimtime="00:03:05.71" />
                    <SPLIT distance="225" swimtime="00:03:32.21" />
                    <SPLIT distance="250" swimtime="00:03:58.61" />
                    <SPLIT distance="275" swimtime="00:04:25.01" />
                    <SPLIT distance="300" swimtime="00:04:50.84" />
                    <SPLIT distance="325" swimtime="00:05:12.24" />
                    <SPLIT distance="350" swimtime="00:05:33.19" />
                    <SPLIT distance="375" swimtime="00:05:53.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="248" swimtime="00:23:11.34" resultid="3095" lane="5" heatid="6750" entrytime="00:23:30.00" />
                <RESULT eventid="1730" points="238" reactiontime="+68" swimtime="00:01:24.70" resultid="3100" lane="6" heatid="7323" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.37" />
                    <SPLIT distance="50" swimtime="00:00:41.63" />
                    <SPLIT distance="75" swimtime="00:01:03.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="349" reactiontime="+85" swimtime="00:00:38.57" resultid="3096" lane="5" heatid="6861" entrytime="00:00:37.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1928-01-01" firstname="Wacława" gender="F" lastname="Wilczynska" nation="POL" athleteid="3102">
              <RESULTS>
                <RESULT comment="Rekord Polski " eventid="1409" points="20" reactiontime="+107" swimtime="00:08:31.54" resultid="3105" lane="4" heatid="6997" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:53.30" />
                    <SPLIT distance="50" swimtime="00:01:56.22" />
                    <SPLIT distance="75" swimtime="00:03:00.34" />
                    <SPLIT distance="100" swimtime="00:04:05.33" />
                    <SPLIT distance="125" swimtime="00:05:11.99" />
                    <SPLIT distance="150" swimtime="00:06:19.35" />
                    <SPLIT distance="175" swimtime="00:07:26.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="40" reactiontime="+85" swimtime="00:02:33.93" resultid="3103" lane="1" heatid="6822" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:33.78" />
                    <SPLIT distance="50" swimtime="00:01:13.19" />
                    <SPLIT distance="75" swimtime="00:01:55.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="33" reactiontime="+74" swimtime="00:06:27.70" resultid="3104" lane="3" heatid="6875" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:43.59" />
                    <SPLIT distance="50" swimtime="00:01:32.45" />
                    <SPLIT distance="75" swimtime="00:02:20.71" />
                    <SPLIT distance="100" swimtime="00:03:09.51" />
                    <SPLIT distance="125" swimtime="00:03:57.95" />
                    <SPLIT distance="150" swimtime="00:04:47.89" />
                    <SPLIT distance="175" swimtime="00:05:39.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" status="DNS" swimtime="00:00:00.00" resultid="3108" lane="5" heatid="7328" entrytime="00:01:00.00" />
                <RESULT eventid="1679" status="DNS" swimtime="00:00:00.00" resultid="3107" lane="4" heatid="7295" entrytime="00:03:31.00" />
                <RESULT eventid="1547" status="DNS" swimtime="00:00:00.00" resultid="3106" lane="4" heatid="7048" entrytime="00:05:18.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="BALEG" name="Barakuda Legnica" nation="POL" region="DOL">
          <CONTACT email="jmalchar@o2.pl" name="MALCHAR JOWITA" phone="506034671" />
          <ATHLETES>
            <ATHLETE birthdate="1971-01-01" firstname="Sebastian" gender="M" lastname="Hudyka" nation="POL" athleteid="3110">
              <RESULTS>
                <RESULT eventid="1075" points="250" swimtime="00:12:07.94" resultid="3111" lane="2" heatid="6719" entrytime="00:12:20.00" />
                <RESULT eventid="1375" points="256" reactiontime="+91" swimtime="00:05:46.26" resultid="3113" lane="4" heatid="6903" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.46" />
                    <SPLIT distance="50" swimtime="00:00:37.43" />
                    <SPLIT distance="75" swimtime="00:00:58.33" />
                    <SPLIT distance="100" swimtime="00:01:19.34" />
                    <SPLIT distance="125" swimtime="00:01:40.89" />
                    <SPLIT distance="150" swimtime="00:02:03.11" />
                    <SPLIT distance="175" swimtime="00:02:25.68" />
                    <SPLIT distance="200" swimtime="00:02:47.91" />
                    <SPLIT distance="225" swimtime="00:03:10.25" />
                    <SPLIT distance="250" swimtime="00:03:32.64" />
                    <SPLIT distance="275" swimtime="00:03:55.20" />
                    <SPLIT distance="300" swimtime="00:04:17.76" />
                    <SPLIT distance="325" swimtime="00:04:40.62" />
                    <SPLIT distance="350" swimtime="00:05:03.62" />
                    <SPLIT distance="375" swimtime="00:05:25.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="275" reactiontime="+102" swimtime="00:01:12.35" resultid="3112" lane="1" heatid="6835" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.29" />
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                    <SPLIT distance="75" swimtime="00:00:53.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="270" reactiontime="+102" swimtime="00:00:32.90" resultid="3115" lane="3" heatid="7340" entrytime="00:00:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="3114" lane="5" heatid="7057" entrytime="00:02:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-12-28" firstname="Jowita" gender="F" lastname="Malchar" nation="POL" athleteid="3116">
              <RESULTS>
                <RESULT eventid="1126" points="338" swimtime="00:22:32.84" resultid="3117" lane="2" heatid="6747" entrytime="00:23:00.00" />
                <RESULT eventid="1358" points="346" reactiontime="+77" swimtime="00:05:44.00" resultid="3119" lane="6" heatid="6897" entrytime="00:05:48.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.92" />
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                    <SPLIT distance="75" swimtime="00:00:58.46" />
                    <SPLIT distance="100" swimtime="00:01:19.62" />
                    <SPLIT distance="125" swimtime="00:01:41.34" />
                    <SPLIT distance="150" swimtime="00:02:03.25" />
                    <SPLIT distance="175" swimtime="00:02:25.28" />
                    <SPLIT distance="200" swimtime="00:02:47.26" />
                    <SPLIT distance="225" swimtime="00:03:09.15" />
                    <SPLIT distance="250" swimtime="00:03:31.08" />
                    <SPLIT distance="275" swimtime="00:03:53.79" />
                    <SPLIT distance="300" swimtime="00:04:15.83" />
                    <SPLIT distance="325" swimtime="00:04:38.22" />
                    <SPLIT distance="350" swimtime="00:05:00.78" />
                    <SPLIT distance="375" swimtime="00:05:22.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="355" reactiontime="+82" swimtime="00:02:42.01" resultid="3121" lane="8" heatid="7052" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.23" />
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                    <SPLIT distance="75" swimtime="00:00:56.64" />
                    <SPLIT distance="100" swimtime="00:01:17.30" />
                    <SPLIT distance="125" swimtime="00:01:38.74" />
                    <SPLIT distance="150" swimtime="00:02:00.35" />
                    <SPLIT distance="175" swimtime="00:02:22.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="394" reactiontime="+82" swimtime="00:01:12.08" resultid="3118" lane="2" heatid="6827" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.46" />
                    <SPLIT distance="50" swimtime="00:00:34.14" />
                    <SPLIT distance="75" swimtime="00:00:52.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="352" reactiontime="+69" swimtime="00:00:39.18" resultid="3120" lane="2" heatid="7029" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="353" reactiontime="+79" swimtime="00:00:36.02" resultid="3122" lane="8" heatid="7279" entrytime="00:00:36.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="384" reactiontime="+80" swimtime="00:00:32.96" resultid="3123" heatid="7334" entrytime="00:00:32.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MACHE" name="Masters Chełm" nation="POL" region="LBL">
          <CONTACT city="Chełm" email="elzbietadz@gmail.com" name="Dziwisz Elżbieta" phone="660429651" state="LUB" street="Lubelska 139D/13" zip="22-100" />
          <ATHLETES>
            <ATHLETE birthdate="1937-01-01" firstname="Tadeusz" gender="M" lastname="Wosk" nation="POL" athleteid="3125">
              <RESULTS>
                <RESULT eventid="1564" points="26" reactiontime="+134" swimtime="00:05:44.47" resultid="3128" lane="1" heatid="7054">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.47" />
                    <SPLIT distance="50" swimtime="00:01:14.98" />
                    <SPLIT distance="75" swimtime="00:01:58.92" />
                    <SPLIT distance="100" swimtime="00:02:43.98" />
                    <SPLIT distance="125" swimtime="00:03:29.72" />
                    <SPLIT distance="150" swimtime="00:04:15.12" />
                    <SPLIT distance="175" swimtime="00:04:58.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="28" reactiontime="+155" swimtime="00:02:33.89" resultid="3126" lane="3" heatid="6829">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:31.51" />
                    <SPLIT distance="50" swimtime="00:01:09.28" />
                    <SPLIT distance="75" swimtime="00:01:50.89" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="M 4" eventid="1598" reactiontime="+111" status="DSQ" swimtime="00:00:00.00" resultid="3129" lane="5" heatid="7071">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:48.77" />
                    <SPLIT distance="50" swimtime="00:01:49.69" />
                    <SPLIT distance="75" swimtime="00:02:49.17" />
                    <SPLIT distance="100" swimtime="00:03:45.74" />
                    <SPLIT distance="125" swimtime="00:04:42.17" />
                    <SPLIT distance="150" swimtime="00:05:38.73" />
                    <SPLIT distance="175" swimtime="00:06:21.83" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="przekroczony limit 10:00:00" eventid="1375" reactiontime="+112" status="DSQ" swimtime="00:00:00.00" resultid="3127" lane="2" heatid="6899">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.10" />
                    <SPLIT distance="50" swimtime="00:01:14.52" />
                    <SPLIT distance="75" swimtime="00:01:57.59" />
                    <SPLIT distance="100" swimtime="00:02:43.52" />
                    <SPLIT distance="125" swimtime="00:03:29.40" />
                    <SPLIT distance="150" swimtime="00:04:17.75" />
                    <SPLIT distance="175" swimtime="00:05:05.53" />
                    <SPLIT distance="200" swimtime="00:05:52.02" />
                    <SPLIT distance="225" swimtime="00:06:41.13" />
                    <SPLIT distance="250" swimtime="00:07:30.85" />
                    <SPLIT distance="275" swimtime="00:08:20.08" />
                    <SPLIT distance="300" swimtime="00:09:09.86" />
                    <SPLIT distance="325" swimtime="00:09:59.55" />
                    <SPLIT distance="350" swimtime="00:10:49.01" />
                    <SPLIT distance="375" swimtime="00:11:35.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1941-01-01" firstname="Janusz" gender="M" lastname="Golik" nation="POL" athleteid="3130">
              <RESULTS>
                <RESULT eventid="1462" points="79" reactiontime="+106" swimtime="00:01:57.02" resultid="3134" lane="1" heatid="7016" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.28" />
                    <SPLIT distance="50" swimtime="00:00:52.45" />
                    <SPLIT distance="75" swimtime="00:01:23.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="68" reactiontime="+125" swimtime="00:04:34.09" resultid="3132" lane="8" heatid="6870" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.82" />
                    <SPLIT distance="50" swimtime="00:00:58.12" />
                    <SPLIT distance="75" swimtime="00:01:30.26" />
                    <SPLIT distance="100" swimtime="00:02:04.79" />
                    <SPLIT distance="125" swimtime="00:02:40.25" />
                    <SPLIT distance="150" swimtime="00:03:15.73" />
                    <SPLIT distance="175" swimtime="00:03:53.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="107" reactiontime="+106" swimtime="00:00:48.30" resultid="3135" heatid="7282" entrytime="00:00:46.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="141" reactiontime="+110" swimtime="00:04:04.55" resultid="3133" lane="3" heatid="7003" entrytime="00:04:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.74" />
                    <SPLIT distance="50" swimtime="00:00:55.74" />
                    <SPLIT distance="75" swimtime="00:01:26.66" />
                    <SPLIT distance="100" swimtime="00:01:58.06" />
                    <SPLIT distance="125" swimtime="00:02:30.84" />
                    <SPLIT distance="150" swimtime="00:03:03.35" />
                    <SPLIT distance="175" swimtime="00:03:34.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="207" reactiontime="+114" swimtime="00:00:45.93" resultid="3131" lane="1" heatid="6856" entrytime="00:00:45.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="166" reactiontime="+111" swimtime="00:01:47.01" resultid="3136" lane="6" heatid="7304" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.27" />
                    <SPLIT distance="50" swimtime="00:00:50.57" />
                    <SPLIT distance="75" swimtime="00:01:19.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="Leszek" gender="M" lastname="Masłowski" nation="POL" athleteid="3140">
              <RESULTS>
                <RESULT eventid="1462" points="35" reactiontime="+119" swimtime="00:02:34.07" resultid="3144" lane="5" heatid="7015">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.57" />
                    <SPLIT distance="50" swimtime="00:01:02.43" />
                    <SPLIT distance="75" swimtime="00:01:45.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="59" reactiontime="+120" swimtime="00:04:51.83" resultid="3145" lane="4" heatid="7071">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.67" />
                    <SPLIT distance="50" swimtime="00:01:10.16" />
                    <SPLIT distance="75" swimtime="00:01:48.21" />
                    <SPLIT distance="100" swimtime="00:02:27.71" />
                    <SPLIT distance="125" swimtime="00:03:06.80" />
                    <SPLIT distance="150" swimtime="00:03:45.59" />
                    <SPLIT distance="175" swimtime="00:04:19.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="50" reactiontime="+67" swimtime="00:02:21.75" resultid="3147" lane="7" heatid="7318">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.43" />
                    <SPLIT distance="50" swimtime="00:01:09.28" />
                    <SPLIT distance="75" swimtime="00:01:45.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="50" reactiontime="+71" swimtime="00:05:09.00" resultid="3143" lane="5" heatid="6880">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:33.46" />
                    <SPLIT distance="50" swimtime="00:01:08.29" />
                    <SPLIT distance="75" swimtime="00:01:46.94" />
                    <SPLIT distance="100" swimtime="00:02:25.69" />
                    <SPLIT distance="125" swimtime="00:03:06.38" />
                    <SPLIT distance="150" swimtime="00:03:47.68" />
                    <SPLIT distance="175" swimtime="00:04:29.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="77" reactiontime="+110" swimtime="00:01:50.31" resultid="3142" lane="4" heatid="6829">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.39" />
                    <SPLIT distance="50" swimtime="00:00:50.51" />
                    <SPLIT distance="75" swimtime="00:01:20.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="61" reactiontime="+106" swimtime="00:00:58.32" resultid="3146" lane="8" heatid="7281">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="54" swimtime="00:02:15.16" resultid="3141" lane="2" heatid="6730">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.57" />
                    <SPLIT distance="50" swimtime="00:01:08.00" />
                    <SPLIT distance="75" swimtime="00:01:45.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Wiesław" gender="M" lastname="Wepa" nation="POL" athleteid="3148">
              <RESULTS>
                <RESULT eventid="1645" points="77" reactiontime="+86" swimtime="00:00:53.92" resultid="3154" lane="3" heatid="7282" entrytime="00:00:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="98" reactiontime="+101" swimtime="00:04:07.64" resultid="3153" lane="2" heatid="7073" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.69" />
                    <SPLIT distance="50" swimtime="00:00:49.80" />
                    <SPLIT distance="75" swimtime="00:01:24.76" />
                    <SPLIT distance="100" swimtime="00:02:00.14" />
                    <SPLIT distance="125" swimtime="00:02:35.78" />
                    <SPLIT distance="150" swimtime="00:03:08.75" />
                    <SPLIT distance="175" swimtime="00:03:38.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="154" reactiontime="+104" swimtime="00:03:57.81" resultid="3152" lane="4" heatid="7003" entrytime="00:04:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.42" />
                    <SPLIT distance="50" swimtime="00:00:53.39" />
                    <SPLIT distance="75" swimtime="00:01:23.99" />
                    <SPLIT distance="100" swimtime="00:01:54.39" />
                    <SPLIT distance="125" swimtime="00:02:25.38" />
                    <SPLIT distance="150" swimtime="00:02:57.35" />
                    <SPLIT distance="175" swimtime="00:03:28.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="154" reactiontime="+88" swimtime="00:01:49.86" resultid="3155" heatid="7303" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.74" />
                    <SPLIT distance="50" swimtime="00:00:53.37" />
                    <SPLIT distance="75" swimtime="00:01:22.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="177" reactiontime="+98" swimtime="00:00:48.34" resultid="3150" lane="2" heatid="6856" entrytime="00:00:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" status="DNS" swimtime="00:00:00.00" resultid="3151" lane="6" heatid="6900" entrytime="00:07:30.00" />
                <RESULT comment="przekroczony limit 30:00:00" eventid="1143" status="DSQ" swimtime="00:33:09.00" resultid="3149" lane="7" heatid="6749" entrytime="00:29:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1926-01-01" firstname="Barbara" gender="F" lastname="Korol" nation="POL" athleteid="3156">
              <RESULTS>
                <RESULT eventid="1187" points="6" swimtime="00:04:44.20" resultid="3157" lane="4" heatid="6821">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:01:04.95" />
                    <SPLIT distance="50" swimtime="00:02:18.47" />
                    <SPLIT distance="75" swimtime="00:03:26.46" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1479" points="19" reactiontime="+99" swimtime="00:01:43.40" resultid="3158" lane="5" heatid="7024">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:49.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="10" swimtime="00:01:48.30" resultid="3160" heatid="7328">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:49.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="18" reactiontime="+107" swimtime="00:03:43.31" resultid="3159" lane="5" heatid="7312">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:51.85" />
                    <SPLIT distance="50" swimtime="00:01:49.27" />
                    <SPLIT distance="75" swimtime="00:02:47.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-01" firstname="Alicja" gender="F" lastname="Wątrobińska" nation="POL" athleteid="3161">
              <RESULTS>
                <RESULT eventid="1641" points="47" reactiontime="+117" swimtime="00:01:10.49" resultid="3167" lane="5" heatid="7275" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1409" points="75" reactiontime="+127" swimtime="00:05:31.09" resultid="3165" lane="5" heatid="6997">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:38.49" />
                    <SPLIT distance="50" swimtime="00:01:19.98" />
                    <SPLIT distance="75" swimtime="00:02:03.20" />
                    <SPLIT distance="100" swimtime="00:02:45.12" />
                    <SPLIT distance="125" swimtime="00:03:28.13" />
                    <SPLIT distance="150" swimtime="00:04:09.79" />
                    <SPLIT distance="175" swimtime="00:04:51.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="43" reactiontime="+95" swimtime="00:01:18.48" resultid="3166" lane="8" heatid="7026" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:39.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="62" reactiontime="+122" swimtime="00:02:28.29" resultid="3162" lane="5" heatid="6723">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.58" />
                    <SPLIT distance="50" swimtime="00:01:14.87" />
                    <SPLIT distance="75" swimtime="00:01:54.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="81" reactiontime="+103" swimtime="00:01:09.92" resultid="3164" lane="4" heatid="6847">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="72" reactiontime="+107" swimtime="00:00:57.49" resultid="3168" lane="3" heatid="7328" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="69" reactiontime="+116" swimtime="00:02:08.57" resultid="3163" lane="3" heatid="6821">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.35" />
                    <SPLIT distance="50" swimtime="00:01:01.64" />
                    <SPLIT distance="75" swimtime="00:01:35.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-01" firstname="Dorota" gender="F" lastname="Czerniakiewicz" nation="POL" athleteid="3169">
              <RESULTS>
                <RESULT eventid="1409" points="188" reactiontime="+89" swimtime="00:04:04.54" resultid="3173" lane="2" heatid="6997">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.96" />
                    <SPLIT distance="50" swimtime="00:00:55.13" />
                    <SPLIT distance="75" swimtime="00:01:25.06" />
                    <SPLIT distance="100" swimtime="00:01:56.83" />
                    <SPLIT distance="125" swimtime="00:02:28.52" />
                    <SPLIT distance="150" swimtime="00:03:00.36" />
                    <SPLIT distance="175" swimtime="00:03:32.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="196" reactiontime="+90" swimtime="00:01:51.98" resultid="3175" lane="2" heatid="7295">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.65" />
                    <SPLIT distance="50" swimtime="00:00:52.98" />
                    <SPLIT distance="75" swimtime="00:01:22.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="208" reactiontime="+81" swimtime="00:00:51.11" resultid="3172" heatid="6850" entrytime="00:00:51.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="163" reactiontime="+86" swimtime="00:00:43.85" resultid="3176" lane="4" heatid="7327">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="133" reactiontime="+105" swimtime="00:00:54.11" resultid="3174" lane="3" heatid="7024">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="147" reactiontime="+83" swimtime="00:01:51.39" resultid="3170" lane="1" heatid="6724" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.98" />
                    <SPLIT distance="50" swimtime="00:00:51.59" />
                    <SPLIT distance="75" swimtime="00:01:22.58" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="za nieprawdiłowy strój" eventid="1187" reactiontime="+85" status="DSQ" swimtime="00:00:00.00" resultid="3171" heatid="6822">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.07" />
                    <SPLIT distance="50" swimtime="00:00:49.40" />
                    <SPLIT distance="75" swimtime="00:01:18.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-10-28" firstname="Elżbieta" gender="F" lastname="Dziwisz" nation="POL" athleteid="3177">
              <RESULTS>
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="3181" heatid="7026" entrytime="00:00:59.00" />
                <RESULT eventid="1679" status="DNS" swimtime="00:00:00.00" resultid="3182" lane="5" heatid="7296" entrytime="00:02:01.00" />
                <RESULT eventid="1409" status="DNS" swimtime="00:00:00.00" resultid="3180" lane="4" heatid="6998" entrytime="00:04:29.00" />
                <RESULT eventid="1290" status="DNS" swimtime="00:00:00.00" resultid="3179" lane="6" heatid="6876" entrytime="00:04:30.00" />
                <RESULT eventid="1222" status="DNS" swimtime="00:00:00.00" resultid="3178" lane="4" heatid="6848" entrytime="00:00:58.00" />
                <RESULT eventid="1713" status="DNS" swimtime="00:00:00.00" resultid="3183" lane="8" heatid="7314" entrytime="00:02:02.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1177" status="DNS" swimtime="00:00:00.00" resultid="3188" lane="6" heatid="6807">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3140" number="1" />
                    <RELAYPOSITION athleteid="3148" number="3" />
                    <RELAYPOSITION athleteid="3130" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1341" status="DNS" swimtime="00:00:00.00" resultid="3189" lane="2" heatid="6985">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3148" number="2" />
                    <RELAYPOSITION athleteid="3130" number="3" />
                    <RELAYPOSITION athleteid="3148" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="3186" heatid="6813">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.53" />
                    <SPLIT distance="100" swimtime="00:03:04.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3156" number="1" />
                    <RELAYPOSITION athleteid="3177" number="2" />
                    <RELAYPOSITION athleteid="3161" number="3" />
                    <RELAYPOSITION athleteid="3169" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1324" points="48" reactiontime="+90" swimtime="00:04:57.18" resultid="3187" lane="8" heatid="6979">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:50.01" />
                    <SPLIT distance="50" swimtime="00:01:04.63" />
                    <SPLIT distance="75" swimtime="00:02:22.44" />
                    <SPLIT distance="100" swimtime="00:01:26.35" />
                    <SPLIT distance="125" swimtime="00:03:32.46" />
                    <SPLIT distance="150" swimtime="00:03:07.76" />
                    <SPLIT distance="175" swimtime="00:04:28.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3156" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="3177" number="2" />
                    <RELAYPOSITION athleteid="3161" number="3" />
                    <RELAYPOSITION athleteid="3169" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="319" agemin="280" agetotalmax="-1" agetotalmin="-1" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1615" swimtime="00:04:55.81" resultid="3190" lane="5" heatid="7440">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:53.79" />
                    <SPLIT distance="50" swimtime="00:01:53.21" />
                    <SPLIT distance="75" swimtime="00:02:19.59" />
                    <SPLIT distance="100" swimtime="00:02:54.77" />
                    <SPLIT distance="125" swimtime="00:03:20.09" />
                    <SPLIT distance="150" swimtime="00:03:47.74" />
                    <SPLIT distance="175" swimtime="00:04:20.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3156" number="1" />
                    <RELAYPOSITION athleteid="3161" number="2" />
                    <RELAYPOSITION athleteid="3130" number="3" reactiontime="+138" />
                    <RELAYPOSITION athleteid="3125" number="4" reactiontime="+104" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1815" status="DNS" swimtime="00:00:00.00" resultid="3191" lane="5" heatid="7502">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3156" number="1" />
                    <RELAYPOSITION athleteid="3161" number="2" />
                    <RELAYPOSITION athleteid="3130" number="3" />
                    <RELAYPOSITION athleteid="3125" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="1615" reactiontime="+99" swimtime="00:03:31.49" resultid="3184" lane="7" heatid="7441">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.87" />
                    <SPLIT distance="50" swimtime="00:00:45.26" />
                    <SPLIT distance="75" swimtime="00:01:05.24" />
                    <SPLIT distance="100" swimtime="00:01:26.71" />
                    <SPLIT distance="125" swimtime="00:01:47.38" />
                    <SPLIT distance="150" swimtime="00:02:12.17" />
                    <SPLIT distance="175" swimtime="00:02:49.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3177" number="1" reactiontime="+99" />
                    <RELAYPOSITION athleteid="3148" number="2" reactiontime="+102" />
                    <RELAYPOSITION athleteid="3140" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="3169" number="4" reactiontime="+191" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1815" status="DNS" swimtime="00:00:00.00" resultid="3185" lane="6" heatid="7502">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3177" number="1" />
                    <RELAYPOSITION athleteid="3148" number="2" />
                    <RELAYPOSITION athleteid="3140" number="3" />
                    <RELAYPOSITION athleteid="3169" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="CPCHO" name="Centrum Park Chojnice" nation="POL">
          <CONTACT city="Chojnice" name="Centrum Park Chojnice" state="POMOR" street="Huberta Wagnera 1" zip="89-604" />
          <ATHLETES>
            <ATHLETE birthdate="1986-09-12" firstname="Tomasz" gender="M" lastname="Żmiejko" nation="POL" athleteid="3204">
              <RESULTS>
                <RESULT eventid="1462" points="306" reactiontime="+77" swimtime="00:01:14.73" resultid="3207" lane="1" heatid="7020" entrytime="00:01:15.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.67" />
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                    <SPLIT distance="75" swimtime="00:00:53.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="410" reactiontime="+74" swimtime="00:01:03.29" resultid="3206" lane="6" heatid="6841" entrytime="00:01:03.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.43" />
                    <SPLIT distance="50" swimtime="00:00:30.15" />
                    <SPLIT distance="75" swimtime="00:00:46.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="433" reactiontime="+73" swimtime="00:00:30.33" resultid="3208" lane="3" heatid="7290" entrytime="00:00:29.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="298" reactiontime="+75" swimtime="00:01:16.57" resultid="3205" lane="4" heatid="6738" entrytime="00:01:15.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.17" />
                    <SPLIT distance="50" swimtime="00:00:36.51" />
                    <SPLIT distance="75" swimtime="00:00:59.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="418" reactiontime="+71" swimtime="00:00:28.44" resultid="3209" lane="6" heatid="7348" entrytime="00:00:27.99">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-03-08" firstname="Barbara" gender="F" lastname="Błaszkowska" nation="POL" athleteid="3210">
              <RESULTS>
                <RESULT eventid="1126" points="91" swimtime="00:34:54.28" resultid="3211" lane="6" heatid="6746" entrytime="00:37:40.20" />
                <RESULT eventid="1358" points="86" reactiontime="+141" swimtime="00:09:05.09" resultid="3213" lane="7" heatid="6894" entrytime="00:09:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.49" />
                    <SPLIT distance="50" swimtime="00:00:58.91" />
                    <SPLIT distance="75" swimtime="00:01:32.18" />
                    <SPLIT distance="100" swimtime="00:02:05.52" />
                    <SPLIT distance="125" swimtime="00:02:40.26" />
                    <SPLIT distance="150" swimtime="00:03:15.00" />
                    <SPLIT distance="175" swimtime="00:03:50.00" />
                    <SPLIT distance="200" swimtime="00:04:23.99" />
                    <SPLIT distance="225" swimtime="00:04:59.31" />
                    <SPLIT distance="250" swimtime="00:05:33.72" />
                    <SPLIT distance="275" swimtime="00:06:09.29" />
                    <SPLIT distance="300" swimtime="00:06:43.62" />
                    <SPLIT distance="325" swimtime="00:07:19.06" />
                    <SPLIT distance="350" swimtime="00:07:54.88" />
                    <SPLIT distance="375" swimtime="00:08:31.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="78" reactiontime="+111" swimtime="00:02:31.87" resultid="3215" lane="1" heatid="7296" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:33.11" />
                    <SPLIT distance="50" swimtime="00:01:09.85" />
                    <SPLIT distance="75" swimtime="00:01:50.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="75" reactiontime="+125" swimtime="00:04:31.57" resultid="3214" lane="8" heatid="7049" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.52" />
                    <SPLIT distance="50" swimtime="00:00:59.75" />
                    <SPLIT distance="75" swimtime="00:01:34.46" />
                    <SPLIT distance="100" swimtime="00:02:09.72" />
                    <SPLIT distance="125" swimtime="00:02:44.78" />
                    <SPLIT distance="150" swimtime="00:03:20.61" />
                    <SPLIT distance="175" swimtime="00:03:56.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="69" reactiontime="+133" swimtime="00:02:08.49" resultid="3212" lane="3" heatid="6822" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.18" />
                    <SPLIT distance="50" swimtime="00:00:58.02" />
                    <SPLIT distance="75" swimtime="00:01:32.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DEGDY" name="KS Delfin Gdynia" nation="POL" region="GD">
          <ATHLETES>
            <ATHLETE birthdate="1971-11-04" firstname="Jakub" gender="M" lastname="Mańczak" nation="POL" license="S01910200065" athleteid="3217">
              <RESULTS>
                <RESULT eventid="1645" points="484" reactiontime="+76" swimtime="00:00:29.24" resultid="3220" lane="8" heatid="7291" entrytime="00:00:29.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="444" reactiontime="+75" swimtime="00:01:06.05" resultid="3219" lane="1" heatid="7021" entrytime="00:01:09.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.80" />
                    <SPLIT distance="50" swimtime="00:00:30.64" />
                    <SPLIT distance="75" swimtime="00:00:48.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="506" reactiontime="+75" swimtime="00:00:26.69" resultid="3221" lane="5" heatid="7348" entrytime="00:00:27.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.99" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="M 10" eventid="1273" reactiontime="+88" status="DSQ" swimtime="00:02:41.36" resultid="3218" lane="3" heatid="6873" entrytime="00:02:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.12" />
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                    <SPLIT distance="75" swimtime="00:00:52.79" />
                    <SPLIT distance="100" swimtime="00:01:12.87" />
                    <SPLIT distance="125" swimtime="00:01:35.09" />
                    <SPLIT distance="150" swimtime="00:01:57.34" />
                    <SPLIT distance="175" swimtime="00:02:19.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-24" firstname="Aleksandra" gender="F" lastname="Sypniewska" nation="POL" license="S01910100045" athleteid="3222">
              <RESULTS>
                <RESULT eventid="1058" points="368" swimtime="00:11:28.93" resultid="3223" lane="2" heatid="6715" entrytime="00:11:30.00" />
                <RESULT eventid="1358" points="376" reactiontime="+96" swimtime="00:05:34.54" resultid="3224" lane="8" heatid="6898" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.35" />
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                    <SPLIT distance="75" swimtime="00:00:53.19" />
                    <SPLIT distance="100" swimtime="00:01:12.90" />
                    <SPLIT distance="125" swimtime="00:01:33.48" />
                    <SPLIT distance="150" swimtime="00:01:54.14" />
                    <SPLIT distance="175" swimtime="00:02:15.40" />
                    <SPLIT distance="200" swimtime="00:02:37.29" />
                    <SPLIT distance="225" swimtime="00:02:59.24" />
                    <SPLIT distance="250" swimtime="00:03:21.29" />
                    <SPLIT distance="275" swimtime="00:03:43.73" />
                    <SPLIT distance="300" swimtime="00:04:05.98" />
                    <SPLIT distance="325" swimtime="00:04:28.16" />
                    <SPLIT distance="350" swimtime="00:04:50.36" />
                    <SPLIT distance="375" swimtime="00:05:12.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="413" reactiontime="+90" swimtime="00:02:34.11" resultid="3225" lane="8" heatid="7053" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.17" />
                    <SPLIT distance="50" swimtime="00:00:34.04" />
                    <SPLIT distance="75" swimtime="00:00:52.63" />
                    <SPLIT distance="100" swimtime="00:01:11.80" />
                    <SPLIT distance="125" swimtime="00:01:31.59" />
                    <SPLIT distance="150" swimtime="00:01:52.19" />
                    <SPLIT distance="175" swimtime="00:02:13.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ENTRE" name="ENTRE.PL Team" nation="POL">
          <CONTACT name="Paweł Zach" />
          <ATHLETES>
            <ATHLETE birthdate="1968-06-21" firstname="Paweł" gender="M" lastname="Zach" nation="POL" athleteid="3227">
              <RESULTS>
                <RESULT eventid="1696" points="137" reactiontime="+88" swimtime="00:01:54.10" resultid="3233" heatid="7304" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.35" />
                    <SPLIT distance="50" swimtime="00:00:50.90" />
                    <SPLIT distance="75" swimtime="00:01:23.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="197" reactiontime="+89" swimtime="00:06:17.71" resultid="3230" lane="2" heatid="6902" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.51" />
                    <SPLIT distance="50" swimtime="00:00:41.95" />
                    <SPLIT distance="75" swimtime="00:01:05.58" />
                    <SPLIT distance="100" swimtime="00:01:29.49" />
                    <SPLIT distance="125" swimtime="00:01:53.73" />
                    <SPLIT distance="150" swimtime="00:02:17.83" />
                    <SPLIT distance="175" swimtime="00:02:42.14" />
                    <SPLIT distance="200" swimtime="00:03:06.43" />
                    <SPLIT distance="225" swimtime="00:03:29.79" />
                    <SPLIT distance="250" swimtime="00:03:54.66" />
                    <SPLIT distance="275" swimtime="00:04:18.69" />
                    <SPLIT distance="300" swimtime="00:04:43.06" />
                    <SPLIT distance="325" swimtime="00:05:06.98" />
                    <SPLIT distance="350" swimtime="00:05:31.37" />
                    <SPLIT distance="375" swimtime="00:05:55.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="211" reactiontime="+84" swimtime="00:02:52.92" resultid="3232" lane="3" heatid="7057" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.48" />
                    <SPLIT distance="50" swimtime="00:00:39.63" />
                    <SPLIT distance="75" swimtime="00:01:01.07" />
                    <SPLIT distance="100" swimtime="00:01:23.42" />
                    <SPLIT distance="125" swimtime="00:01:45.93" />
                    <SPLIT distance="150" swimtime="00:02:09.03" />
                    <SPLIT distance="175" swimtime="00:02:31.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="226" reactiontime="+89" swimtime="00:00:34.89" resultid="3234" lane="5" heatid="7338" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="191" reactiontime="+96" swimtime="00:01:21.58" resultid="3229" heatid="6833" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.27" />
                    <SPLIT distance="50" swimtime="00:00:38.66" />
                    <SPLIT distance="75" swimtime="00:01:00.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" status="DNS" swimtime="00:00:00.00" resultid="3231" heatid="7035" entrytime="00:00:47.00" />
                <RESULT eventid="1143" status="DNF" swimtime="00:00:00.00" resultid="3228" lane="7" heatid="6750" entrytime="00:24:20.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SOKOL" name="Sokół Kolbuszowa" nation="POL">
          <CONTACT email="bartek_swim@interia.pl" name="Pietryka Bartosz" phone="604620876" />
          <ATHLETES>
            <ATHLETE birthdate="1972-02-11" firstname="Witold" gender="M" lastname="Rado" nation="POL" athleteid="3236">
              <RESULTS>
                <RESULT eventid="1143" points="378" swimtime="00:20:09.00" resultid="3237" lane="3" heatid="6752" entrytime="00:19:15.00" />
                <RESULT eventid="1462" points="391" reactiontime="+85" swimtime="00:01:08.92" resultid="3240" lane="5" heatid="7022" entrytime="00:01:05.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.13" />
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                    <SPLIT distance="75" swimtime="00:00:50.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="386" reactiontime="+94" swimtime="00:05:02.03" resultid="3239" lane="7" heatid="6909" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.69" />
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                    <SPLIT distance="75" swimtime="00:00:50.99" />
                    <SPLIT distance="100" swimtime="00:01:09.62" />
                    <SPLIT distance="125" swimtime="00:01:28.53" />
                    <SPLIT distance="150" swimtime="00:01:47.92" />
                    <SPLIT distance="175" swimtime="00:02:07.57" />
                    <SPLIT distance="200" swimtime="00:02:27.13" />
                    <SPLIT distance="225" swimtime="00:02:46.68" />
                    <SPLIT distance="250" swimtime="00:03:06.14" />
                    <SPLIT distance="275" swimtime="00:03:25.65" />
                    <SPLIT distance="300" swimtime="00:03:45.11" />
                    <SPLIT distance="325" swimtime="00:04:04.59" />
                    <SPLIT distance="350" swimtime="00:04:24.35" />
                    <SPLIT distance="375" swimtime="00:04:43.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="310" reactiontime="+80" swimtime="00:01:17.61" resultid="3243" lane="8" heatid="7325" entrytime="00:01:10.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.40" />
                    <SPLIT distance="50" swimtime="00:00:37.77" />
                    <SPLIT distance="75" swimtime="00:00:57.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="379" reactiontime="+89" swimtime="00:02:22.25" resultid="3241" lane="1" heatid="7065" entrytime="00:02:10.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.17" />
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                    <SPLIT distance="75" swimtime="00:00:49.84" />
                    <SPLIT distance="100" swimtime="00:01:08.26" />
                    <SPLIT distance="125" swimtime="00:01:26.34" />
                    <SPLIT distance="150" swimtime="00:01:45.20" />
                    <SPLIT distance="175" swimtime="00:02:04.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="376" reactiontime="+80" swimtime="00:01:05.17" resultid="3238" heatid="6843" entrytime="00:01:00.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.63" />
                    <SPLIT distance="50" swimtime="00:00:31.03" />
                    <SPLIT distance="75" swimtime="00:00:47.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="3242" lane="6" heatid="7292" entrytime="00:00:28.85" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-07-20" firstname="Bartosz" gender="M" lastname="Pietryka" nation="POL" athleteid="3244">
              <RESULTS>
                <RESULT eventid="1730" points="480" reactiontime="+82" swimtime="00:01:07.07" resultid="3248" lane="7" heatid="7326" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.27" />
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                    <SPLIT distance="75" swimtime="00:00:50.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="490" reactiontime="+77" swimtime="00:00:31.02" resultid="3246" lane="1" heatid="7042" entrytime="00:00:30.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="469" reactiontime="+81" swimtime="00:01:04.84" resultid="3245" lane="8" heatid="7023" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.17" />
                    <SPLIT distance="50" swimtime="00:00:29.23" />
                    <SPLIT distance="75" swimtime="00:00:46.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="3247" heatid="7293" entrytime="00:00:28.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" name="niezrzeszeni" nation="POL" region="LOD">
          <CONTACT city="łódź" name="Ewa Cieplucha" phone="604627966" street="Retkińska 74 m 18" zip="94-004" />
          <ATHLETES>
            <ATHLETE birthdate="1981-05-26" firstname="Ewa" gender="F" lastname="Cieplucha" nation="POL" athleteid="3250">
              <RESULTS>
                <RESULT eventid="1479" points="471" reactiontime="+64" swimtime="00:00:35.54" resultid="3252" lane="4" heatid="7029" entrytime="00:00:39.13">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="431" reactiontime="+69" swimtime="00:01:17.79" resultid="3253" lane="2" heatid="7316" entrytime="00:01:25.13">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.97" />
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                    <SPLIT distance="75" swimtime="00:00:56.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="356" reactiontime="+87" swimtime="00:01:14.55" resultid="3251" heatid="6827" entrytime="00:01:13.13">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.44" />
                    <SPLIT distance="50" swimtime="00:00:34.92" />
                    <SPLIT distance="75" swimtime="00:00:54.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-07-29" firstname="Magdalena" gender="F" lastname="Piątkiewicz" nation="POL" athleteid="3254">
              <RESULTS>
                <RESULT eventid="1713" points="402" reactiontime="+78" swimtime="00:01:19.61" resultid="3257" lane="5" heatid="7316" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.27" />
                    <SPLIT distance="50" swimtime="00:00:39.38" />
                    <SPLIT distance="75" swimtime="00:00:59.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="448" reactiontime="+74" swimtime="00:00:36.14" resultid="3256" heatid="7030" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="444" reactiontime="+90" swimtime="00:00:31.41" resultid="3258" lane="4" heatid="7332" entrytime="00:00:34.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="393" reactiontime="+95" swimtime="00:01:12.16" resultid="3255" lane="6" heatid="6827" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.84" />
                    <SPLIT distance="50" swimtime="00:00:35.23" />
                    <SPLIT distance="75" swimtime="00:00:53.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="VIELB" name="Victory Masters Elbląg 1" nation="POL" region="WAR">
          <CONTACT city="ELBLĄG" email="lateccy@o2.pl" name="Latecki Grzegorz" state="WAR" zip="82-300" />
          <ATHLETES>
            <ATHLETE birthdate="1965-03-12" firstname="Grzegorz" gender="M" lastname="Latecki" nation="POL" athleteid="3260">
              <RESULTS>
                <RESULT eventid="1645" points="500" reactiontime="+75" swimtime="00:00:28.92" resultid="3266" lane="4" heatid="7290" entrytime="00:00:29.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="421" reactiontime="+80" swimtime="00:02:32.31" resultid="3265" lane="3" heatid="7078" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.20" />
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                    <SPLIT distance="75" swimtime="00:00:52.17" />
                    <SPLIT distance="100" swimtime="00:01:12.05" />
                    <SPLIT distance="125" swimtime="00:01:34.13" />
                    <SPLIT distance="150" swimtime="00:01:57.43" />
                    <SPLIT distance="175" swimtime="00:02:15.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="438" reactiontime="+70" swimtime="00:00:32.22" resultid="3264" lane="3" heatid="7040" entrytime="00:00:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="484" reactiontime="+76" swimtime="00:00:27.09" resultid="3267" lane="4" heatid="7348" entrytime="00:00:27.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="448" reactiontime="+85" swimtime="00:00:35.51" resultid="3263" lane="2" heatid="6863" entrytime="00:00:36.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="414" reactiontime="+80" swimtime="00:01:08.62" resultid="3261" lane="1" heatid="6741" entrytime="00:01:10.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.27" />
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                    <SPLIT distance="75" swimtime="00:00:51.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="478" reactiontime="+78" swimtime="00:01:00.17" resultid="3262" lane="4" heatid="6842" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.73" />
                    <SPLIT distance="50" swimtime="00:00:29.24" />
                    <SPLIT distance="75" swimtime="00:00:44.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-08-31" firstname="Karolina" gender="F" lastname="Karaś" nation="POL" athleteid="3268">
              <RESULTS>
                <RESULT eventid="1358" points="139" reactiontime="+111" swimtime="00:07:45.70" resultid="3270" lane="7" heatid="6895" entrytime="00:07:26.23">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.60" />
                    <SPLIT distance="50" swimtime="00:00:53.93" />
                    <SPLIT distance="75" swimtime="00:01:22.25" />
                    <SPLIT distance="100" swimtime="00:01:51.68" />
                    <SPLIT distance="125" swimtime="00:02:21.02" />
                    <SPLIT distance="150" swimtime="00:02:50.91" />
                    <SPLIT distance="175" swimtime="00:03:20.65" />
                    <SPLIT distance="200" swimtime="00:03:49.96" />
                    <SPLIT distance="225" swimtime="00:04:20.52" />
                    <SPLIT distance="250" swimtime="00:04:50.16" />
                    <SPLIT distance="275" swimtime="00:05:20.30" />
                    <SPLIT distance="300" swimtime="00:05:50.32" />
                    <SPLIT distance="325" swimtime="00:06:20.36" />
                    <SPLIT distance="350" swimtime="00:06:49.34" />
                    <SPLIT distance="375" swimtime="00:07:17.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="120" reactiontime="+108" swimtime="00:01:46.97" resultid="3269" heatid="6824" entrytime="00:01:37.65">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.15" />
                    <SPLIT distance="50" swimtime="00:00:53.05" />
                    <SPLIT distance="75" swimtime="00:01:20.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="150" reactiontime="+87" swimtime="00:00:45.07" resultid="3272" lane="2" heatid="7330" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="134" reactiontime="+99" swimtime="00:03:44.35" resultid="3271" lane="8" heatid="7050" entrytime="00:03:35.76">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.43" />
                    <SPLIT distance="50" swimtime="00:00:52.74" />
                    <SPLIT distance="75" swimtime="00:01:20.73" />
                    <SPLIT distance="100" swimtime="00:01:50.27" />
                    <SPLIT distance="125" swimtime="00:02:19.98" />
                    <SPLIT distance="150" swimtime="00:02:48.97" />
                    <SPLIT distance="175" swimtime="00:03:17.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-05-05" firstname="Beata" gender="F" lastname="Karaś" nation="POL" athleteid="3273">
              <RESULTS>
                <RESULT eventid="1126" points="191" swimtime="00:27:16.56" resultid="3274" lane="1" heatid="6747" entrytime="00:26:00.00" />
                <RESULT eventid="1781" points="141" reactiontime="+106" swimtime="00:08:37.01" resultid="3279" lane="4" heatid="7355" entrytime="00:08:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.53" />
                    <SPLIT distance="50" swimtime="00:00:53.18" />
                    <SPLIT distance="75" swimtime="00:01:25.63" />
                    <SPLIT distance="100" swimtime="00:01:58.59" />
                    <SPLIT distance="125" swimtime="00:02:32.97" />
                    <SPLIT distance="150" swimtime="00:03:06.29" />
                    <SPLIT distance="175" swimtime="00:03:38.63" />
                    <SPLIT distance="200" swimtime="00:04:11.77" />
                    <SPLIT distance="225" swimtime="00:04:49.97" />
                    <SPLIT distance="250" swimtime="00:05:29.27" />
                    <SPLIT distance="275" swimtime="00:06:10.41" />
                    <SPLIT distance="300" swimtime="00:06:50.96" />
                    <SPLIT distance="325" swimtime="00:07:18.98" />
                    <SPLIT distance="350" swimtime="00:07:45.85" />
                    <SPLIT distance="375" swimtime="00:08:12.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1445" points="118" reactiontime="+102" swimtime="00:01:55.34" resultid="3277" lane="1" heatid="7013" entrytime="00:01:47.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.26" />
                    <SPLIT distance="50" swimtime="00:00:52.36" />
                    <SPLIT distance="75" swimtime="00:01:23.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="124" reactiontime="+109" swimtime="00:04:09.00" resultid="3275" lane="6" heatid="6868" entrytime="00:03:54.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.18" />
                    <SPLIT distance="50" swimtime="00:00:54.84" />
                    <SPLIT distance="75" swimtime="00:01:25.60" />
                    <SPLIT distance="100" swimtime="00:01:57.28" />
                    <SPLIT distance="125" swimtime="00:02:29.46" />
                    <SPLIT distance="150" swimtime="00:03:01.84" />
                    <SPLIT distance="175" swimtime="00:03:35.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1581" points="142" reactiontime="+104" swimtime="00:04:05.87" resultid="3278" lane="6" heatid="7068" entrytime="00:03:51.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.22" />
                    <SPLIT distance="50" swimtime="00:00:52.90" />
                    <SPLIT distance="75" swimtime="00:01:27.35" />
                    <SPLIT distance="100" swimtime="00:02:00.10" />
                    <SPLIT distance="125" swimtime="00:02:37.10" />
                    <SPLIT distance="150" swimtime="00:03:14.92" />
                    <SPLIT distance="175" swimtime="00:03:41.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="187" reactiontime="+115" swimtime="00:07:01.66" resultid="3276" heatid="6896" entrytime="00:06:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.21" />
                    <SPLIT distance="50" swimtime="00:00:48.02" />
                    <SPLIT distance="75" swimtime="00:01:13.82" />
                    <SPLIT distance="100" swimtime="00:01:40.56" />
                    <SPLIT distance="125" swimtime="00:02:07.61" />
                    <SPLIT distance="150" swimtime="00:02:34.90" />
                    <SPLIT distance="175" swimtime="00:03:01.65" />
                    <SPLIT distance="200" swimtime="00:03:28.72" />
                    <SPLIT distance="225" swimtime="00:03:55.71" />
                    <SPLIT distance="250" swimtime="00:04:23.26" />
                    <SPLIT distance="275" swimtime="00:04:50.66" />
                    <SPLIT distance="300" swimtime="00:05:17.75" />
                    <SPLIT distance="325" swimtime="00:05:43.89" />
                    <SPLIT distance="350" swimtime="00:06:10.72" />
                    <SPLIT distance="375" swimtime="00:06:37.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-03-30" firstname="Henryk" gender="M" lastname="Iszoro" nation="POL" athleteid="3280">
              <RESULTS>
                <RESULT eventid="1411" points="110" reactiontime="+115" swimtime="00:04:26.03" resultid="3282" heatid="7003" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.69" />
                    <SPLIT distance="50" swimtime="00:00:59.62" />
                    <SPLIT distance="75" swimtime="00:01:31.80" />
                    <SPLIT distance="100" swimtime="00:02:06.87" />
                    <SPLIT distance="125" swimtime="00:02:40.17" />
                    <SPLIT distance="150" swimtime="00:03:14.98" />
                    <SPLIT distance="175" swimtime="00:03:49.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="196" reactiontime="+124" swimtime="00:00:46.78" resultid="3281" lane="1" heatid="6855" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="144" reactiontime="+87" swimtime="00:01:52.38" resultid="3283" lane="1" heatid="7303" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.86" />
                    <SPLIT distance="50" swimtime="00:00:51.16" />
                    <SPLIT distance="75" swimtime="00:01:20.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-06-30" firstname="Andrzej" gender="M" lastname="Pasieczny" nation="POL" athleteid="3284">
              <RESULTS>
                <RESULT comment="Rekord Polski " eventid="1273" points="474" reactiontime="+93" swimtime="00:02:23.62" resultid="3285" lane="1" heatid="6874" entrytime="00:02:31.87">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.56" />
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                    <SPLIT distance="75" swimtime="00:00:49.42" />
                    <SPLIT distance="100" swimtime="00:01:07.51" />
                    <SPLIT distance="125" swimtime="00:01:25.59" />
                    <SPLIT distance="150" swimtime="00:01:44.15" />
                    <SPLIT distance="175" swimtime="00:02:02.85" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1462" points="480" reactiontime="+80" swimtime="00:01:04.35" resultid="3287" heatid="7022" entrytime="00:01:07.09">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.92" />
                    <SPLIT distance="50" swimtime="00:00:30.45" />
                    <SPLIT distance="75" swimtime="00:00:47.14" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1564" points="496" reactiontime="+86" swimtime="00:02:10.03" resultid="3288" heatid="7065" entrytime="00:02:12.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.30" />
                    <SPLIT distance="50" swimtime="00:00:30.64" />
                    <SPLIT distance="75" swimtime="00:00:46.92" />
                    <SPLIT distance="100" swimtime="00:01:03.83" />
                    <SPLIT distance="125" swimtime="00:01:20.42" />
                    <SPLIT distance="150" swimtime="00:01:37.23" />
                    <SPLIT distance="175" swimtime="00:01:53.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="468" reactiontime="+78" swimtime="00:00:29.56" resultid="3289" lane="7" heatid="7289" entrytime="00:00:31.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" status="DNS" swimtime="00:00:00.00" resultid="3286" lane="2" heatid="6908" entrytime="00:04:50.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-11-18" firstname="Tomasz" gender="M" lastname="Gleb" nation="POL" athleteid="3290">
              <RESULTS>
                <RESULT eventid="1075" points="321" swimtime="00:11:09.85" resultid="3291" lane="1" heatid="6721" entrytime="00:11:15.00" />
                <RESULT eventid="1375" points="347" reactiontime="+87" swimtime="00:05:13.12" resultid="3293" lane="8" heatid="6907" entrytime="00:05:22.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.96" />
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                    <SPLIT distance="75" swimtime="00:00:51.21" />
                    <SPLIT distance="100" swimtime="00:01:10.20" />
                    <SPLIT distance="125" swimtime="00:01:29.40" />
                    <SPLIT distance="150" swimtime="00:01:48.85" />
                    <SPLIT distance="175" swimtime="00:02:08.96" />
                    <SPLIT distance="200" swimtime="00:02:29.55" />
                    <SPLIT distance="225" swimtime="00:02:50.06" />
                    <SPLIT distance="250" swimtime="00:03:10.27" />
                    <SPLIT distance="275" swimtime="00:03:30.66" />
                    <SPLIT distance="300" swimtime="00:03:51.10" />
                    <SPLIT distance="325" swimtime="00:04:11.76" />
                    <SPLIT distance="350" swimtime="00:04:32.24" />
                    <SPLIT distance="375" swimtime="00:04:52.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="348" reactiontime="+85" swimtime="00:02:26.28" resultid="3294" lane="6" heatid="7061" entrytime="00:02:30.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.89" />
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                    <SPLIT distance="75" swimtime="00:00:50.09" />
                    <SPLIT distance="100" swimtime="00:01:08.19" />
                    <SPLIT distance="125" swimtime="00:01:26.88" />
                    <SPLIT distance="150" swimtime="00:01:46.34" />
                    <SPLIT distance="175" swimtime="00:02:06.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="391" reactiontime="+85" swimtime="00:00:29.08" resultid="3295" heatid="7344" entrytime="00:00:30.01">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="378" reactiontime="+91" swimtime="00:01:05.05" resultid="3292" heatid="6840" entrytime="00:01:06.01">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.89" />
                    <SPLIT distance="50" swimtime="00:00:31.47" />
                    <SPLIT distance="75" swimtime="00:00:48.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-11-18" firstname="Danuta" gender="F" lastname="Gojlik" nation="POL" athleteid="3296">
              <RESULTS>
                <RESULT eventid="1679" points="211" reactiontime="+92" swimtime="00:01:49.20" resultid="3299" lane="3" heatid="7297" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.77" />
                    <SPLIT distance="50" swimtime="00:00:52.23" />
                    <SPLIT distance="75" swimtime="00:01:20.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1409" points="207" reactiontime="+98" swimtime="00:03:57.00" resultid="3298" lane="2" heatid="7001" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.05" />
                    <SPLIT distance="50" swimtime="00:00:52.92" />
                    <SPLIT distance="75" swimtime="00:01:22.78" />
                    <SPLIT distance="100" swimtime="00:01:53.13" />
                    <SPLIT distance="125" swimtime="00:02:23.52" />
                    <SPLIT distance="150" swimtime="00:02:55.24" />
                    <SPLIT distance="175" swimtime="00:03:26.69" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="04 K-15" eventid="1222" reactiontime="+68" status="DSQ" swimtime="00:00:49.17" resultid="3297" lane="5" heatid="6850" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-03-21" firstname="Tomasz" gender="M" lastname="Wysocki" nation="POL" athleteid="3300">
              <RESULTS>
                <RESULT eventid="1109" points="484" reactiontime="+89" swimtime="00:01:05.13" resultid="3301" lane="2" heatid="6743" entrytime="00:01:07.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.80" />
                    <SPLIT distance="50" swimtime="00:00:28.70" />
                    <SPLIT distance="75" swimtime="00:00:49.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="403" reactiontime="+84" swimtime="00:02:34.22" resultid="3303" lane="8" heatid="6887" entrytime="00:02:33.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.55" />
                    <SPLIT distance="50" swimtime="00:00:35.13" />
                    <SPLIT distance="75" swimtime="00:00:54.35" />
                    <SPLIT distance="100" swimtime="00:01:14.53" />
                    <SPLIT distance="125" swimtime="00:01:34.71" />
                    <SPLIT distance="150" swimtime="00:01:55.12" />
                    <SPLIT distance="175" swimtime="00:02:15.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="567" reactiontime="+84" swimtime="00:00:25.70" resultid="3306" lane="6" heatid="7352" entrytime="00:00:26.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="611" reactiontime="+73" swimtime="00:00:28.83" resultid="3304" lane="2" heatid="7043" entrytime="00:00:28.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="597" reactiontime="+84" swimtime="00:00:27.26" resultid="3305" lane="2" heatid="7291" entrytime="00:00:29.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="491" reactiontime="+87" swimtime="00:00:34.44" resultid="3302" lane="6" heatid="6863" entrytime="00:00:36.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-08-29" firstname="Mirosław" gender="M" lastname="Radomski" nation="POL" athleteid="3307">
              <RESULTS>
                <RESULT eventid="1075" points="279" swimtime="00:11:41.50" resultid="3308" lane="3" heatid="6720" entrytime="00:12:00.00" />
                <RESULT eventid="1273" points="243" reactiontime="+113" swimtime="00:02:59.30" resultid="3309" lane="1" heatid="6872" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.37" />
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                    <SPLIT distance="75" swimtime="00:01:00.61" />
                    <SPLIT distance="100" swimtime="00:01:23.39" />
                    <SPLIT distance="125" swimtime="00:01:47.24" />
                    <SPLIT distance="150" swimtime="00:02:11.53" />
                    <SPLIT distance="175" swimtime="00:02:35.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="257" reactiontime="+110" swimtime="00:06:23.21" resultid="3312" lane="8" heatid="7361" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.75" />
                    <SPLIT distance="50" swimtime="00:00:39.69" />
                    <SPLIT distance="75" swimtime="00:01:03.01" />
                    <SPLIT distance="100" swimtime="00:01:27.26" />
                    <SPLIT distance="125" swimtime="00:01:56.73" />
                    <SPLIT distance="150" swimtime="00:03:18.64" />
                    <SPLIT distance="175" swimtime="00:02:52.14" />
                    <SPLIT distance="200" swimtime="00:04:11.26" />
                    <SPLIT distance="225" swimtime="00:03:45.25" />
                    <SPLIT distance="250" swimtime="00:05:04.30" />
                    <SPLIT distance="275" swimtime="00:04:37.67" />
                    <SPLIT distance="300" swimtime="00:05:47.35" />
                    <SPLIT distance="325" swimtime="00:06:05.83" />
                    <SPLIT distance="350" swimtime="00:06:23.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="303" reactiontime="+90" swimtime="00:03:09.67" resultid="3310" lane="6" heatid="7007" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.24" />
                    <SPLIT distance="50" swimtime="00:00:44.44" />
                    <SPLIT distance="75" swimtime="00:01:08.93" />
                    <SPLIT distance="100" swimtime="00:01:33.92" />
                    <SPLIT distance="125" swimtime="00:01:58.16" />
                    <SPLIT distance="150" swimtime="00:02:24.29" />
                    <SPLIT distance="175" swimtime="00:02:47.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" status="DNS" swimtime="00:00:00.00" resultid="3311" lane="3" heatid="7075" entrytime="00:03:10.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1177" status="DNS" swimtime="00:00:00.00" resultid="6670" lane="2" heatid="6807" />
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1177" status="DNS" swimtime="00:00:00.00" resultid="3313" lane="2" heatid="6809" entrytime="00:01:55.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3260" number="1" />
                    <RELAYPOSITION athleteid="3300" number="2" />
                    <RELAYPOSITION athleteid="3290" number="3" />
                    <RELAYPOSITION athleteid="3284" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="MKSZC" name="MKP Szczecin" nation="POL" region="ZAC">
          <CONTACT name="g" />
          <ATHLETES>
            <ATHLETE birthdate="1966-08-10" firstname="Małgorzata" gender="F" lastname="Serbin" nation="POL" athleteid="3318">
              <RESULTS>
                <RESULT comment="Rekord Polski " eventid="1713" points="457" reactiontime="+78" swimtime="00:01:16.28" resultid="3322" lane="6" heatid="7317" entrytime="00:01:16.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.58" />
                    <SPLIT distance="50" swimtime="00:00:37.48" />
                    <SPLIT distance="75" swimtime="00:00:56.93" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1547" points="517" reactiontime="+71" swimtime="00:02:22.99" resultid="3321" lane="3" heatid="7053" entrytime="00:02:25.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.79" />
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                    <SPLIT distance="75" swimtime="00:00:51.51" />
                    <SPLIT distance="100" swimtime="00:01:09.90" />
                    <SPLIT distance="125" swimtime="00:01:28.26" />
                    <SPLIT distance="150" swimtime="00:01:46.93" />
                    <SPLIT distance="175" swimtime="00:02:05.47" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1358" points="510" reactiontime="+74" swimtime="00:05:02.25" resultid="3320" lane="4" heatid="6898" entrytime="00:05:09.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.13" />
                    <SPLIT distance="50" swimtime="00:00:34.76" />
                    <SPLIT distance="75" swimtime="00:00:53.61" />
                    <SPLIT distance="100" swimtime="00:01:12.88" />
                    <SPLIT distance="125" swimtime="00:01:32.10" />
                    <SPLIT distance="150" swimtime="00:01:51.51" />
                    <SPLIT distance="175" swimtime="00:02:10.63" />
                    <SPLIT distance="200" swimtime="00:02:29.90" />
                    <SPLIT distance="225" swimtime="00:02:49.06" />
                    <SPLIT distance="250" swimtime="00:03:08.48" />
                    <SPLIT distance="275" swimtime="00:03:27.61" />
                    <SPLIT distance="300" swimtime="00:03:46.81" />
                    <SPLIT distance="325" swimtime="00:04:06.00" />
                    <SPLIT distance="350" swimtime="00:04:25.14" />
                    <SPLIT distance="375" swimtime="00:04:44.01" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1126" points="472" swimtime="00:20:09.90" resultid="3319" lane="3" heatid="6747" entrytime="00:20:30.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1935-09-01" firstname="Stefania" gender="F" lastname="Noetzel" nation="POL" athleteid="3323">
              <RESULTS>
                <RESULT comment="Rekord Polski " eventid="1679" points="109" swimtime="00:02:15.99" resultid="3326" lane="2" heatid="7296" entrytime="00:02:09.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:31.98" />
                    <SPLIT distance="50" swimtime="00:01:06.00" />
                    <SPLIT distance="75" swimtime="00:01:41.60" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1409" points="119" swimtime="00:04:44.75" resultid="3325" lane="1" heatid="6998" entrytime="00:04:42.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.54" />
                    <SPLIT distance="50" swimtime="00:01:07.23" />
                    <SPLIT distance="75" swimtime="00:01:43.35" />
                    <SPLIT distance="100" swimtime="00:02:19.21" />
                    <SPLIT distance="125" swimtime="00:02:55.98" />
                    <SPLIT distance="150" swimtime="00:03:33.09" />
                    <SPLIT distance="175" swimtime="00:04:09.73" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1222" points="105" swimtime="00:01:04.15" resultid="3324" lane="6" heatid="6848" entrytime="00:01:01.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:31.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-10-02" firstname="Piotr" gender="M" lastname="Kowalczyk" nation="POL" athleteid="3327">
              <RESULTS>
                <RESULT eventid="1075" points="406" swimtime="00:10:19.31" resultid="3328" lane="7" heatid="6722" entrytime="00:10:20.00" entrycourse="SCM" />
                <RESULT eventid="1375" points="438" reactiontime="+79" swimtime="00:04:49.67" resultid="3329" lane="6" heatid="6908" entrytime="00:04:54.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.00" />
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                    <SPLIT distance="75" swimtime="00:00:50.26" />
                    <SPLIT distance="100" swimtime="00:01:08.50" />
                    <SPLIT distance="125" swimtime="00:01:26.77" />
                    <SPLIT distance="150" swimtime="00:01:45.62" />
                    <SPLIT distance="175" swimtime="00:02:04.26" />
                    <SPLIT distance="200" swimtime="00:02:22.46" />
                    <SPLIT distance="225" swimtime="00:02:40.85" />
                    <SPLIT distance="250" swimtime="00:02:59.28" />
                    <SPLIT distance="275" swimtime="00:03:17.86" />
                    <SPLIT distance="300" swimtime="00:03:36.74" />
                    <SPLIT distance="325" swimtime="00:03:55.54" />
                    <SPLIT distance="350" swimtime="00:04:13.83" />
                    <SPLIT distance="375" swimtime="00:04:32.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="455" reactiontime="+76" swimtime="00:02:13.79" resultid="3330" lane="1" heatid="7064" entrytime="00:02:15.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.39" />
                    <SPLIT distance="50" swimtime="00:00:30.39" />
                    <SPLIT distance="75" swimtime="00:00:47.34" />
                    <SPLIT distance="100" swimtime="00:01:04.29" />
                    <SPLIT distance="125" swimtime="00:01:21.78" />
                    <SPLIT distance="150" swimtime="00:01:39.37" />
                    <SPLIT distance="175" swimtime="00:01:56.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-03-03" firstname="Agnieszka" gender="F" lastname="Kalska" nation="POL" athleteid="3331">
              <RESULTS>
                <RESULT eventid="1187" points="517" reactiontime="+74" swimtime="00:01:05.85" resultid="3332" lane="3" heatid="6828" entrytime="00:01:04.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.95" />
                    <SPLIT distance="50" swimtime="00:00:31.39" />
                    <SPLIT distance="75" swimtime="00:00:48.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="532" reactiontime="+73" swimtime="00:00:29.57" resultid="3334" lane="5" heatid="7335" entrytime="00:00:29.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="479" reactiontime="+77" swimtime="00:02:26.73" resultid="3333" lane="2" heatid="7053" entrytime="00:02:29.86">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.60" />
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                    <SPLIT distance="75" swimtime="00:00:51.84" />
                    <SPLIT distance="100" swimtime="00:01:10.49" />
                    <SPLIT distance="125" swimtime="00:01:29.20" />
                    <SPLIT distance="150" swimtime="00:01:48.61" />
                    <SPLIT distance="175" swimtime="00:02:07.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-01" firstname="Marcin" gender="M" lastname="Gargas" nation="POL" athleteid="4490">
              <RESULTS>
                <RESULT eventid="1564" points="172" reactiontime="+87" swimtime="00:03:04.78" resultid="4492" lane="2" heatid="7056" entrytime="00:03:03.91">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.42" />
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                    <SPLIT distance="75" swimtime="00:01:02.32" />
                    <SPLIT distance="100" swimtime="00:01:24.76" />
                    <SPLIT distance="125" swimtime="00:01:48.48" />
                    <SPLIT distance="150" swimtime="00:02:13.90" />
                    <SPLIT distance="175" swimtime="00:02:39.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="204" reactiontime="+93" swimtime="00:01:19.85" resultid="4491" lane="2" heatid="6832" entrytime="00:01:25.88">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.54" />
                    <SPLIT distance="50" swimtime="00:00:37.38" />
                    <SPLIT distance="75" swimtime="00:00:58.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOSZC" name="MOSRiR Szczecin" nation="POL" region="ZAC">
          <CONTACT name="Olszewski Bartosz" />
          <ATHLETES>
            <ATHLETE birthdate="1962-10-01" firstname="Aleksy" gender="M" lastname="Wierzchoń" nation="POL" athleteid="3336">
              <RESULTS>
                <RESULT eventid="1143" points="214" swimtime="00:24:20.37" resultid="3337" heatid="6751" entrytime="00:23:01.00" />
                <RESULT eventid="1411" points="286" reactiontime="+97" swimtime="00:03:13.38" resultid="3340" lane="4" heatid="7008" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.67" />
                    <SPLIT distance="50" swimtime="00:00:42.50" />
                    <SPLIT distance="75" swimtime="00:01:06.31" />
                    <SPLIT distance="100" swimtime="00:01:31.26" />
                    <SPLIT distance="125" swimtime="00:01:56.84" />
                    <SPLIT distance="150" swimtime="00:02:21.98" />
                    <SPLIT distance="175" swimtime="00:02:47.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="312" reactiontime="+101" swimtime="00:00:40.07" resultid="3338" lane="2" heatid="6858" entrytime="00:00:41.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" status="DNS" swimtime="00:00:00.00" resultid="3339" heatid="6908" entrytime="00:05:03.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="OMPOZ" name="One Man Team" nation="POL">
          <CONTACT email="gmo@o2.pl" name="MONCZAK, Grzegorz" />
          <ATHLETES>
            <ATHLETE birthdate="1973-05-25" firstname="Grzegorz" gender="M" lastname="Monczak" nation="POL" athleteid="3346">
              <RESULTS>
                <RESULT eventid="1375" points="473" reactiontime="+74" swimtime="00:04:42.31" resultid="3349" lane="5" heatid="6908" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.07" />
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                    <SPLIT distance="75" swimtime="00:00:49.76" />
                    <SPLIT distance="100" swimtime="00:01:07.57" />
                    <SPLIT distance="125" swimtime="00:01:25.58" />
                    <SPLIT distance="150" swimtime="00:01:43.75" />
                    <SPLIT distance="175" swimtime="00:02:01.81" />
                    <SPLIT distance="200" swimtime="00:02:19.93" />
                    <SPLIT distance="225" swimtime="00:02:38.21" />
                    <SPLIT distance="250" swimtime="00:02:56.61" />
                    <SPLIT distance="275" swimtime="00:03:15.09" />
                    <SPLIT distance="300" swimtime="00:03:33.49" />
                    <SPLIT distance="325" swimtime="00:03:51.68" />
                    <SPLIT distance="350" swimtime="00:04:09.67" />
                    <SPLIT distance="375" swimtime="00:04:26.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="464" swimtime="00:09:52.12" resultid="3347" lane="6" heatid="6722" entrytime="00:09:59.00" entrycourse="SCM" />
                <RESULT eventid="1798" points="393" reactiontime="+77" swimtime="00:05:32.76" resultid="3353" lane="7" heatid="7364" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.36" />
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                    <SPLIT distance="75" swimtime="00:00:53.84" />
                    <SPLIT distance="100" swimtime="00:01:14.22" />
                    <SPLIT distance="125" swimtime="00:01:36.57" />
                    <SPLIT distance="150" swimtime="00:01:58.21" />
                    <SPLIT distance="175" swimtime="00:02:20.15" />
                    <SPLIT distance="200" swimtime="00:02:41.91" />
                    <SPLIT distance="225" swimtime="00:03:06.52" />
                    <SPLIT distance="250" swimtime="00:03:30.61" />
                    <SPLIT distance="275" swimtime="00:03:54.65" />
                    <SPLIT distance="300" swimtime="00:04:18.89" />
                    <SPLIT distance="325" swimtime="00:04:38.20" />
                    <SPLIT distance="350" swimtime="00:04:56.87" />
                    <SPLIT distance="375" swimtime="00:05:15.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="413" reactiontime="+73" swimtime="00:02:33.27" resultid="3351" lane="4" heatid="7077" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.59" />
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                    <SPLIT distance="75" swimtime="00:00:52.82" />
                    <SPLIT distance="100" swimtime="00:01:13.21" />
                    <SPLIT distance="125" swimtime="00:01:35.63" />
                    <SPLIT distance="150" swimtime="00:01:58.45" />
                    <SPLIT distance="175" swimtime="00:02:16.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="505" reactiontime="+73" swimtime="00:02:09.29" resultid="3350" lane="3" heatid="7064" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.47" />
                    <SPLIT distance="50" swimtime="00:00:30.44" />
                    <SPLIT distance="75" swimtime="00:00:46.89" />
                    <SPLIT distance="100" swimtime="00:01:03.42" />
                    <SPLIT distance="125" swimtime="00:01:20.02" />
                    <SPLIT distance="150" swimtime="00:01:36.58" />
                    <SPLIT distance="175" swimtime="00:01:52.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="491" reactiontime="+71" swimtime="00:00:59.61" resultid="3348" heatid="6844" entrytime="00:00:59.99">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.84" />
                    <SPLIT distance="50" swimtime="00:00:29.06" />
                    <SPLIT distance="75" swimtime="00:00:44.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" status="DNS" swimtime="00:00:00.00" resultid="3352" lane="7" heatid="7309" entrytime="00:01:22.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KONST" name="Konstancin-Jeziorna" nation="POL">
          <CONTACT name="Obiedziński" />
          <ATHLETES>
            <ATHLETE birthdate="1969-04-11" firstname="Paweł" gender="M" lastname="Obiedziński" nation="POL" athleteid="3355">
              <RESULTS>
                <RESULT eventid="1411" points="346" reactiontime="+80" swimtime="00:03:01.53" resultid="3358" lane="8" heatid="7010" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.12" />
                    <SPLIT distance="50" swimtime="00:00:39.69" />
                    <SPLIT distance="75" swimtime="00:01:01.93" />
                    <SPLIT distance="100" swimtime="00:01:25.02" />
                    <SPLIT distance="125" swimtime="00:01:49.03" />
                    <SPLIT distance="150" swimtime="00:02:13.55" />
                    <SPLIT distance="175" swimtime="00:02:37.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="424" reactiontime="+74" swimtime="00:02:17.04" resultid="3359" lane="5" heatid="7063" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.26" />
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                    <SPLIT distance="75" swimtime="00:00:46.62" />
                    <SPLIT distance="100" swimtime="00:01:04.04" />
                    <SPLIT distance="125" swimtime="00:01:21.44" />
                    <SPLIT distance="150" swimtime="00:01:39.93" />
                    <SPLIT distance="175" swimtime="00:01:58.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="455" reactiontime="+71" swimtime="00:01:01.16" resultid="3356" lane="1" heatid="6842" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.79" />
                    <SPLIT distance="50" swimtime="00:00:29.06" />
                    <SPLIT distance="75" swimtime="00:00:45.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="429" reactiontime="+71" swimtime="00:00:30.43" resultid="3360" lane="3" heatid="7289" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="495" reactiontime="+73" swimtime="00:00:26.89" resultid="3361" lane="3" heatid="7348" entrytime="00:00:27.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="397" reactiontime="+70" swimtime="00:00:36.98" resultid="3357" lane="6" heatid="6862" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MTLUB" name="MTP Lublinianka" nation="POL" region="LBL">
          <CONTACT city="Lublin" email="jerzy.paleolog@up.lublin.pl" internet="http://www.lublinianka.website.pl/index.html" name="Jerzy Demetraki_paleolog" phone="+48602 725175" state="LUBEL" street="Doswiadczalna 50C/5" zip="20-280" />
          <ATHLETES>
            <ATHLETE birthdate="1955-03-07" firstname="Jerzy" gender="M" lastname="Demetraki-Paleolog" nation="POL" athleteid="3363">
              <RESULTS>
                <RESULT eventid="1798" points="206" reactiontime="+107" swimtime="00:06:52.84" resultid="3368" lane="4" heatid="7360" entrytime="00:06:59.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.45" />
                    <SPLIT distance="50" swimtime="00:00:46.71" />
                    <SPLIT distance="75" swimtime="00:01:13.12" />
                    <SPLIT distance="100" swimtime="00:01:41.64" />
                    <SPLIT distance="125" swimtime="00:02:09.31" />
                    <SPLIT distance="150" swimtime="00:02:36.99" />
                    <SPLIT distance="175" swimtime="00:03:04.74" />
                    <SPLIT distance="200" swimtime="00:03:31.19" />
                    <SPLIT distance="225" swimtime="00:03:59.36" />
                    <SPLIT distance="250" swimtime="00:04:27.12" />
                    <SPLIT distance="275" swimtime="00:04:56.02" />
                    <SPLIT distance="300" swimtime="00:05:26.23" />
                    <SPLIT distance="325" swimtime="00:05:49.80" />
                    <SPLIT distance="350" swimtime="00:06:12.02" />
                    <SPLIT distance="375" swimtime="00:06:32.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="167" reactiontime="+111" swimtime="00:03:23.17" resultid="3365" lane="2" heatid="6871" entrytime="00:03:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.49" />
                    <SPLIT distance="50" swimtime="00:00:47.48" />
                    <SPLIT distance="75" swimtime="00:01:15.06" />
                    <SPLIT distance="100" swimtime="00:01:42.64" />
                    <SPLIT distance="125" swimtime="00:02:08.29" />
                    <SPLIT distance="150" swimtime="00:02:33.45" />
                    <SPLIT distance="175" swimtime="00:02:58.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="222" swimtime="00:12:37.30" resultid="3364" heatid="6721" entrytime="00:11:19.20" entrycourse="SCM" />
                <RESULT eventid="1462" points="189" reactiontime="+109" swimtime="00:01:27.76" resultid="3367" lane="8" heatid="7018" entrytime="00:01:28.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.74" />
                    <SPLIT distance="50" swimtime="00:00:41.63" />
                    <SPLIT distance="75" swimtime="00:01:04.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="237" reactiontime="+132" swimtime="00:05:55.58" resultid="3366" lane="8" heatid="6904" entrytime="00:05:54.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.48" />
                    <SPLIT distance="50" swimtime="00:00:41.24" />
                    <SPLIT distance="75" swimtime="00:01:03.42" />
                    <SPLIT distance="100" swimtime="00:01:26.79" />
                    <SPLIT distance="125" swimtime="00:01:48.81" />
                    <SPLIT distance="150" swimtime="00:02:10.96" />
                    <SPLIT distance="175" swimtime="00:02:34.20" />
                    <SPLIT distance="200" swimtime="00:02:57.18" />
                    <SPLIT distance="225" swimtime="00:03:19.56" />
                    <SPLIT distance="250" swimtime="00:03:41.13" />
                    <SPLIT distance="275" swimtime="00:04:03.71" />
                    <SPLIT distance="300" swimtime="00:04:26.29" />
                    <SPLIT distance="325" swimtime="00:04:48.28" />
                    <SPLIT distance="350" swimtime="00:05:10.90" />
                    <SPLIT distance="375" swimtime="00:05:33.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SUWAR" name="Sródmiejski U.K.S.Polna Warszawa" nation="POL">
          <CONTACT city="Warszawa" name="Przybylski Piotr" phone="501-704-665" street="Polna7a" zip="00-625" />
          <ATHLETES>
            <ATHLETE birthdate="1975-01-05" firstname="Bartłomiej" gender="M" lastname="Pawłowski" nation="POL" athleteid="3370">
              <RESULTS>
                <RESULT eventid="1239" points="439" reactiontime="+84" swimtime="00:00:35.74" resultid="3373" lane="8" heatid="6860" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="456" reactiontime="+80" swimtime="00:00:27.63" resultid="3374" lane="8" heatid="7339" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="323" reactiontime="+84" swimtime="00:01:14.51" resultid="3371" lane="7" heatid="6738" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.65" />
                    <SPLIT distance="50" swimtime="00:00:34.76" />
                    <SPLIT distance="75" swimtime="00:00:56.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="3372" lane="4" heatid="6836" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="NZWAW" name="K.S. niezrzeszeni.pl" nation="POL" region="WA">
          <CONTACT city="Warszawa" email="niezrzeszenipl@gmail.com" internet="niezrzeszeni.pl" name="Wawer Matylda Katarzyna" phone="501701359" />
          <ATHLETES>
            <ATHLETE birthdate="1954-04-08" firstname="Wojciech" gender="M" lastname="Staruch" nation="POL" athleteid="3384">
              <RESULTS>
                <RESULT eventid="1239" points="330" reactiontime="+89" swimtime="00:00:39.33" resultid="3386" lane="8" heatid="6859" entrytime="00:00:40.17">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="262" reactiontime="+85" swimtime="00:01:31.96" resultid="3390" lane="5" heatid="7306" entrytime="00:01:31.12">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.58" />
                    <SPLIT distance="50" swimtime="00:00:42.82" />
                    <SPLIT distance="75" swimtime="00:01:07.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="210" reactiontime="+89" swimtime="00:01:26.05" resultid="3385" lane="4" heatid="6734" entrytime="00:01:27.88">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.60" />
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                    <SPLIT distance="75" swimtime="00:01:05.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="149" reactiontime="+94" swimtime="00:03:14.04" resultid="3389" heatid="7057" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.56" />
                    <SPLIT distance="50" swimtime="00:00:41.79" />
                    <SPLIT distance="75" swimtime="00:01:04.76" />
                    <SPLIT distance="100" swimtime="00:01:29.36" />
                    <SPLIT distance="125" swimtime="00:01:55.03" />
                    <SPLIT distance="150" swimtime="00:02:21.27" />
                    <SPLIT distance="175" swimtime="00:02:48.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="213" reactiontime="+102" swimtime="00:03:33.43" resultid="3388" lane="5" heatid="7006" entrytime="00:03:29.01">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.02" />
                    <SPLIT distance="50" swimtime="00:00:46.49" />
                    <SPLIT distance="75" swimtime="00:01:12.93" />
                    <SPLIT distance="100" swimtime="00:01:40.50" />
                    <SPLIT distance="125" swimtime="00:02:09.00" />
                    <SPLIT distance="150" swimtime="00:02:37.83" />
                    <SPLIT distance="175" swimtime="00:03:06.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="273" reactiontime="+86" swimtime="00:00:32.79" resultid="3391" lane="7" heatid="7341" entrytime="00:00:32.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="148" reactiontime="+103" swimtime="00:06:55.45" resultid="3387" heatid="6901" entrytime="00:07:04.99">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.00" />
                    <SPLIT distance="50" swimtime="00:00:43.04" />
                    <SPLIT distance="75" swimtime="00:01:06.54" />
                    <SPLIT distance="100" swimtime="00:01:31.29" />
                    <SPLIT distance="125" swimtime="00:01:57.22" />
                    <SPLIT distance="150" swimtime="00:02:23.37" />
                    <SPLIT distance="175" swimtime="00:02:50.11" />
                    <SPLIT distance="200" swimtime="00:03:17.08" />
                    <SPLIT distance="225" swimtime="00:03:43.90" />
                    <SPLIT distance="250" swimtime="00:04:11.58" />
                    <SPLIT distance="275" swimtime="00:04:38.96" />
                    <SPLIT distance="300" swimtime="00:05:06.65" />
                    <SPLIT distance="325" swimtime="00:05:34.50" />
                    <SPLIT distance="350" swimtime="00:06:03.03" />
                    <SPLIT distance="375" swimtime="00:06:30.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-12-27" firstname="Wojciech" gender="M" lastname="Korpetta" nation="POL" athleteid="3392">
              <RESULTS>
                <RESULT eventid="1307" points="191" reactiontime="+66" swimtime="00:03:17.54" resultid="3395" lane="2" heatid="6883" entrytime="00:03:25.04">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.17" />
                    <SPLIT distance="50" swimtime="00:02:30.29" />
                    <SPLIT distance="75" swimtime="00:01:12.40" />
                    <SPLIT distance="100" swimtime="00:03:17.54" />
                    <SPLIT distance="125" swimtime="00:02:04.06" />
                    <SPLIT distance="175" swimtime="00:02:55.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="147" reactiontime="+118" swimtime="00:03:36.14" resultid="3397" lane="5" heatid="7073" entrytime="00:03:35.67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.03" />
                    <SPLIT distance="50" swimtime="00:00:49.68" />
                    <SPLIT distance="75" swimtime="00:01:18.05" />
                    <SPLIT distance="100" swimtime="00:01:44.19" />
                    <SPLIT distance="125" swimtime="00:02:16.02" />
                    <SPLIT distance="150" swimtime="00:02:47.42" />
                    <SPLIT distance="175" swimtime="00:03:12.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="224" reactiontime="+64" swimtime="00:00:40.26" resultid="3396" lane="5" heatid="7036" entrytime="00:00:41.26">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="203" reactiontime="+60" swimtime="00:01:29.30" resultid="3398" lane="3" heatid="7321" entrytime="00:01:32.05">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.93" />
                    <SPLIT distance="50" swimtime="00:00:43.34" />
                    <SPLIT distance="75" swimtime="00:01:06.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="215" reactiontime="+102" swimtime="00:00:45.31" resultid="3394" lane="6" heatid="6856" entrytime="00:00:45.16">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="172" reactiontime="+121" swimtime="00:01:31.94" resultid="3393" lane="6" heatid="6733" entrytime="00:01:32.31">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.90" />
                    <SPLIT distance="50" swimtime="00:00:44.12" />
                    <SPLIT distance="75" swimtime="00:01:10.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-14" firstname="Andrzej" gender="M" lastname="Miński" nation="POL" athleteid="3400">
              <RESULTS>
                <RESULT eventid="1143" points="191" swimtime="00:25:16.85" resultid="3401" lane="3" heatid="6749" entrytime="00:25:45.38" />
                <RESULT eventid="1375" points="184" reactiontime="+108" swimtime="00:06:26.36" resultid="3403" lane="1" heatid="6902" entrytime="00:06:17.72">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.80" />
                    <SPLIT distance="50" swimtime="00:00:42.22" />
                    <SPLIT distance="75" swimtime="00:01:05.57" />
                    <SPLIT distance="100" swimtime="00:01:29.93" />
                    <SPLIT distance="125" swimtime="00:01:54.92" />
                    <SPLIT distance="150" swimtime="00:02:20.14" />
                    <SPLIT distance="175" swimtime="00:02:45.43" />
                    <SPLIT distance="200" swimtime="00:03:10.67" />
                    <SPLIT distance="225" swimtime="00:03:36.17" />
                    <SPLIT distance="250" swimtime="00:04:00.88" />
                    <SPLIT distance="275" swimtime="00:04:26.09" />
                    <SPLIT distance="300" swimtime="00:04:50.91" />
                    <SPLIT distance="325" swimtime="00:05:15.70" />
                    <SPLIT distance="350" swimtime="00:05:40.23" />
                    <SPLIT distance="375" swimtime="00:06:03.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="214" reactiontime="+110" swimtime="00:01:38.40" resultid="3406" lane="1" heatid="7305" entrytime="00:01:38.17">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.88" />
                    <SPLIT distance="50" swimtime="00:00:46.66" />
                    <SPLIT distance="75" swimtime="00:01:12.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="186" reactiontime="+110" swimtime="00:03:43.36" resultid="3404" lane="2" heatid="7006" entrytime="00:03:29.71">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.50" />
                    <SPLIT distance="50" swimtime="00:00:51.78" />
                    <SPLIT distance="75" swimtime="00:01:19.80" />
                    <SPLIT distance="100" swimtime="00:01:48.00" />
                    <SPLIT distance="125" swimtime="00:02:16.85" />
                    <SPLIT distance="150" swimtime="00:02:45.94" />
                    <SPLIT distance="175" swimtime="00:03:15.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="135" reactiontime="+116" swimtime="00:07:54.99" resultid="3407" lane="3" heatid="7358">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.06" />
                    <SPLIT distance="50" swimtime="00:00:54.78" />
                    <SPLIT distance="75" swimtime="00:01:25.17" />
                    <SPLIT distance="100" swimtime="00:01:56.88" />
                    <SPLIT distance="125" swimtime="00:02:33.61" />
                    <SPLIT distance="150" swimtime="00:03:10.36" />
                    <SPLIT distance="175" swimtime="00:03:45.45" />
                    <SPLIT distance="200" swimtime="00:04:21.65" />
                    <SPLIT distance="225" swimtime="00:04:50.95" />
                    <SPLIT distance="250" swimtime="00:05:20.69" />
                    <SPLIT distance="275" swimtime="00:05:50.50" />
                    <SPLIT distance="300" swimtime="00:06:20.67" />
                    <SPLIT distance="325" swimtime="00:06:44.57" />
                    <SPLIT distance="350" swimtime="00:07:08.74" />
                    <SPLIT distance="375" swimtime="00:07:33.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="186" reactiontime="+106" swimtime="00:01:22.33" resultid="3402" lane="7" heatid="6833" entrytime="00:01:20.98">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.26" />
                    <SPLIT distance="50" swimtime="00:00:38.60" />
                    <SPLIT distance="75" swimtime="00:01:00.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="3405" lane="1" heatid="7057" entrytime="00:02:59.19" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-07-16" firstname="Matylda Katarzyna" gender="F" lastname="Wawer" nation="POL" athleteid="3408">
              <RESULTS>
                <RESULT eventid="1547" points="189" reactiontime="+92" swimtime="00:03:19.94" resultid="3412" lane="2" heatid="7050" entrytime="00:03:15.89">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.48" />
                    <SPLIT distance="50" swimtime="00:00:45.56" />
                    <SPLIT distance="75" swimtime="00:01:10.19" />
                    <SPLIT distance="100" swimtime="00:01:36.12" />
                    <SPLIT distance="125" swimtime="00:02:02.38" />
                    <SPLIT distance="150" swimtime="00:02:29.30" />
                    <SPLIT distance="175" swimtime="00:02:56.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="216" reactiontime="+84" swimtime="00:00:42.39" resultid="3413" lane="3" heatid="7277" entrytime="00:00:43.29">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1445" points="135" reactiontime="+91" swimtime="00:01:50.23" resultid="3411" lane="4" heatid="7012" entrytime="00:01:52.47">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.78" />
                    <SPLIT distance="50" swimtime="00:00:51.79" />
                    <SPLIT distance="75" swimtime="00:01:22.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="254" reactiontime="+89" swimtime="00:01:23.44" resultid="3409" heatid="6825" entrytime="00:01:23.37">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.34" />
                    <SPLIT distance="50" swimtime="00:00:40.22" />
                    <SPLIT distance="75" swimtime="00:01:02.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="293" reactiontime="+88" swimtime="00:00:36.06" resultid="3414" lane="3" heatid="7331" entrytime="00:00:36.33">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOSTA" name="MOTYL SENIOR MOSiR Stalowa Wola" nation="POL" region="PDK">
          <CONTACT city="Stalowa Wola" email="lorkowska@wp.pl" name="Chmielewski Andrzej" phone="15-8422562 wew.45" state="PODK" street="Hutnicza 15" zip="37-450-" />
          <ATHLETES>
            <ATHLETE birthdate="1975-03-19" firstname="Robert" gender="M" lastname="Baran" nation="POL" athleteid="3416">
              <RESULTS>
                <RESULT eventid="1730" points="501" reactiontime="+70" swimtime="00:01:06.13" resultid="3422" lane="4" heatid="7325" entrytime="00:01:07.77">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.38" />
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                    <SPLIT distance="75" swimtime="00:00:49.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="477" reactiontime="+75" swimtime="00:02:25.82" resultid="3419" lane="7" heatid="6887" entrytime="00:02:29.57">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.42" />
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                    <SPLIT distance="75" swimtime="00:00:52.23" />
                    <SPLIT distance="100" swimtime="00:01:11.05" />
                    <SPLIT distance="125" swimtime="00:01:29.50" />
                    <SPLIT distance="150" swimtime="00:01:48.57" />
                    <SPLIT distance="175" swimtime="00:02:07.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="519" reactiontime="+70" swimtime="00:00:30.43" resultid="3420" heatid="7042" entrytime="00:00:30.92">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="520" reactiontime="+86" swimtime="00:00:58.50" resultid="3418" lane="1" heatid="6843" entrytime="00:01:00.35">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.26" />
                    <SPLIT distance="50" swimtime="00:00:28.00" />
                    <SPLIT distance="75" swimtime="00:00:43.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="517" reactiontime="+84" swimtime="00:00:26.50" resultid="3423" lane="1" heatid="7350" entrytime="00:00:27.42">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="383" reactiontime="+87" swimtime="00:02:37.21" resultid="3421" heatid="7079" entrytime="00:02:34.34">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.38" />
                    <SPLIT distance="50" swimtime="00:00:31.92" />
                    <SPLIT distance="75" swimtime="00:00:50.89" />
                    <SPLIT distance="100" swimtime="00:01:09.09" />
                    <SPLIT distance="125" swimtime="00:01:33.69" />
                    <SPLIT distance="150" swimtime="00:01:58.69" />
                    <SPLIT distance="175" swimtime="00:02:18.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="425" reactiontime="+96" swimtime="00:01:08.02" resultid="3417" lane="3" heatid="6742" entrytime="00:01:09.08">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.21" />
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                    <SPLIT distance="75" swimtime="00:00:52.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-14" firstname="Arkadiusz" gender="M" lastname="Berwecki" nation="POL" athleteid="3424">
              <RESULTS>
                <RESULT eventid="1109" points="492" swimtime="00:01:04.78" resultid="3425" lane="1" heatid="6745" entrytime="00:01:03.51" />
                <RESULT eventid="1239" points="534" reactiontime="+72" swimtime="00:00:33.50" resultid="3427" heatid="6865" entrytime="00:00:34.01">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="565" reactiontime="+72" swimtime="00:00:56.88" resultid="3426" heatid="6846" entrytime="00:00:57.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.75" />
                    <SPLIT distance="50" swimtime="00:00:27.10" />
                    <SPLIT distance="75" swimtime="00:00:41.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="565" reactiontime="+70" swimtime="00:00:25.74" resultid="3431" lane="7" heatid="7353" entrytime="00:00:26.01">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="571" reactiontime="+70" swimtime="00:01:00.75" resultid="3428" lane="6" heatid="7023" entrytime="00:01:00.11">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.07" />
                    <SPLIT distance="50" swimtime="00:00:28.39" />
                    <SPLIT distance="75" swimtime="00:00:44.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="544" reactiontime="+74" swimtime="00:02:06.09" resultid="3429" lane="7" heatid="7066" entrytime="00:02:04.51">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.57" />
                    <SPLIT distance="50" swimtime="00:00:28.64" />
                    <SPLIT distance="75" swimtime="00:00:44.20" />
                    <SPLIT distance="100" swimtime="00:01:00.31" />
                    <SPLIT distance="125" swimtime="00:01:16.56" />
                    <SPLIT distance="150" swimtime="00:01:33.24" />
                    <SPLIT distance="175" swimtime="00:01:49.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="598" reactiontime="+69" swimtime="00:00:27.25" resultid="3430" lane="7" heatid="7294" entrytime="00:00:26.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-15" firstname="Paweł" gender="M" lastname="Cieśliński" nation="POL" athleteid="3432">
              <RESULTS>
                <RESULT eventid="1273" points="216" reactiontime="+94" swimtime="00:03:06.45" resultid="3435" lane="6" heatid="6872" entrytime="00:03:10.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.03" />
                    <SPLIT distance="50" swimtime="00:00:43.08" />
                    <SPLIT distance="75" swimtime="00:01:07.30" />
                    <SPLIT distance="100" swimtime="00:01:31.02" />
                    <SPLIT distance="125" swimtime="00:01:55.91" />
                    <SPLIT distance="150" swimtime="00:02:20.21" />
                    <SPLIT distance="175" swimtime="00:02:44.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="330" reactiontime="+99" swimtime="00:03:04.45" resultid="3436" lane="6" heatid="7008" entrytime="00:03:10.11">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.66" />
                    <SPLIT distance="50" swimtime="00:00:42.54" />
                    <SPLIT distance="75" swimtime="00:01:05.85" />
                    <SPLIT distance="100" swimtime="00:01:29.83" />
                    <SPLIT distance="125" swimtime="00:01:53.91" />
                    <SPLIT distance="150" swimtime="00:02:18.26" />
                    <SPLIT distance="175" swimtime="00:02:41.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="249" reactiontime="+91" swimtime="00:06:27.09" resultid="3439" lane="4" heatid="7361" entrytime="00:06:30.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.05" />
                    <SPLIT distance="50" swimtime="00:00:44.13" />
                    <SPLIT distance="75" swimtime="00:01:09.45" />
                    <SPLIT distance="100" swimtime="00:01:35.53" />
                    <SPLIT distance="125" swimtime="00:02:01.11" />
                    <SPLIT distance="150" swimtime="00:02:25.67" />
                    <SPLIT distance="175" swimtime="00:02:50.70" />
                    <SPLIT distance="200" swimtime="00:03:15.80" />
                    <SPLIT distance="225" swimtime="00:03:42.30" />
                    <SPLIT distance="250" swimtime="00:04:07.24" />
                    <SPLIT distance="275" swimtime="00:04:32.66" />
                    <SPLIT distance="300" swimtime="00:04:58.95" />
                    <SPLIT distance="325" swimtime="00:05:22.01" />
                    <SPLIT distance="350" swimtime="00:05:44.82" />
                    <SPLIT distance="375" swimtime="00:06:07.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="365" reactiontime="+77" swimtime="00:01:22.42" resultid="3438" lane="6" heatid="7308" entrytime="00:01:25.11">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.26" />
                    <SPLIT distance="50" swimtime="00:00:39.32" />
                    <SPLIT distance="75" swimtime="00:01:01.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="395" reactiontime="+70" swimtime="00:00:37.03" resultid="3434" lane="3" heatid="6860" entrytime="00:00:38.05">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="277" reactiontime="+80" swimtime="00:01:18.46" resultid="3433" lane="3" heatid="6736" entrytime="00:01:20.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.89" />
                    <SPLIT distance="50" swimtime="00:00:37.49" />
                    <SPLIT distance="75" swimtime="00:00:59.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" status="DNS" swimtime="00:00:00.00" resultid="3437" lane="2" heatid="7075" entrytime="00:03:10.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-02-07" firstname="Paweł" gender="M" lastname="Ciurko" nation="POL" athleteid="3440">
              <RESULTS>
                <RESULT eventid="1798" points="289" reactiontime="+87" swimtime="00:06:08.71" resultid="3447" lane="2" heatid="7363" entrytime="00:06:05.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.36" />
                    <SPLIT distance="50" swimtime="00:00:41.11" />
                    <SPLIT distance="75" swimtime="00:01:05.15" />
                    <SPLIT distance="100" swimtime="00:01:30.49" />
                    <SPLIT distance="125" swimtime="00:01:57.06" />
                    <SPLIT distance="150" swimtime="00:02:22.17" />
                    <SPLIT distance="175" swimtime="00:02:46.81" />
                    <SPLIT distance="200" swimtime="00:03:11.70" />
                    <SPLIT distance="225" swimtime="00:03:35.54" />
                    <SPLIT distance="250" swimtime="00:03:58.90" />
                    <SPLIT distance="275" swimtime="00:04:22.08" />
                    <SPLIT distance="300" swimtime="00:04:45.43" />
                    <SPLIT distance="325" swimtime="00:05:06.67" />
                    <SPLIT distance="350" swimtime="00:05:28.00" />
                    <SPLIT distance="375" swimtime="00:05:48.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="224" reactiontime="+89" swimtime="00:03:04.22" resultid="3443" lane="8" heatid="6873" entrytime="00:03:01.11">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.92" />
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                    <SPLIT distance="75" swimtime="00:00:58.25" />
                    <SPLIT distance="100" swimtime="00:01:21.08" />
                    <SPLIT distance="125" swimtime="00:01:45.02" />
                    <SPLIT distance="150" swimtime="00:02:11.65" />
                    <SPLIT distance="175" swimtime="00:02:37.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="425" reactiontime="+85" swimtime="00:01:18.32" resultid="3446" lane="8" heatid="7310" entrytime="00:01:18.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.01" />
                    <SPLIT distance="50" swimtime="00:00:37.16" />
                    <SPLIT distance="75" swimtime="00:00:57.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="379" reactiontime="+89" swimtime="00:02:56.19" resultid="3444" heatid="7008" entrytime="00:03:10.89">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.13" />
                    <SPLIT distance="50" swimtime="00:00:40.35" />
                    <SPLIT distance="75" swimtime="00:01:02.25" />
                    <SPLIT distance="100" swimtime="00:01:24.76" />
                    <SPLIT distance="125" swimtime="00:01:48.39" />
                    <SPLIT distance="150" swimtime="00:02:11.11" />
                    <SPLIT distance="175" swimtime="00:02:34.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="303" reactiontime="+88" swimtime="00:02:50.00" resultid="3445" lane="4" heatid="7076" entrytime="00:02:59.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.20" />
                    <SPLIT distance="50" swimtime="00:00:36.25" />
                    <SPLIT distance="75" swimtime="00:01:01.14" />
                    <SPLIT distance="100" swimtime="00:01:25.12" />
                    <SPLIT distance="125" swimtime="00:01:46.88" />
                    <SPLIT distance="150" swimtime="00:02:09.69" />
                    <SPLIT distance="175" swimtime="00:02:30.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="347" reactiontime="+79" swimtime="00:01:06.91" resultid="3442" lane="3" heatid="6836" entrytime="00:01:10.03">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.42" />
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                    <SPLIT distance="75" swimtime="00:00:49.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="283" reactiontime="+90" swimtime="00:01:17.90" resultid="3441" lane="2" heatid="6737" entrytime="00:01:19.11">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.75" />
                    <SPLIT distance="50" swimtime="00:00:38.31" />
                    <SPLIT distance="75" swimtime="00:00:58.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-08-09" firstname="Włodzimierz" gender="M" lastname="Jarzyna" nation="POL" athleteid="3448">
              <RESULTS>
                <RESULT eventid="1598" points="186" reactiontime="+97" swimtime="00:03:19.96" resultid="3453" heatid="7075" entrytime="00:03:17.18">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.23" />
                    <SPLIT distance="50" swimtime="00:00:46.05" />
                    <SPLIT distance="75" swimtime="00:01:12.31" />
                    <SPLIT distance="100" swimtime="00:01:38.98" />
                    <SPLIT distance="125" swimtime="00:02:08.22" />
                    <SPLIT distance="150" swimtime="00:02:36.65" />
                    <SPLIT distance="175" swimtime="00:03:00.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="188" reactiontime="+92" swimtime="00:07:05.32" resultid="3455" lane="6" heatid="7359" entrytime="00:07:37.42">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.97" />
                    <SPLIT distance="50" swimtime="00:00:47.79" />
                    <SPLIT distance="75" swimtime="00:01:15.85" />
                    <SPLIT distance="100" swimtime="00:01:43.17" />
                    <SPLIT distance="125" swimtime="00:02:12.01" />
                    <SPLIT distance="150" swimtime="00:02:40.17" />
                    <SPLIT distance="175" swimtime="00:03:07.39" />
                    <SPLIT distance="200" swimtime="00:03:33.74" />
                    <SPLIT distance="225" swimtime="00:04:03.34" />
                    <SPLIT distance="250" swimtime="00:04:33.26" />
                    <SPLIT distance="275" swimtime="00:05:02.81" />
                    <SPLIT distance="300" swimtime="00:05:32.64" />
                    <SPLIT distance="325" swimtime="00:05:57.38" />
                    <SPLIT distance="350" swimtime="00:06:21.12" />
                    <SPLIT distance="375" swimtime="00:06:44.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="177" reactiontime="+92" swimtime="00:03:22.61" resultid="3450" lane="4" heatid="6882" entrytime="00:03:41.41">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.33" />
                    <SPLIT distance="50" swimtime="00:00:47.83" />
                    <SPLIT distance="75" swimtime="00:01:13.05" />
                    <SPLIT distance="100" swimtime="00:01:39.69" />
                    <SPLIT distance="125" swimtime="00:02:06.79" />
                    <SPLIT distance="150" swimtime="00:02:34.17" />
                    <SPLIT distance="175" swimtime="00:02:59.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="197" reactiontime="+96" swimtime="00:06:17.68" resultid="3451" lane="2" heatid="6901" entrytime="00:06:38.81">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.07" />
                    <SPLIT distance="50" swimtime="00:00:40.77" />
                    <SPLIT distance="75" swimtime="00:01:03.42" />
                    <SPLIT distance="100" swimtime="00:01:26.62" />
                    <SPLIT distance="125" swimtime="00:01:50.29" />
                    <SPLIT distance="150" swimtime="00:02:14.54" />
                    <SPLIT distance="175" swimtime="00:02:38.96" />
                    <SPLIT distance="200" swimtime="00:03:03.44" />
                    <SPLIT distance="225" swimtime="00:03:27.93" />
                    <SPLIT distance="250" swimtime="00:03:52.84" />
                    <SPLIT distance="275" swimtime="00:04:17.41" />
                    <SPLIT distance="300" swimtime="00:04:41.47" />
                    <SPLIT distance="325" swimtime="00:05:04.82" />
                    <SPLIT distance="350" swimtime="00:05:26.30" />
                    <SPLIT distance="375" swimtime="00:05:55.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="176" swimtime="00:13:37.58" resultid="3449" lane="8" heatid="6718" entrytime="00:14:07.27" />
                <RESULT eventid="1411" points="208" reactiontime="+91" swimtime="00:03:35.01" resultid="3452" lane="3" heatid="7004" entrytime="00:03:49.17">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.25" />
                    <SPLIT distance="50" swimtime="00:00:48.53" />
                    <SPLIT distance="75" swimtime="00:01:15.48" />
                    <SPLIT distance="100" swimtime="00:01:43.19" />
                    <SPLIT distance="125" swimtime="00:02:12.02" />
                    <SPLIT distance="150" swimtime="00:02:40.45" />
                    <SPLIT distance="175" swimtime="00:03:08.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="196" reactiontime="+76" swimtime="00:01:30.40" resultid="3454" lane="4" heatid="7320" entrytime="00:01:41.38">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.49" />
                    <SPLIT distance="50" swimtime="00:00:45.82" />
                    <SPLIT distance="75" swimtime="00:01:09.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-18" firstname="Waldemar" gender="M" lastname="Kalbarczyk" nation="POL" athleteid="3456">
              <RESULTS>
                <RESULT eventid="1273" points="192" reactiontime="+91" swimtime="00:03:13.91" resultid="3459" lane="5" heatid="6872" entrytime="00:03:08.25">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.60" />
                    <SPLIT distance="50" swimtime="00:00:42.11" />
                    <SPLIT distance="75" swimtime="00:01:07.21" />
                    <SPLIT distance="100" swimtime="00:01:32.43" />
                    <SPLIT distance="125" swimtime="00:01:57.46" />
                    <SPLIT distance="150" swimtime="00:02:22.59" />
                    <SPLIT distance="175" swimtime="00:02:46.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="300" reactiontime="+69" swimtime="00:00:36.53" resultid="3461" lane="1" heatid="7037" entrytime="00:00:38.51">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="301" reactiontime="+86" swimtime="00:01:16.32" resultid="3457" lane="7" heatid="6736" entrytime="00:01:22.15">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.43" />
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                    <SPLIT distance="75" swimtime="00:00:58.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="291" reactiontime="+87" swimtime="00:03:12.25" resultid="3460" lane="1" heatid="7005" entrytime="00:03:37.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.05" />
                    <SPLIT distance="50" swimtime="00:00:41.93" />
                    <SPLIT distance="75" swimtime="00:01:06.28" />
                    <SPLIT distance="100" swimtime="00:01:31.09" />
                    <SPLIT distance="125" swimtime="00:01:56.19" />
                    <SPLIT distance="150" swimtime="00:02:22.06" />
                    <SPLIT distance="175" swimtime="00:02:47.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="317" reactiontime="+86" swimtime="00:00:33.67" resultid="3462" lane="4" heatid="7286" entrytime="00:00:34.25">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="385" reactiontime="+82" swimtime="00:00:29.23" resultid="3463" lane="4" heatid="7344" entrytime="00:00:29.99">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="355" reactiontime="+85" swimtime="00:01:06.39" resultid="3458" lane="5" heatid="6836" entrytime="00:01:10.52">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.38" />
                    <SPLIT distance="50" swimtime="00:00:30.80" />
                    <SPLIT distance="75" swimtime="00:00:48.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-02-27" firstname="Robert" gender="M" lastname="Lorkowski" nation="POL" athleteid="3464">
              <RESULTS>
                <RESULT eventid="1564" points="316" reactiontime="+87" swimtime="00:02:31.04" resultid="3468" lane="1" heatid="7061" entrytime="00:02:32.45">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.54" />
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                    <SPLIT distance="75" swimtime="00:00:51.43" />
                    <SPLIT distance="100" swimtime="00:01:10.97" />
                    <SPLIT distance="125" swimtime="00:01:30.89" />
                    <SPLIT distance="150" swimtime="00:01:51.35" />
                    <SPLIT distance="175" swimtime="00:02:11.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="303" reactiontime="+79" swimtime="00:02:49.95" resultid="3469" lane="2" heatid="7077" entrytime="00:02:53.71">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.19" />
                    <SPLIT distance="50" swimtime="00:00:37.88" />
                    <SPLIT distance="75" swimtime="00:00:59.77" />
                    <SPLIT distance="100" swimtime="00:01:21.52" />
                    <SPLIT distance="125" swimtime="00:01:46.67" />
                    <SPLIT distance="150" swimtime="00:02:11.99" />
                    <SPLIT distance="175" swimtime="00:02:31.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="279" reactiontime="+82" swimtime="00:06:13.04" resultid="3471" lane="3" heatid="7362" entrytime="00:06:18.24">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.66" />
                    <SPLIT distance="50" swimtime="00:00:39.85" />
                    <SPLIT distance="75" swimtime="00:01:04.00" />
                    <SPLIT distance="100" swimtime="00:01:28.98" />
                    <SPLIT distance="125" swimtime="00:01:53.70" />
                    <SPLIT distance="150" swimtime="00:02:17.66" />
                    <SPLIT distance="175" swimtime="00:02:41.72" />
                    <SPLIT distance="200" swimtime="00:03:05.43" />
                    <SPLIT distance="225" swimtime="00:03:32.36" />
                    <SPLIT distance="250" swimtime="00:03:58.68" />
                    <SPLIT distance="275" swimtime="00:04:25.22" />
                    <SPLIT distance="300" swimtime="00:04:51.58" />
                    <SPLIT distance="325" swimtime="00:05:12.70" />
                    <SPLIT distance="350" swimtime="00:05:33.55" />
                    <SPLIT distance="375" swimtime="00:05:54.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="204" reactiontime="+101" swimtime="00:03:10.21" resultid="3466" lane="7" heatid="6872" entrytime="00:03:13.74">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.78" />
                    <SPLIT distance="50" swimtime="00:00:39.72" />
                    <SPLIT distance="75" swimtime="00:01:03.41" />
                    <SPLIT distance="100" swimtime="00:01:27.56" />
                    <SPLIT distance="125" swimtime="00:01:53.18" />
                    <SPLIT distance="150" swimtime="00:02:18.82" />
                    <SPLIT distance="175" swimtime="00:02:44.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="280" swimtime="00:11:40.56" resultid="3465" lane="5" heatid="6719" entrytime="00:12:17.10" />
                <RESULT eventid="1730" status="DNS" swimtime="00:00:00.00" resultid="3470" lane="5" heatid="7322" entrytime="00:01:23.70" />
                <RESULT eventid="1375" status="DNS" swimtime="00:00:00.00" resultid="3467" lane="4" heatid="6904" entrytime="00:05:46.11" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-11-29" firstname="Jarosław" gender="M" lastname="Niedbałowski" nation="POL" athleteid="3472">
              <RESULTS>
                <RESULT eventid="1696" points="344" reactiontime="+79" swimtime="00:01:24.03" resultid="3476" heatid="7308" entrytime="00:01:25.87">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.16" />
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                    <SPLIT distance="75" swimtime="00:01:00.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="292" reactiontime="+82" swimtime="00:03:11.99" resultid="3475" lane="5" heatid="7007" entrytime="00:03:16.17">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.13" />
                    <SPLIT distance="50" swimtime="00:00:42.42" />
                    <SPLIT distance="75" swimtime="00:01:06.30" />
                    <SPLIT distance="100" swimtime="00:01:31.38" />
                    <SPLIT distance="125" swimtime="00:01:56.33" />
                    <SPLIT distance="150" swimtime="00:02:22.09" />
                    <SPLIT distance="175" swimtime="00:02:47.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="380" reactiontime="+79" swimtime="00:00:37.50" resultid="3474" lane="5" heatid="6860" entrytime="00:00:38.12">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="292" reactiontime="+77" swimtime="00:00:32.06" resultid="3477" heatid="7342" entrytime="00:00:31.53">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="3473" lane="2" heatid="6735" entrytime="00:01:25.01" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-06-04" firstname="Paweł" gender="M" lastname="Opaliński" nation="POL" athleteid="3478">
              <RESULTS>
                <RESULT eventid="1696" points="455" reactiontime="+78" swimtime="00:01:16.56" resultid="3485" lane="4" heatid="7309" entrytime="00:01:19.77">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.35" />
                    <SPLIT distance="50" swimtime="00:00:35.62" />
                    <SPLIT distance="75" swimtime="00:00:55.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="419" reactiontime="+84" swimtime="00:04:54.10" resultid="3481" lane="1" heatid="6907" entrytime="00:05:15.95">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.09" />
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                    <SPLIT distance="75" swimtime="00:00:50.04" />
                    <SPLIT distance="100" swimtime="00:01:08.17" />
                    <SPLIT distance="125" swimtime="00:01:26.74" />
                    <SPLIT distance="150" swimtime="00:01:45.48" />
                    <SPLIT distance="175" swimtime="00:02:04.11" />
                    <SPLIT distance="200" swimtime="00:02:23.31" />
                    <SPLIT distance="225" swimtime="00:02:42.24" />
                    <SPLIT distance="250" swimtime="00:03:01.48" />
                    <SPLIT distance="275" swimtime="00:03:20.33" />
                    <SPLIT distance="300" swimtime="00:03:39.71" />
                    <SPLIT distance="325" swimtime="00:03:58.74" />
                    <SPLIT distance="350" swimtime="00:04:18.73" />
                    <SPLIT distance="375" swimtime="00:04:37.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="360" reactiontime="+84" swimtime="00:01:10.79" resultid="3482" heatid="7021" entrytime="00:01:11.73">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.42" />
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                    <SPLIT distance="75" swimtime="00:00:51.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="336" swimtime="00:10:59.32" resultid="3479" lane="7" heatid="6721" entrytime="00:11:16.27" />
                <RESULT eventid="1564" points="444" reactiontime="+82" swimtime="00:02:14.90" resultid="3483" lane="3" heatid="7063" entrytime="00:02:18.77">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.39" />
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                    <SPLIT distance="75" swimtime="00:00:46.97" />
                    <SPLIT distance="100" swimtime="00:01:04.08" />
                    <SPLIT distance="125" swimtime="00:01:21.74" />
                    <SPLIT distance="150" swimtime="00:01:39.89" />
                    <SPLIT distance="175" swimtime="00:01:57.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="419" reactiontime="+79" swimtime="00:00:30.68" resultid="3484" lane="8" heatid="7289" entrytime="00:00:31.72">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="447" reactiontime="+79" swimtime="00:01:01.49" resultid="3480" lane="8" heatid="6842" entrytime="00:01:02.76">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.63" />
                    <SPLIT distance="50" swimtime="00:00:28.91" />
                    <SPLIT distance="75" swimtime="00:00:45.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-06-26" firstname="Krzysztof" gender="M" lastname="Pawłowski" nation="POL" athleteid="3486">
              <RESULTS>
                <RESULT eventid="1798" points="287" reactiontime="+79" swimtime="00:06:09.38" resultid="3493" lane="2" heatid="7362" entrytime="00:06:20.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.89" />
                    <SPLIT distance="50" swimtime="00:00:40.11" />
                    <SPLIT distance="75" swimtime="00:01:03.97" />
                    <SPLIT distance="100" swimtime="00:01:29.72" />
                    <SPLIT distance="125" swimtime="00:01:54.28" />
                    <SPLIT distance="150" swimtime="00:02:18.27" />
                    <SPLIT distance="175" swimtime="00:02:41.90" />
                    <SPLIT distance="200" swimtime="00:03:05.87" />
                    <SPLIT distance="225" swimtime="00:03:30.74" />
                    <SPLIT distance="250" swimtime="00:03:56.43" />
                    <SPLIT distance="275" swimtime="00:04:22.00" />
                    <SPLIT distance="300" swimtime="00:04:48.27" />
                    <SPLIT distance="325" swimtime="00:05:09.33" />
                    <SPLIT distance="350" swimtime="00:05:29.95" />
                    <SPLIT distance="375" swimtime="00:05:50.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="274" swimtime="00:11:45.53" resultid="3487" lane="7" heatid="6720" entrytime="00:12:05.30" />
                <RESULT eventid="1411" points="324" reactiontime="+78" swimtime="00:03:05.58" resultid="3490" lane="7" heatid="7008" entrytime="00:03:10.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.63" />
                    <SPLIT distance="50" swimtime="00:00:42.22" />
                    <SPLIT distance="75" swimtime="00:01:05.98" />
                    <SPLIT distance="100" swimtime="00:01:30.00" />
                    <SPLIT distance="125" swimtime="00:01:54.32" />
                    <SPLIT distance="150" swimtime="00:02:18.88" />
                    <SPLIT distance="175" swimtime="00:02:42.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="299" reactiontime="+74" swimtime="00:02:50.32" resultid="3488" lane="4" heatid="6884" entrytime="00:02:57.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.51" />
                    <SPLIT distance="50" swimtime="00:00:40.27" />
                    <SPLIT distance="75" swimtime="00:01:01.92" />
                    <SPLIT distance="100" swimtime="00:01:23.75" />
                    <SPLIT distance="125" swimtime="00:01:45.85" />
                    <SPLIT distance="150" swimtime="00:02:07.78" />
                    <SPLIT distance="175" swimtime="00:02:29.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="356" reactiontime="+81" swimtime="00:01:23.09" resultid="3492" lane="3" heatid="7307" entrytime="00:01:26.45">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.92" />
                    <SPLIT distance="50" swimtime="00:00:39.16" />
                    <SPLIT distance="75" swimtime="00:01:00.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="310" reactiontime="+84" swimtime="00:02:48.68" resultid="3491" lane="7" heatid="7077" entrytime="00:02:55.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.46" />
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                    <SPLIT distance="75" swimtime="00:00:59.54" />
                    <SPLIT distance="100" swimtime="00:01:21.62" />
                    <SPLIT distance="125" swimtime="00:01:46.16" />
                    <SPLIT distance="150" swimtime="00:02:10.31" />
                    <SPLIT distance="175" swimtime="00:02:30.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="303" reactiontime="+82" swimtime="00:05:27.41" resultid="3489" heatid="6905" entrytime="00:05:45.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.12" />
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                    <SPLIT distance="75" swimtime="00:00:56.21" />
                    <SPLIT distance="100" swimtime="00:01:16.92" />
                    <SPLIT distance="125" swimtime="00:01:37.46" />
                    <SPLIT distance="150" swimtime="00:01:58.63" />
                    <SPLIT distance="175" swimtime="00:02:19.33" />
                    <SPLIT distance="200" swimtime="00:02:40.53" />
                    <SPLIT distance="225" swimtime="00:03:01.59" />
                    <SPLIT distance="250" swimtime="00:03:23.17" />
                    <SPLIT distance="275" swimtime="00:03:44.26" />
                    <SPLIT distance="300" swimtime="00:04:05.38" />
                    <SPLIT distance="325" swimtime="00:04:25.67" />
                    <SPLIT distance="350" swimtime="00:04:46.72" />
                    <SPLIT distance="375" swimtime="00:05:06.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-04-17" firstname="Maria" gender="F" lastname="Petecka" nation="POL" athleteid="3494">
              <RESULTS>
                <RESULT eventid="1679" points="305" reactiontime="+76" swimtime="00:01:36.68" resultid="3500" lane="5" heatid="7299" entrytime="00:01:36.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.37" />
                    <SPLIT distance="50" swimtime="00:00:45.82" />
                    <SPLIT distance="75" swimtime="00:01:11.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="298" reactiontime="+89" swimtime="00:00:38.08" resultid="3499" lane="2" heatid="7278" entrytime="00:00:39.11">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1581" points="275" reactiontime="+87" swimtime="00:03:17.45" resultid="3498" lane="4" heatid="7069" entrytime="00:03:16.05">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.46" />
                    <SPLIT distance="50" swimtime="00:00:41.28" />
                    <SPLIT distance="75" swimtime="00:01:09.31" />
                    <SPLIT distance="100" swimtime="00:01:35.49" />
                    <SPLIT distance="125" swimtime="00:02:03.22" />
                    <SPLIT distance="150" swimtime="00:02:30.51" />
                    <SPLIT distance="175" swimtime="00:02:55.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="313" reactiontime="+86" swimtime="00:00:44.64" resultid="3496" lane="7" heatid="6851" entrytime="00:00:46.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="290" reactiontime="+88" swimtime="00:01:28.75" resultid="3495" heatid="6727" entrytime="00:01:28.01">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.06" />
                    <SPLIT distance="50" swimtime="00:00:41.82" />
                    <SPLIT distance="75" swimtime="00:01:07.08" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K 11" eventid="1409" reactiontime="+89" status="DSQ" swimtime="00:00:00.00" resultid="3497" lane="6" heatid="7000" entrytime="00:03:28.03">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.82" />
                    <SPLIT distance="50" swimtime="00:00:46.90" />
                    <SPLIT distance="75" swimtime="00:01:13.04" />
                    <SPLIT distance="100" swimtime="00:01:40.16" />
                    <SPLIT distance="125" swimtime="00:02:07.96" />
                    <SPLIT distance="150" swimtime="00:02:35.26" />
                    <SPLIT distance="175" swimtime="00:03:02.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-03-12" firstname="Adam" gender="M" lastname="Przybylski" nation="POL" athleteid="3501">
              <RESULTS>
                <RESULT eventid="1598" points="249" reactiontime="+89" swimtime="00:03:01.50" resultid="3506" lane="7" heatid="7075" entrytime="00:03:15.11">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.29" />
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                    <SPLIT distance="75" swimtime="00:01:01.47" />
                    <SPLIT distance="100" swimtime="00:01:24.88" />
                    <SPLIT distance="125" swimtime="00:01:52.63" />
                    <SPLIT distance="150" swimtime="00:02:19.90" />
                    <SPLIT distance="175" swimtime="00:02:41.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="259" reactiontime="+56" swimtime="00:01:22.41" resultid="3507" lane="1" heatid="7321" entrytime="00:01:38.83">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.22" />
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                    <SPLIT distance="75" swimtime="00:01:01.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="254" swimtime="00:12:03.75" resultid="3502" lane="8" heatid="6720" entrytime="00:12:10.73" />
                <RESULT eventid="1564" points="288" reactiontime="+84" swimtime="00:02:35.83" resultid="3505" heatid="7059" entrytime="00:02:41.31">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.45" />
                    <SPLIT distance="50" swimtime="00:00:33.97" />
                    <SPLIT distance="75" swimtime="00:00:52.97" />
                    <SPLIT distance="100" swimtime="00:01:13.18" />
                    <SPLIT distance="125" swimtime="00:01:33.58" />
                    <SPLIT distance="150" swimtime="00:01:55.01" />
                    <SPLIT distance="175" swimtime="00:02:15.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="361" reactiontime="+84" swimtime="00:00:29.88" resultid="3508" lane="1" heatid="7345" entrytime="00:00:29.02">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="325" reactiontime="+87" swimtime="00:01:08.39" resultid="3503" lane="1" heatid="6833" entrytime="00:01:20.11">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.01" />
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                    <SPLIT distance="75" swimtime="00:00:51.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="3504" lane="3" heatid="6871" entrytime="00:03:21.12" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-04-15" firstname="Michał" gender="M" lastname="Skrok" nation="POL" athleteid="3509">
              <RESULTS>
                <RESULT eventid="1411" points="453" reactiontime="+82" swimtime="00:02:45.92" resultid="3513" lane="3" heatid="7010" entrytime="00:02:53.11">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.04" />
                    <SPLIT distance="50" swimtime="00:00:37.43" />
                    <SPLIT distance="75" swimtime="00:00:58.09" />
                    <SPLIT distance="100" swimtime="00:01:18.90" />
                    <SPLIT distance="125" swimtime="00:01:39.91" />
                    <SPLIT distance="150" swimtime="00:02:01.27" />
                    <SPLIT distance="175" swimtime="00:02:23.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="534" reactiontime="+77" swimtime="00:00:33.50" resultid="3511" lane="8" heatid="6865" entrytime="00:00:34.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="440" reactiontime="+84" swimtime="00:02:30.14" resultid="3514" lane="1" heatid="7079" entrytime="00:02:33.53">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.02" />
                    <SPLIT distance="50" swimtime="00:00:31.10" />
                    <SPLIT distance="75" swimtime="00:00:51.62" />
                    <SPLIT distance="100" swimtime="00:01:11.75" />
                    <SPLIT distance="125" swimtime="00:01:32.46" />
                    <SPLIT distance="150" swimtime="00:01:53.68" />
                    <SPLIT distance="175" swimtime="00:02:12.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="485" reactiontime="+73" swimtime="00:01:14.95" resultid="3515" lane="5" heatid="7310" entrytime="00:01:15.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.86" />
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                    <SPLIT distance="75" swimtime="00:00:54.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="404" reactiontime="+69" swimtime="00:02:34.10" resultid="3512" heatid="6886" entrytime="00:02:40.11">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.77" />
                    <SPLIT distance="50" swimtime="00:00:36.50" />
                    <SPLIT distance="75" swimtime="00:00:55.77" />
                    <SPLIT distance="100" swimtime="00:01:15.23" />
                    <SPLIT distance="125" swimtime="00:01:35.14" />
                    <SPLIT distance="150" swimtime="00:01:54.92" />
                    <SPLIT distance="175" swimtime="00:02:14.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="450" reactiontime="+73" swimtime="00:01:06.73" resultid="3510" heatid="6743" entrytime="00:01:08.33">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.66" />
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                    <SPLIT distance="75" swimtime="00:00:50.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" status="DNS" swimtime="00:00:00.00" resultid="3516" lane="7" heatid="7363" entrytime="00:06:10.70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-06-07" firstname="Wiesław" gender="M" lastname="Bar" nation="POL" athleteid="3517">
              <RESULTS>
                <RESULT eventid="1143" points="319" swimtime="00:21:19.24" resultid="3518" lane="1" heatid="6752" entrytime="00:21:01.10" />
                <RESULT eventid="1375" points="380" reactiontime="+95" swimtime="00:05:03.60" resultid="3520" lane="6" heatid="6907" entrytime="00:05:13.11">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.09" />
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                    <SPLIT distance="75" swimtime="00:00:50.25" />
                    <SPLIT distance="100" swimtime="00:01:08.42" />
                    <SPLIT distance="125" swimtime="00:01:27.32" />
                    <SPLIT distance="150" swimtime="00:01:46.43" />
                    <SPLIT distance="175" swimtime="00:02:05.82" />
                    <SPLIT distance="200" swimtime="00:02:25.13" />
                    <SPLIT distance="225" swimtime="00:02:44.97" />
                    <SPLIT distance="250" swimtime="00:03:04.68" />
                    <SPLIT distance="275" swimtime="00:03:24.87" />
                    <SPLIT distance="300" swimtime="00:03:45.05" />
                    <SPLIT distance="325" swimtime="00:04:04.71" />
                    <SPLIT distance="350" swimtime="00:04:24.89" />
                    <SPLIT distance="375" swimtime="00:04:45.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="342" reactiontime="+91" swimtime="00:05:48.41" resultid="3524" lane="4" heatid="7362" entrytime="00:06:15.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.15" />
                    <SPLIT distance="50" swimtime="00:00:34.00" />
                    <SPLIT distance="75" swimtime="00:00:54.44" />
                    <SPLIT distance="100" swimtime="00:01:16.49" />
                    <SPLIT distance="125" swimtime="00:01:39.11" />
                    <SPLIT distance="150" swimtime="00:02:01.52" />
                    <SPLIT distance="175" swimtime="00:02:24.44" />
                    <SPLIT distance="200" swimtime="00:02:47.25" />
                    <SPLIT distance="225" swimtime="00:03:12.83" />
                    <SPLIT distance="250" swimtime="00:03:38.61" />
                    <SPLIT distance="275" swimtime="00:04:04.03" />
                    <SPLIT distance="300" swimtime="00:04:29.93" />
                    <SPLIT distance="325" swimtime="00:04:50.27" />
                    <SPLIT distance="350" swimtime="00:05:10.92" />
                    <SPLIT distance="375" swimtime="00:05:30.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="407" reactiontime="+83" swimtime="00:02:18.88" resultid="3522" lane="2" heatid="7063" entrytime="00:02:19.11">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.46" />
                    <SPLIT distance="50" swimtime="00:00:30.70" />
                    <SPLIT distance="75" swimtime="00:00:47.81" />
                    <SPLIT distance="100" swimtime="00:01:05.00" />
                    <SPLIT distance="125" swimtime="00:01:23.21" />
                    <SPLIT distance="150" swimtime="00:01:41.87" />
                    <SPLIT distance="175" swimtime="00:02:00.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="466" reactiontime="+83" swimtime="00:00:27.44" resultid="3523" lane="3" heatid="7349" entrytime="00:00:27.51">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="451" reactiontime="+84" swimtime="00:01:01.32" resultid="3519" heatid="6842" entrytime="00:01:02.18">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.86" />
                    <SPLIT distance="50" swimtime="00:00:29.32" />
                    <SPLIT distance="75" swimtime="00:00:45.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="342" reactiontime="+83" swimtime="00:01:12.03" resultid="3521" lane="7" heatid="7022" entrytime="00:01:07.01">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.47" />
                    <SPLIT distance="50" swimtime="00:00:32.26" />
                    <SPLIT distance="75" swimtime="00:00:51.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1177" points="512" reactiontime="+87" swimtime="00:01:48.44" resultid="3525" lane="8" heatid="6810" entrytime="00:01:51.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.06" />
                    <SPLIT distance="50" swimtime="00:00:26.58" />
                    <SPLIT distance="75" swimtime="00:00:39.99" />
                    <SPLIT distance="100" swimtime="00:00:54.47" />
                    <SPLIT distance="125" swimtime="00:01:07.77" />
                    <SPLIT distance="150" swimtime="00:01:21.92" />
                    <SPLIT distance="175" swimtime="00:01:34.63" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3416" number="1" reactiontime="+87" />
                    <RELAYPOSITION athleteid="3509" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="3478" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="3424" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1177" points="404" reactiontime="+82" swimtime="00:01:57.30" resultid="3526" lane="6" heatid="6809" entrytime="00:01:55.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.03" />
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                    <SPLIT distance="75" swimtime="00:00:44.35" />
                    <SPLIT distance="100" swimtime="00:01:00.53" />
                    <SPLIT distance="125" swimtime="00:01:13.83" />
                    <SPLIT distance="150" swimtime="00:01:28.59" />
                    <SPLIT distance="175" swimtime="00:01:42.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3456" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="3432" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="3517" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="3501" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1177" points="360" reactiontime="+82" swimtime="00:02:01.95" resultid="3527" lane="6" heatid="6808" entrytime="00:02:05.11">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.61" />
                    <SPLIT distance="50" swimtime="00:00:30.31" />
                    <SPLIT distance="75" swimtime="00:00:45.45" />
                    <SPLIT distance="100" swimtime="00:01:01.73" />
                    <SPLIT distance="125" swimtime="00:01:15.17" />
                    <SPLIT distance="150" swimtime="00:01:30.45" />
                    <SPLIT distance="175" swimtime="00:01:45.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3464" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="3472" number="2" reactiontime="+33" />
                    <RELAYPOSITION athleteid="3486" number="3" reactiontime="+15" />
                    <RELAYPOSITION athleteid="3448" number="4" reactiontime="+18" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1341" points="502" reactiontime="+71" swimtime="00:02:00.13" resultid="3528" lane="3" heatid="6987" entrytime="00:02:05.41">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.80" />
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                    <SPLIT distance="75" swimtime="00:00:46.86" />
                    <SPLIT distance="100" swimtime="00:01:04.95" />
                    <SPLIT distance="125" swimtime="00:01:17.82" />
                    <SPLIT distance="150" swimtime="00:01:32.85" />
                    <SPLIT distance="175" swimtime="00:01:45.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3416" number="1" reactiontime="+71" />
                    <RELAYPOSITION athleteid="3509" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="3424" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="3478" number="4" reactiontime="+70" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="5">
              <RESULTS>
                <RESULT eventid="1341" points="351" reactiontime="+77" swimtime="00:02:15.34" resultid="3529" heatid="6987" entrytime="00:02:15.11">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.12" />
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                    <SPLIT distance="75" swimtime="00:00:54.63" />
                    <SPLIT distance="100" swimtime="00:01:15.32" />
                    <SPLIT distance="125" swimtime="00:01:29.45" />
                    <SPLIT distance="150" swimtime="00:01:46.74" />
                    <SPLIT distance="175" swimtime="00:02:00.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3456" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="3432" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="3517" number="3" reactiontime="+49" />
                    <RELAYPOSITION athleteid="3501" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" number="6">
              <RESULTS>
                <RESULT eventid="1341" points="300" reactiontime="+92" swimtime="00:02:22.52" resultid="3530" lane="6" heatid="6986" entrytime="00:02:23.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.97" />
                    <SPLIT distance="50" swimtime="00:00:38.04" />
                    <SPLIT distance="75" swimtime="00:00:55.31" />
                    <SPLIT distance="100" swimtime="00:00:58.46" />
                    <SPLIT distance="125" swimtime="00:01:31.37" />
                    <SPLIT distance="150" swimtime="00:01:50.20" />
                    <SPLIT distance="175" swimtime="00:02:06.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3464" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="3472" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="3486" number="3" />
                    <RELAYPOSITION athleteid="3448" number="4" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="RESWIE" name="Klub Sportowy &quot;Rekin&quot; Świebodzice" nation="POL" region="DOL">
          <CONTACT city="ŚWIEBODZICE" name="WINIARCZYK" phone="606626274" state="DOLNO" street="MIESZKA STAREGO 4" zip="58-160" />
          <ATHLETES>
            <ATHLETE birthdate="1982-01-01" firstname="Tomasz" gender="M" lastname="Karch" nation="POL" athleteid="3555">
              <RESULTS>
                <RESULT comment="przekroczony limit 20:00:00" eventid="1143" status="DSQ" swimtime="00:22:26.66" resultid="3556" lane="8" heatid="6752" entrytime="00:21:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SAKIE" name="Salos Kielce" nation="POL">
          <CONTACT name="Kijewska" phone="606 760616" street="Iwona" />
          <ATHLETES>
            <ATHLETE birthdate="1957-07-30" firstname="Stefan" gender="M" lastname="Najgeburski" nation="POL" athleteid="3562">
              <RESULTS>
                <RESULT eventid="1143" points="249" swimtime="00:23:09.62" resultid="3563" lane="7" heatid="6751" entrytime="00:23:00.00" />
                <RESULT eventid="1564" points="234" reactiontime="+79" swimtime="00:02:47.06" resultid="3566" lane="1" heatid="7058" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.46" />
                    <SPLIT distance="50" swimtime="00:00:37.14" />
                    <SPLIT distance="75" swimtime="00:00:57.76" />
                    <SPLIT distance="100" swimtime="00:01:19.49" />
                    <SPLIT distance="125" swimtime="00:01:41.24" />
                    <SPLIT distance="150" swimtime="00:02:03.83" />
                    <SPLIT distance="175" swimtime="00:02:26.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="162" reactiontime="+84" swimtime="00:01:32.45" resultid="3565" lane="1" heatid="7018" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.83" />
                    <SPLIT distance="50" swimtime="00:00:42.78" />
                    <SPLIT distance="75" swimtime="00:01:07.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="245" reactiontime="+75" swimtime="00:05:51.55" resultid="3564" lane="8" heatid="6905" entrytime="00:05:46.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.84" />
                    <SPLIT distance="50" swimtime="00:00:38.00" />
                    <SPLIT distance="75" swimtime="00:00:59.48" />
                    <SPLIT distance="100" swimtime="00:01:20.90" />
                    <SPLIT distance="125" swimtime="00:01:43.12" />
                    <SPLIT distance="150" swimtime="00:02:05.49" />
                    <SPLIT distance="175" swimtime="00:02:28.19" />
                    <SPLIT distance="200" swimtime="00:02:51.18" />
                    <SPLIT distance="225" swimtime="00:03:14.47" />
                    <SPLIT distance="250" swimtime="00:03:36.82" />
                    <SPLIT distance="275" swimtime="00:03:59.40" />
                    <SPLIT distance="300" swimtime="00:04:22.17" />
                    <SPLIT distance="325" swimtime="00:04:44.79" />
                    <SPLIT distance="350" swimtime="00:05:07.60" />
                    <SPLIT distance="375" swimtime="00:05:30.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="216" reactiontime="+77" swimtime="00:06:45.80" resultid="3567" lane="1" heatid="7361" entrytime="00:06:46.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.61" />
                    <SPLIT distance="50" swimtime="00:00:45.13" />
                    <SPLIT distance="75" swimtime="00:01:11.66" />
                    <SPLIT distance="100" swimtime="00:01:39.43" />
                    <SPLIT distance="125" swimtime="00:02:07.36" />
                    <SPLIT distance="150" swimtime="00:02:34.19" />
                    <SPLIT distance="175" swimtime="00:03:00.71" />
                    <SPLIT distance="200" swimtime="00:03:26.63" />
                    <SPLIT distance="225" swimtime="00:03:54.49" />
                    <SPLIT distance="250" swimtime="00:04:22.43" />
                    <SPLIT distance="275" swimtime="00:04:50.20" />
                    <SPLIT distance="300" swimtime="00:05:18.24" />
                    <SPLIT distance="325" swimtime="00:05:40.89" />
                    <SPLIT distance="350" swimtime="00:06:02.93" />
                    <SPLIT distance="375" swimtime="00:06:25.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-05-17" firstname="Iwona" gender="F" lastname="Kijewska" nation="POL" athleteid="3568">
              <RESULTS>
                <RESULT eventid="1679" points="324" reactiontime="+88" swimtime="00:01:34.75" resultid="3575" lane="2" heatid="7299" entrytime="00:01:36.78">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.65" />
                    <SPLIT distance="50" swimtime="00:00:44.80" />
                    <SPLIT distance="75" swimtime="00:01:09.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="309" reactiontime="+88" swimtime="00:00:37.65" resultid="3574" lane="3" heatid="7278" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1445" points="232" reactiontime="+98" swimtime="00:01:32.05" resultid="3572" lane="4" heatid="7013" entrytime="00:01:27.67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.40" />
                    <SPLIT distance="50" swimtime="00:00:43.39" />
                    <SPLIT distance="75" swimtime="00:01:07.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1581" points="294" reactiontime="+91" swimtime="00:03:13.03" resultid="3573" lane="6" heatid="7070" entrytime="00:03:08.32">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.07" />
                    <SPLIT distance="50" swimtime="00:00:39.89" />
                    <SPLIT distance="75" swimtime="00:01:06.61" />
                    <SPLIT distance="100" swimtime="00:01:32.68" />
                    <SPLIT distance="125" swimtime="00:01:59.45" />
                    <SPLIT distance="150" swimtime="00:02:26.30" />
                    <SPLIT distance="175" swimtime="00:02:50.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="339" reactiontime="+91" swimtime="00:00:43.45" resultid="3570" lane="4" heatid="6851" entrytime="00:00:44.32">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="322" reactiontime="+96" swimtime="00:01:25.78" resultid="3569" lane="7" heatid="6727" entrytime="00:01:27.56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.64" />
                    <SPLIT distance="50" swimtime="00:00:40.51" />
                    <SPLIT distance="75" swimtime="00:01:05.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" status="DNS" swimtime="00:00:00.00" resultid="3571" lane="3" heatid="6896" entrytime="00:06:10.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SIGLI" name="Sikret Gliwice" nation="POL">
          <CONTACT city="GLIWICE" email="J.ZAGALA@ECOTRADE.PL" name="ZAGAŁA JOANNA" phone="601427257" street="JAGIELOŃSKA 21" zip="44-100" />
          <ATHLETES>
            <ATHLETE birthdate="1958-02-05" firstname="Zofia" gender="F" lastname="Dąbrowska" nation="POL" athleteid="3577">
              <RESULTS>
                <RESULT eventid="1222" points="212" reactiontime="+89" swimtime="00:00:50.76" resultid="3579" lane="3" heatid="6849" entrytime="00:00:52.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1581" points="139" reactiontime="+97" swimtime="00:04:07.71" resultid="3581" lane="8" heatid="7068" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.39" />
                    <SPLIT distance="50" swimtime="00:00:50.56" />
                    <SPLIT distance="75" swimtime="00:01:24.93" />
                    <SPLIT distance="100" swimtime="00:02:00.60" />
                    <SPLIT distance="125" swimtime="00:02:32.87" />
                    <SPLIT distance="150" swimtime="00:03:06.26" />
                    <SPLIT distance="175" swimtime="00:03:39.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="160" reactiontime="+83" swimtime="00:01:48.21" resultid="3578" heatid="6725" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.52" />
                    <SPLIT distance="50" swimtime="00:00:51.48" />
                    <SPLIT distance="75" swimtime="00:01:20.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="155" reactiontime="+93" swimtime="00:00:47.31" resultid="3582" lane="1" heatid="7277" entrytime="00:00:46.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="209" reactiontime="+89" swimtime="00:00:40.36" resultid="3583" lane="5" heatid="7330" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.11" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="przekroczony limit 8:30:00" eventid="1358" reactiontime="+107" status="DSQ" swimtime="00:00:00.00" resultid="3580" lane="4" heatid="6894" entrytime="00:07:42.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.96" />
                    <SPLIT distance="50" swimtime="00:00:45.59" />
                    <SPLIT distance="75" swimtime="00:01:12.70" />
                    <SPLIT distance="100" swimtime="00:01:41.47" />
                    <SPLIT distance="125" swimtime="00:02:12.27" />
                    <SPLIT distance="150" swimtime="00:02:43.18" />
                    <SPLIT distance="175" swimtime="00:03:14.57" />
                    <SPLIT distance="200" swimtime="00:03:45.24" />
                    <SPLIT distance="225" swimtime="00:04:16.82" />
                    <SPLIT distance="250" swimtime="00:04:49.12" />
                    <SPLIT distance="275" swimtime="00:05:22.20" />
                    <SPLIT distance="300" swimtime="00:05:57.77" />
                    <SPLIT distance="325" swimtime="00:07:31.17" />
                    <SPLIT distance="350" swimtime="00:07:00.87" />
                    <SPLIT distance="375" swimtime="00:08:32.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SIWAR" name="Sinnet T.C. Warszawa" nation="POL">
          <CONTACT city="Warszawa" email="piotrbarski@uw.edu.pl" name="Barski" phone="603976435" street="Polinezyjska 5/71" zip="02-777" />
          <ATHLETES>
            <ATHLETE birthdate="1965-01-01" firstname="Piotr" gender="M" lastname="Barski" nation="POL" athleteid="3590">
              <RESULTS>
                <RESULT comment="Rekord Polski " eventid="1205" points="551" reactiontime="+80" swimtime="00:00:57.39" resultid="3592" lane="6" heatid="6830" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.41" />
                    <SPLIT distance="50" swimtime="00:00:28.06" />
                    <SPLIT distance="75" swimtime="00:00:42.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="520" reactiontime="+80" swimtime="00:00:26.45" resultid="3596" lane="2" heatid="7353" entrytime="00:00:25.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="476" reactiontime="+73" swimtime="00:01:15.41" resultid="3595" lane="8" heatid="7311" entrytime="00:01:12.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.90" />
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                    <SPLIT distance="75" swimtime="00:00:55.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="476" reactiontime="+83" swimtime="00:02:43.20" resultid="3594" heatid="7011" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.18" />
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                    <SPLIT distance="75" swimtime="00:00:57.72" />
                    <SPLIT distance="100" swimtime="00:01:18.87" />
                    <SPLIT distance="125" swimtime="00:01:40.13" />
                    <SPLIT distance="150" swimtime="00:02:01.34" />
                    <SPLIT distance="175" swimtime="00:02:22.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="589" reactiontime="+77" swimtime="00:00:32.42" resultid="3593" lane="1" heatid="6866" entrytime="00:00:31.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="429" reactiontime="+81" swimtime="00:01:07.80" resultid="3591" lane="6" heatid="6744" entrytime="00:01:06.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.84" />
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                    <SPLIT distance="75" swimtime="00:00:52.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="JSJEL" name="MUKP Just Swim Jelenia Góra" nation="POL" region="WR">
          <CONTACT city="Jelenia Góra" email="szymon.kurowski@justswim.pl" fax="+48 75 64 523 01" internet="www.justswim.pl" name="Szymon Kurowski" phone="+48 609 669 129" state="DOL" street="al. Wojska Polskiego 21" zip="58-500" />
          <ATHLETES>
            <ATHLETE birthdate="1983-05-01" firstname="Andrei" gender="M" lastname="Vashkevich" nation="POL" athleteid="3598">
              <RESULTS>
                <RESULT eventid="1645" points="687" reactiontime="+89" swimtime="00:00:26.01" resultid="3600" lane="6" heatid="7294" entrytime="00:00:26.24">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="692" reactiontime="+85" swimtime="00:00:24.05" resultid="3601" lane="2" heatid="7354" entrytime="00:00:24.44">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" status="DNS" swimtime="00:00:00.00" resultid="3599" lane="6" heatid="7041" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TOTOR" name="Toruńczyk Masters Toruń" nation="POL" region="KUJ">
          <CONTACT city="Toruń" email="szufar@o2.pl" name="Szufarski Andrzej" phone="600898866" state="KUJ-P" street="Matejki 60/7" zip="87-100" />
          <ATHLETES>
            <ATHLETE birthdate="1940-01-01" firstname="Edward" gender="M" lastname="Korolko" nation="POL" athleteid="3603">
              <RESULTS>
                <RESULT eventid="1205" points="126" reactiontime="+98" swimtime="00:01:33.63" resultid="3604" lane="2" heatid="6831" entrytime="00:01:33.25">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.08" />
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                    <SPLIT distance="75" swimtime="00:01:07.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="89" reactiontime="+106" swimtime="00:03:50.26" resultid="3607" heatid="7055" entrytime="00:03:40.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.13" />
                    <SPLIT distance="50" swimtime="00:00:49.07" />
                    <SPLIT distance="75" swimtime="00:01:18.29" />
                    <SPLIT distance="100" swimtime="00:01:49.25" />
                    <SPLIT distance="125" swimtime="00:02:19.62" />
                    <SPLIT distance="150" swimtime="00:02:49.82" />
                    <SPLIT distance="175" swimtime="00:03:19.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="75" reactiontime="+68" swimtime="00:00:57.78" resultid="3606" lane="1" heatid="7033" entrytime="00:00:56.25">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="68" reactiontime="+77" swimtime="00:02:08.11" resultid="3608" lane="7" heatid="7319" entrytime="00:02:07.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.59" />
                    <SPLIT distance="50" swimtime="00:01:01.33" />
                    <SPLIT distance="75" swimtime="00:01:36.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" status="DNS" swimtime="00:00:00.00" resultid="3605" lane="1" heatid="6881" entrytime="00:04:35.36" />
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="3609" lane="7" heatid="7337" entrytime="00:00:40.10" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-01" firstname="Jan" gender="M" lastname="Bantkowski" nation="POL" athleteid="3610">
              <RESULTS>
                <RESULT eventid="1564" points="99" reactiontime="+111" swimtime="00:03:42.32" resultid="3615" lane="3" heatid="7055" entrytime="00:03:28.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.52" />
                    <SPLIT distance="50" swimtime="00:00:47.61" />
                    <SPLIT distance="75" swimtime="00:01:15.98" />
                    <SPLIT distance="100" swimtime="00:01:44.48" />
                    <SPLIT distance="125" swimtime="00:02:14.86" />
                    <SPLIT distance="150" swimtime="00:02:45.08" />
                    <SPLIT distance="175" swimtime="00:03:14.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="119" reactiontime="+128" swimtime="00:01:59.47" resultid="3616" lane="2" heatid="7302" entrytime="00:02:03.54">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.72" />
                    <SPLIT distance="50" swimtime="00:00:56.73" />
                    <SPLIT distance="75" swimtime="00:01:27.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="53" reactiontime="+100" swimtime="00:05:01.90" resultid="3613" lane="6" heatid="6881" entrytime="00:04:32.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.29" />
                    <SPLIT distance="50" swimtime="00:01:10.94" />
                    <SPLIT distance="75" swimtime="00:01:49.29" />
                    <SPLIT distance="100" swimtime="00:02:28.26" />
                    <SPLIT distance="125" swimtime="00:03:06.22" />
                    <SPLIT distance="150" swimtime="00:03:44.95" />
                    <SPLIT distance="175" swimtime="00:04:23.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="100" reactiontime="+123" swimtime="00:04:34.71" resultid="3614" lane="1" heatid="7003" entrytime="00:04:15.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.95" />
                    <SPLIT distance="50" swimtime="00:01:03.51" />
                    <SPLIT distance="75" swimtime="00:01:38.93" />
                    <SPLIT distance="100" swimtime="00:02:14.01" />
                    <SPLIT distance="125" swimtime="00:02:49.99" />
                    <SPLIT distance="150" swimtime="00:03:24.89" />
                    <SPLIT distance="175" swimtime="00:04:00.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="3611" lane="5" heatid="6731" entrytime="00:01:48.60" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="3612" lane="5" heatid="6869" entrytime="00:04:38.42" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-01-01" firstname="Henryk" gender="M" lastname="Zientara" nation="POL" athleteid="3617">
              <RESULTS>
                <RESULT eventid="1411" points="134" reactiontime="+107" swimtime="00:04:08.57" resultid="3619" lane="5" heatid="7003" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.49" />
                    <SPLIT distance="50" swimtime="00:00:50.65" />
                    <SPLIT distance="75" swimtime="00:01:20.72" />
                    <SPLIT distance="100" swimtime="00:01:52.85" />
                    <SPLIT distance="125" swimtime="00:02:26.07" />
                    <SPLIT distance="150" swimtime="00:03:00.22" />
                    <SPLIT distance="175" swimtime="00:03:34.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="146" reactiontime="+132" swimtime="00:01:51.64" resultid="3621" lane="5" heatid="7303" entrytime="00:01:54.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.24" />
                    <SPLIT distance="50" swimtime="00:00:51.17" />
                    <SPLIT distance="75" swimtime="00:01:21.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="84" reactiontime="+86" swimtime="00:01:59.61" resultid="3622" lane="1" heatid="7319" entrytime="00:02:04.21">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.45" />
                    <SPLIT distance="50" swimtime="00:00:56.42" />
                    <SPLIT distance="75" swimtime="00:01:28.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="176" reactiontime="+107" swimtime="00:00:48.42" resultid="3618" lane="5" heatid="6855" entrytime="00:00:49.17">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="106" reactiontime="+95" swimtime="00:00:51.69" resultid="3620" lane="6" heatid="7034" entrytime="00:00:49.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Jarosław" gender="M" lastname="Wysocki" nation="POL" athleteid="3623">
              <RESULTS>
                <RESULT eventid="1239" points="278" reactiontime="+84" swimtime="00:00:41.64" resultid="3625" lane="8" heatid="6858" entrytime="00:00:42.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="257" reactiontime="+86" swimtime="00:01:32.62" resultid="3627" heatid="7306" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.20" />
                    <SPLIT distance="50" swimtime="00:00:43.84" />
                    <SPLIT distance="75" swimtime="00:01:07.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="219" reactiontime="+86" swimtime="00:03:31.32" resultid="3626" lane="5" heatid="7005" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.05" />
                    <SPLIT distance="50" swimtime="00:00:46.62" />
                    <SPLIT distance="75" swimtime="00:01:13.29" />
                    <SPLIT distance="100" swimtime="00:01:40.72" />
                    <SPLIT distance="125" swimtime="00:02:09.38" />
                    <SPLIT distance="150" swimtime="00:02:36.73" />
                    <SPLIT distance="175" swimtime="00:03:04.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="163" reactiontime="+83" swimtime="00:01:33.51" resultid="3624" lane="4" heatid="6732" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.32" />
                    <SPLIT distance="50" swimtime="00:00:45.19" />
                    <SPLIT distance="75" swimtime="00:01:09.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-01" firstname="Krzysztof" gender="M" lastname="Lietz" nation="POL" athleteid="3628">
              <RESULTS>
                <RESULT eventid="1645" points="294" reactiontime="+76" swimtime="00:00:34.52" resultid="3634" lane="6" heatid="7286" entrytime="00:00:34.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="323" reactiontime="+78" swimtime="00:00:30.99" resultid="3635" lane="1" heatid="7342" entrytime="00:00:31.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="222" reactiontime="+79" swimtime="00:01:24.41" resultid="3629" lane="2" heatid="6736" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.99" />
                    <SPLIT distance="50" swimtime="00:00:40.36" />
                    <SPLIT distance="75" swimtime="00:01:05.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="195" reactiontime="+89" swimtime="00:03:16.68" resultid="3633" lane="4" heatid="7074" entrytime="00:03:19.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.19" />
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                    <SPLIT distance="75" swimtime="00:01:07.47" />
                    <SPLIT distance="100" swimtime="00:01:35.97" />
                    <SPLIT distance="125" swimtime="00:02:05.35" />
                    <SPLIT distance="150" swimtime="00:02:33.58" />
                    <SPLIT distance="175" swimtime="00:02:56.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="275" reactiontime="+76" swimtime="00:00:41.76" resultid="3631" lane="3" heatid="6858" entrytime="00:00:40.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="185" reactiontime="+86" swimtime="00:01:28.39" resultid="3632" lane="4" heatid="7017" entrytime="00:01:29.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.96" />
                    <SPLIT distance="50" swimtime="00:00:40.88" />
                    <SPLIT distance="75" swimtime="00:01:05.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="279" reactiontime="+78" swimtime="00:01:11.92" resultid="3630" lane="3" heatid="6835" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.98" />
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="75" swimtime="00:00:53.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-01" firstname="Marcin" gender="M" lastname="Mykowski" nation="POL" athleteid="3636">
              <RESULTS>
                <RESULT eventid="1205" points="568" reactiontime="+75" swimtime="00:00:56.81" resultid="3637" lane="6" heatid="6843" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.10" />
                    <SPLIT distance="50" swimtime="00:00:27.37" />
                    <SPLIT distance="75" swimtime="00:00:42.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="554" reactiontime="+73" swimtime="00:00:25.91" resultid="3639" lane="8" heatid="7351" entrytime="00:00:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" status="DNS" swimtime="00:00:00.00" resultid="3638" lane="7" heatid="7041" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-01" firstname="Grzegorz" gender="M" lastname="Arentewicz" nation="POL" athleteid="3640">
              <RESULTS>
                <RESULT eventid="1564" points="299" reactiontime="+81" swimtime="00:02:33.91" resultid="3645" lane="6" heatid="7062" entrytime="00:02:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.95" />
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                    <SPLIT distance="75" swimtime="00:00:52.17" />
                    <SPLIT distance="100" swimtime="00:01:11.42" />
                    <SPLIT distance="125" swimtime="00:02:14.65" />
                    <SPLIT distance="150" swimtime="00:01:53.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="309" reactiontime="+85" swimtime="00:01:14.51" resultid="3644" heatid="7020" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.53" />
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                    <SPLIT distance="75" swimtime="00:00:54.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="276" reactiontime="+85" swimtime="00:05:37.91" resultid="3643" lane="3" heatid="6905" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.93" />
                    <SPLIT distance="50" swimtime="00:00:36.04" />
                    <SPLIT distance="75" swimtime="00:00:55.88" />
                    <SPLIT distance="100" swimtime="00:01:17.13" />
                    <SPLIT distance="125" swimtime="00:02:20.38" />
                    <SPLIT distance="150" swimtime="00:01:59.35" />
                    <SPLIT distance="175" swimtime="00:03:04.49" />
                    <SPLIT distance="200" swimtime="00:02:42.47" />
                    <SPLIT distance="225" swimtime="00:03:48.64" />
                    <SPLIT distance="250" swimtime="00:03:26.74" />
                    <SPLIT distance="275" swimtime="00:04:33.05" />
                    <SPLIT distance="300" swimtime="00:04:10.87" />
                    <SPLIT distance="325" swimtime="00:05:16.84" />
                    <SPLIT distance="350" swimtime="00:04:54.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="348" reactiontime="+84" swimtime="00:01:06.85" resultid="3642" lane="2" heatid="6838" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.30" />
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                    <SPLIT distance="75" swimtime="00:00:49.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="356" reactiontime="+78" swimtime="00:00:32.37" resultid="3646" lane="7" heatid="7288" entrytime="00:00:32.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="274" reactiontime="+79" swimtime="00:01:18.73" resultid="3641" lane="2" heatid="6738" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.02" />
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                    <SPLIT distance="75" swimtime="00:01:00.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="364" reactiontime="+80" swimtime="00:00:29.78" resultid="3647" heatid="7345" entrytime="00:00:29.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-01" firstname="Artur" gender="M" lastname="Kłosiński" nation="POL" athleteid="3648">
              <RESULTS>
                <RESULT eventid="1564" points="442" reactiontime="+72" swimtime="00:02:15.14" resultid="3653" lane="1" heatid="7063" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.05" />
                    <SPLIT distance="50" swimtime="00:00:30.59" />
                    <SPLIT distance="75" swimtime="00:00:47.57" />
                    <SPLIT distance="100" swimtime="00:01:04.73" />
                    <SPLIT distance="125" swimtime="00:01:22.33" />
                    <SPLIT distance="150" swimtime="00:01:40.30" />
                    <SPLIT distance="175" swimtime="00:01:58.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="384" reactiontime="+68" swimtime="00:01:12.25" resultid="3654" heatid="7323" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.36" />
                    <SPLIT distance="50" swimtime="00:00:35.25" />
                    <SPLIT distance="75" swimtime="00:00:53.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="531" reactiontime="+79" swimtime="00:00:58.07" resultid="3650" lane="4" heatid="6844" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.15" />
                    <SPLIT distance="50" swimtime="00:00:27.74" />
                    <SPLIT distance="75" swimtime="00:00:42.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="407" reactiontime="+79" swimtime="00:01:09.02" resultid="3649" lane="5" heatid="6741" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.63" />
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                    <SPLIT distance="75" swimtime="00:00:52.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="531" reactiontime="+74" swimtime="00:00:26.27" resultid="3655" lane="8" heatid="7352" entrytime="00:00:26.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="453" reactiontime="+76" swimtime="00:00:35.38" resultid="3651" lane="5" heatid="6862" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" status="DNS" swimtime="00:00:00.00" resultid="3652" lane="5" heatid="7040" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-02-16" firstname="Agnieszka" gender="F" lastname="Kostyra" nation="POL" athleteid="3656">
              <RESULTS>
                <RESULT eventid="1058" points="323" swimtime="00:11:59.94" resultid="3657" lane="5" heatid="6715" entrytime="00:11:20.00" />
                <RESULT eventid="1358" points="341" reactiontime="+75" swimtime="00:05:45.71" resultid="3659" lane="1" heatid="6898" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.13" />
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                    <SPLIT distance="75" swimtime="00:00:55.86" />
                    <SPLIT distance="100" swimtime="00:01:16.13" />
                    <SPLIT distance="125" swimtime="00:01:36.80" />
                    <SPLIT distance="150" swimtime="00:01:57.81" />
                    <SPLIT distance="175" swimtime="00:02:19.48" />
                    <SPLIT distance="200" swimtime="00:02:41.73" />
                    <SPLIT distance="225" swimtime="00:03:04.33" />
                    <SPLIT distance="250" swimtime="00:03:27.18" />
                    <SPLIT distance="275" swimtime="00:03:50.56" />
                    <SPLIT distance="300" swimtime="00:04:13.40" />
                    <SPLIT distance="325" swimtime="00:04:36.78" />
                    <SPLIT distance="350" swimtime="00:05:00.45" />
                    <SPLIT distance="375" swimtime="00:05:23.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1581" points="352" reactiontime="+63" swimtime="00:03:01.85" resultid="3661" lane="4" heatid="7070" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.05" />
                    <SPLIT distance="50" swimtime="00:00:38.31" />
                    <SPLIT distance="75" swimtime="00:01:01.65" />
                    <SPLIT distance="100" swimtime="00:01:23.85" />
                    <SPLIT distance="125" swimtime="00:01:50.03" />
                    <SPLIT distance="150" swimtime="00:02:17.15" />
                    <SPLIT distance="175" swimtime="00:02:40.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1781" points="326" reactiontime="+70" swimtime="00:06:31.19" resultid="3663" lane="3" heatid="7356" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.78" />
                    <SPLIT distance="50" swimtime="00:00:44.54" />
                    <SPLIT distance="75" swimtime="00:01:10.18" />
                    <SPLIT distance="100" swimtime="00:01:38.01" />
                    <SPLIT distance="125" swimtime="00:02:02.72" />
                    <SPLIT distance="150" swimtime="00:02:26.37" />
                    <SPLIT distance="175" swimtime="00:02:50.42" />
                    <SPLIT distance="200" swimtime="00:03:13.85" />
                    <SPLIT distance="225" swimtime="00:03:41.94" />
                    <SPLIT distance="250" swimtime="00:04:09.23" />
                    <SPLIT distance="275" swimtime="00:04:35.18" />
                    <SPLIT distance="300" swimtime="00:05:01.74" />
                    <SPLIT distance="325" swimtime="00:05:25.26" />
                    <SPLIT distance="350" swimtime="00:05:47.36" />
                    <SPLIT distance="375" swimtime="00:06:09.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="353" reactiontime="+73" swimtime="00:02:42.41" resultid="3660" lane="1" heatid="7053" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.45" />
                    <SPLIT distance="50" swimtime="00:00:35.23" />
                    <SPLIT distance="75" swimtime="00:00:54.57" />
                    <SPLIT distance="100" swimtime="00:01:15.51" />
                    <SPLIT distance="125" swimtime="00:01:37.23" />
                    <SPLIT distance="150" swimtime="00:01:59.05" />
                    <SPLIT distance="175" swimtime="00:02:20.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="353" reactiontime="+75" swimtime="00:02:57.20" resultid="3658" lane="1" heatid="6879" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.80" />
                    <SPLIT distance="50" swimtime="00:00:42.29" />
                    <SPLIT distance="75" swimtime="00:01:04.22" />
                    <SPLIT distance="100" swimtime="00:01:26.75" />
                    <SPLIT distance="125" swimtime="00:01:49.08" />
                    <SPLIT distance="150" swimtime="00:02:11.94" />
                    <SPLIT distance="175" swimtime="00:02:34.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="321" reactiontime="+73" swimtime="00:00:37.17" resultid="3662" lane="8" heatid="7280" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-01" firstname="Magdalena" gender="F" lastname="Rogozińska" nation="POL" athleteid="3664">
              <RESULTS>
                <RESULT eventid="1092" points="367" swimtime="00:01:22.07" resultid="3665" lane="2" heatid="6728" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.87" />
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                    <SPLIT distance="75" swimtime="00:01:01.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="391" reactiontime="+90" swimtime="00:00:41.45" resultid="3666" lane="6" heatid="6852" entrytime="00:00:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1409" points="314" reactiontime="+94" swimtime="00:03:26.28" resultid="3667" lane="1" heatid="7000" entrytime="00:03:29.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.64" />
                    <SPLIT distance="50" swimtime="00:00:47.19" />
                    <SPLIT distance="75" swimtime="00:01:13.54" />
                    <SPLIT distance="100" swimtime="00:01:40.22" />
                    <SPLIT distance="125" swimtime="00:02:07.18" />
                    <SPLIT distance="150" swimtime="00:02:34.38" />
                    <SPLIT distance="175" swimtime="00:03:01.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="350" reactiontime="+90" swimtime="00:01:32.30" resultid="3670" lane="6" heatid="7300" entrytime="00:01:29.45">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.40" />
                    <SPLIT distance="50" swimtime="00:00:44.05" />
                    <SPLIT distance="75" swimtime="00:01:08.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="275" reactiontime="+95" swimtime="00:00:39.12" resultid="3669" lane="1" heatid="7278" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="345" reactiontime="+79" swimtime="00:00:39.42" resultid="3668" lane="6" heatid="7029" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-01" firstname="Maciej" gender="M" lastname="Kuras" nation="POL" athleteid="3671">
              <RESULTS>
                <RESULT eventid="1307" points="339" reactiontime="+74" swimtime="00:02:43.26" resultid="3673" lane="2" heatid="6885" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.16" />
                    <SPLIT distance="50" swimtime="00:00:38.22" />
                    <SPLIT distance="75" swimtime="00:00:58.81" />
                    <SPLIT distance="100" swimtime="00:01:19.74" />
                    <SPLIT distance="125" swimtime="00:01:40.93" />
                    <SPLIT distance="150" swimtime="00:02:01.89" />
                    <SPLIT distance="175" swimtime="00:02:22.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="338" reactiontime="+71" swimtime="00:01:15.39" resultid="3677" lane="1" heatid="7324" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.89" />
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                    <SPLIT distance="75" swimtime="00:00:55.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="320" reactiontime="+73" swimtime="00:02:46.87" resultid="3675" heatid="7078" entrytime="00:02:46.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.92" />
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                    <SPLIT distance="75" swimtime="00:00:54.73" />
                    <SPLIT distance="100" swimtime="00:01:15.41" />
                    <SPLIT distance="125" swimtime="00:01:39.67" />
                    <SPLIT distance="150" swimtime="00:02:04.70" />
                    <SPLIT distance="175" swimtime="00:02:26.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="422" reactiontime="+67" swimtime="00:00:30.61" resultid="3676" lane="5" heatid="7289" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="325" reactiontime="+67" swimtime="00:00:35.58" resultid="3674" lane="1" heatid="7038" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="338" reactiontime="+73" swimtime="00:01:13.38" resultid="3672" lane="1" heatid="6740" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.22" />
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                    <SPLIT distance="75" swimtime="00:00:54.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-07-06" firstname="Andrzej" gender="M" lastname="Szufarski" nation="POL" athleteid="3678">
              <RESULTS>
                <RESULT eventid="1645" points="168" reactiontime="+106" swimtime="00:00:41.55" resultid="3682" lane="8" heatid="7283" entrytime="00:00:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="189" reactiontime="+99" swimtime="00:01:42.50" resultid="3683" lane="5" heatid="7305" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.62" />
                    <SPLIT distance="50" swimtime="00:00:47.16" />
                    <SPLIT distance="75" swimtime="00:01:14.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="97" reactiontime="+109" swimtime="00:01:49.58" resultid="3681" lane="4" heatid="7016" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.11" />
                    <SPLIT distance="50" swimtime="00:00:45.13" />
                    <SPLIT distance="75" swimtime="00:01:13.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="203" reactiontime="+100" swimtime="00:00:46.24" resultid="3680" heatid="6857" entrytime="00:00:44.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="140" reactiontime="+102" swimtime="00:01:38.46" resultid="3679" lane="8" heatid="6733" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.43" />
                    <SPLIT distance="50" swimtime="00:00:46.16" />
                    <SPLIT distance="75" swimtime="00:01:14.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1177" points="480" reactiontime="+72" swimtime="00:01:50.77" resultid="3684" lane="3" heatid="6809" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.70" />
                    <SPLIT distance="50" swimtime="00:00:25.93" />
                    <SPLIT distance="75" swimtime="00:00:40.27" />
                    <SPLIT distance="100" swimtime="00:00:55.55" />
                    <SPLIT distance="125" swimtime="00:01:09.41" />
                    <SPLIT distance="150" swimtime="00:01:24.56" />
                    <SPLIT distance="175" swimtime="00:01:37.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3636" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="3640" number="2" reactiontime="+66" />
                    <RELAYPOSITION athleteid="3671" number="3" reactiontime="+31" />
                    <RELAYPOSITION athleteid="3648" number="4" reactiontime="+52" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1341" points="442" reactiontime="+62" swimtime="00:02:05.32" resultid="3685" lane="1" heatid="6987" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.23" />
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                    <SPLIT distance="75" swimtime="00:00:47.08" />
                    <SPLIT distance="100" swimtime="00:01:07.19" />
                    <SPLIT distance="125" swimtime="00:01:21.87" />
                    <SPLIT distance="150" swimtime="00:01:39.00" />
                    <SPLIT distance="175" swimtime="00:01:51.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3636" number="1" reactiontime="+62" />
                    <RELAYPOSITION athleteid="3640" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="3671" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="3648" number="4" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1341" points="173" reactiontime="+55" swimtime="00:02:51.11" resultid="3686" lane="8" heatid="6986" entrytime="00:02:46.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.53" />
                    <SPLIT distance="50" swimtime="00:00:52.34" />
                    <SPLIT distance="75" swimtime="00:01:12.14" />
                    <SPLIT distance="100" swimtime="00:01:35.36" />
                    <SPLIT distance="125" swimtime="00:01:50.94" />
                    <SPLIT distance="150" swimtime="00:02:28.02" />
                    <SPLIT distance="175" swimtime="00:02:27.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3678" number="1" reactiontime="+55" />
                    <RELAYPOSITION athleteid="3623" number="2" reactiontime="+20" />
                    <RELAYPOSITION athleteid="3628" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="3603" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="VIJOZ" name="UKS Victoria Józefów" nation="POL" region="WA">
          <CONTACT email="ali90@o2.pl" name="kowalczyk alicja" />
          <ATHLETES>
            <ATHLETE birthdate="1966-03-01" firstname="Jan" gender="M" lastname="Kośmider" nation="POL" athleteid="3699">
              <RESULTS>
                <RESULT eventid="1798" points="349" reactiontime="+90" swimtime="00:05:46.22" resultid="3705" lane="4" heatid="7363" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.96" />
                    <SPLIT distance="50" swimtime="00:00:37.11" />
                    <SPLIT distance="75" swimtime="00:00:58.42" />
                    <SPLIT distance="100" swimtime="00:01:20.78" />
                    <SPLIT distance="125" swimtime="00:01:45.04" />
                    <SPLIT distance="150" swimtime="00:02:07.99" />
                    <SPLIT distance="175" swimtime="00:02:30.14" />
                    <SPLIT distance="200" swimtime="00:02:52.10" />
                    <SPLIT distance="225" swimtime="00:03:15.69" />
                    <SPLIT distance="250" swimtime="00:03:39.61" />
                    <SPLIT distance="275" swimtime="00:04:04.22" />
                    <SPLIT distance="300" swimtime="00:04:28.41" />
                    <SPLIT distance="325" swimtime="00:04:49.60" />
                    <SPLIT distance="350" swimtime="00:05:09.68" />
                    <SPLIT distance="375" swimtime="00:05:28.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="399" swimtime="00:10:22.70" resultid="3700" lane="8" heatid="6722" entrytime="00:10:45.00" />
                <RESULT eventid="1375" points="427" reactiontime="+80" swimtime="00:04:52.17" resultid="3702" lane="1" heatid="6908" entrytime="00:04:54.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.07" />
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="75" swimtime="00:00:50.45" />
                    <SPLIT distance="100" swimtime="00:01:08.91" />
                    <SPLIT distance="125" swimtime="00:01:27.74" />
                    <SPLIT distance="150" swimtime="00:01:46.61" />
                    <SPLIT distance="175" swimtime="00:02:05.73" />
                    <SPLIT distance="200" swimtime="00:02:24.68" />
                    <SPLIT distance="225" swimtime="00:02:43.18" />
                    <SPLIT distance="250" swimtime="00:03:01.82" />
                    <SPLIT distance="275" swimtime="00:03:20.44" />
                    <SPLIT distance="300" swimtime="00:03:39.12" />
                    <SPLIT distance="325" swimtime="00:03:57.41" />
                    <SPLIT distance="350" swimtime="00:04:15.98" />
                    <SPLIT distance="375" swimtime="00:04:34.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="432" reactiontime="+79" swimtime="00:00:35.95" resultid="3701" lane="5" heatid="6863" entrytime="00:00:36.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="3703" lane="6" heatid="7064" entrytime="00:02:15.50" />
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="3704" lane="3" heatid="7288" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WOSIE" name="Wodnik Siemianowice Śląskie" nation="POL">
          <CONTACT name="Piotr Szymik" />
          <ATHLETES>
            <ATHLETE birthdate="1960-02-18" firstname="Piotr" gender="M" lastname="Szymik" nation="POL" athleteid="3707">
              <RESULTS>
                <RESULT eventid="1143" points="311" swimtime="00:21:29.63" resultid="3708" heatid="6752" entrytime="00:21:21.41" />
                <RESULT eventid="1462" points="217" reactiontime="+88" swimtime="00:01:23.85" resultid="3711" heatid="7019" entrytime="00:01:22.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.15" />
                    <SPLIT distance="50" swimtime="00:00:39.29" />
                    <SPLIT distance="75" swimtime="00:01:01.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="294" reactiontime="+74" swimtime="00:05:30.76" resultid="3710" lane="1" heatid="6906" entrytime="00:05:31.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.94" />
                    <SPLIT distance="50" swimtime="00:00:35.62" />
                    <SPLIT distance="75" swimtime="00:00:54.94" />
                    <SPLIT distance="100" swimtime="00:01:15.24" />
                    <SPLIT distance="125" swimtime="00:01:36.14" />
                    <SPLIT distance="150" swimtime="00:01:57.38" />
                    <SPLIT distance="175" swimtime="00:02:18.48" />
                    <SPLIT distance="200" swimtime="00:02:39.69" />
                    <SPLIT distance="225" swimtime="00:03:01.00" />
                    <SPLIT distance="250" swimtime="00:03:22.87" />
                    <SPLIT distance="275" swimtime="00:03:44.36" />
                    <SPLIT distance="300" swimtime="00:04:05.93" />
                    <SPLIT distance="325" swimtime="00:04:27.18" />
                    <SPLIT distance="350" swimtime="00:04:49.33" />
                    <SPLIT distance="375" swimtime="00:05:10.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="250" reactiontime="+77" swimtime="00:00:36.43" resultid="3713" lane="3" heatid="7284" entrytime="00:00:36.11">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="269" reactiontime="+85" swimtime="00:06:17.30" resultid="3714" lane="6" heatid="7362" entrytime="00:06:21.14">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.00" />
                    <SPLIT distance="50" swimtime="00:00:43.41" />
                    <SPLIT distance="75" swimtime="00:01:07.34" />
                    <SPLIT distance="100" swimtime="00:01:31.33" />
                    <SPLIT distance="125" swimtime="00:01:54.90" />
                    <SPLIT distance="150" swimtime="00:02:18.55" />
                    <SPLIT distance="175" swimtime="00:02:43.09" />
                    <SPLIT distance="200" swimtime="00:03:08.26" />
                    <SPLIT distance="225" swimtime="00:03:35.08" />
                    <SPLIT distance="250" swimtime="00:04:01.70" />
                    <SPLIT distance="275" swimtime="00:04:29.07" />
                    <SPLIT distance="300" swimtime="00:04:55.41" />
                    <SPLIT distance="325" swimtime="00:05:16.01" />
                    <SPLIT distance="350" swimtime="00:05:36.25" />
                    <SPLIT distance="375" swimtime="00:05:57.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="266" reactiontime="+89" swimtime="00:02:57.58" resultid="3712" heatid="7077" entrytime="00:02:55.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.81" />
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                    <SPLIT distance="75" swimtime="00:01:01.81" />
                    <SPLIT distance="100" swimtime="00:01:24.80" />
                    <SPLIT distance="125" swimtime="00:01:50.70" />
                    <SPLIT distance="150" swimtime="00:02:17.06" />
                    <SPLIT distance="175" swimtime="00:02:37.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="3709" lane="8" heatid="6872" entrytime="00:03:15.14" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TROBO" name="UKS Trojka Oborniki" nation="POL" region="WIE">
          <CONTACT city="OBORNIKI" email="jawol@poczta.onet.pl" name="WOLNIEWICZ" phone="791064667" state="WIE" street="PIŁSUDSKIEGO 49/42" zip="64-600" />
          <ATHLETES>
            <ATHLETE birthdate="1948-01-01" firstname="Janusz" gender="M" lastname="Wolniewicz" nation="POL" athleteid="3716">
              <RESULTS>
                <RESULT eventid="1143" points="149" swimtime="00:27:27.28" resultid="3717" lane="6" heatid="6749" entrytime="00:28:44.64" entrycourse="SCM" />
                <RESULT eventid="1564" points="160" reactiontime="+114" swimtime="00:03:09.51" resultid="3719" lane="7" heatid="7056" entrytime="00:03:14.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.87" />
                    <SPLIT distance="50" swimtime="00:00:40.29" />
                    <SPLIT distance="75" swimtime="00:01:03.80" />
                    <SPLIT distance="100" swimtime="00:01:27.69" />
                    <SPLIT distance="125" swimtime="00:01:53.05" />
                    <SPLIT distance="150" swimtime="00:02:19.04" />
                    <SPLIT distance="175" swimtime="00:02:45.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="158" reactiontime="+101" swimtime="00:06:46.52" resultid="3718" lane="6" heatid="6901" entrytime="00:06:50.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.86" />
                    <SPLIT distance="50" swimtime="00:00:44.16" />
                    <SPLIT distance="75" swimtime="00:01:08.39" />
                    <SPLIT distance="100" swimtime="00:01:33.01" />
                    <SPLIT distance="125" swimtime="00:01:58.27" />
                    <SPLIT distance="150" swimtime="00:02:23.99" />
                    <SPLIT distance="175" swimtime="00:02:49.96" />
                    <SPLIT distance="200" swimtime="00:03:16.26" />
                    <SPLIT distance="225" swimtime="00:03:42.60" />
                    <SPLIT distance="250" swimtime="00:04:09.09" />
                    <SPLIT distance="275" swimtime="00:04:35.81" />
                    <SPLIT distance="300" swimtime="00:05:02.25" />
                    <SPLIT distance="325" swimtime="00:05:29.27" />
                    <SPLIT distance="350" swimtime="00:05:55.66" />
                    <SPLIT distance="375" swimtime="00:06:21.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="81" reactiontime="+107" swimtime="00:09:21.70" resultid="3720" lane="5" heatid="7358" entrytime="00:08:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.74" />
                    <SPLIT distance="50" swimtime="00:01:00.81" />
                    <SPLIT distance="75" swimtime="00:01:36.25" />
                    <SPLIT distance="100" swimtime="00:02:13.61" />
                    <SPLIT distance="125" swimtime="00:04:08.57" />
                    <SPLIT distance="150" swimtime="00:03:31.14" />
                    <SPLIT distance="175" swimtime="00:05:28.82" />
                    <SPLIT distance="200" swimtime="00:04:45.41" />
                    <SPLIT distance="225" swimtime="00:06:54.14" />
                    <SPLIT distance="250" swimtime="00:06:12.11" />
                    <SPLIT distance="275" swimtime="00:08:03.11" />
                    <SPLIT distance="300" swimtime="00:07:36.78" />
                    <SPLIT distance="325" swimtime="00:08:56.17" />
                    <SPLIT distance="350" swimtime="00:08:29.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WOZGI" name="Zgiersko-Łęczycki Wopr" nation="POL" region="LOD">
          <CONTACT city="ZGIERZ" email="UJANIN@GMAIL.COM" name="JANISZEWSKA" phone="601326923" state="ŁÓDZK" street="ŻYTNIA 84" zip="95-100" />
          <ATHLETES>
            <ATHLETE birthdate="1964-01-23" firstname="Urszula" gender="F" lastname="Janiszewska" nation="POL" athleteid="3722">
              <RESULTS>
                <RESULT eventid="1126" points="161" swimtime="00:28:49.46" resultid="3723" lane="4" heatid="6746" entrytime="00:29:00.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAKRA" name="Masters Kraśnik" nation="POL" region="LBL">
          <CONTACT name="G.M" />
          <ATHLETES>
            <ATHLETE birthdate="1975-01-01" firstname="Marcin" gender="M" lastname="Mazurek" nation="POL" athleteid="3725">
              <RESULTS>
                <RESULT eventid="1375" points="203" reactiontime="+90" swimtime="00:06:14.15" resultid="3727" lane="2" heatid="6905" entrytime="00:05:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.85" />
                    <SPLIT distance="50" swimtime="00:00:39.21" />
                    <SPLIT distance="75" swimtime="00:01:00.62" />
                    <SPLIT distance="100" swimtime="00:01:23.28" />
                    <SPLIT distance="125" swimtime="00:01:46.46" />
                    <SPLIT distance="150" swimtime="00:02:09.91" />
                    <SPLIT distance="175" swimtime="00:02:33.66" />
                    <SPLIT distance="200" swimtime="00:02:57.39" />
                    <SPLIT distance="225" swimtime="00:03:21.54" />
                    <SPLIT distance="250" swimtime="00:03:46.15" />
                    <SPLIT distance="275" swimtime="00:04:10.53" />
                    <SPLIT distance="300" swimtime="00:04:35.76" />
                    <SPLIT distance="325" swimtime="00:05:00.63" />
                    <SPLIT distance="350" swimtime="00:05:26.10" />
                    <SPLIT distance="375" swimtime="00:05:51.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="235" reactiontime="+95" swimtime="00:01:16.23" resultid="3726" lane="4" heatid="6834" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.84" />
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                    <SPLIT distance="75" swimtime="00:00:56.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="3728" heatid="7060" entrytime="00:02:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Krzysztof" gender="M" lastname="Samonek" nation="POL" athleteid="3729">
              <RESULTS>
                <RESULT eventid="1307" points="137" reactiontime="+86" swimtime="00:03:40.52" resultid="3731" lane="5" heatid="6882" entrytime="00:03:44.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.45" />
                    <SPLIT distance="50" swimtime="00:00:49.08" />
                    <SPLIT distance="75" swimtime="00:01:16.34" />
                    <SPLIT distance="100" swimtime="00:01:44.70" />
                    <SPLIT distance="125" swimtime="00:02:13.39" />
                    <SPLIT distance="150" swimtime="00:02:42.76" />
                    <SPLIT distance="175" swimtime="00:03:12.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="169" reactiontime="+83" swimtime="00:00:44.23" resultid="3732" lane="8" heatid="7036" entrytime="00:00:44.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="146" reactiontime="+80" swimtime="00:01:39.77" resultid="3734" lane="7" heatid="7321" entrytime="00:01:39.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.77" />
                    <SPLIT distance="50" swimtime="00:00:47.08" />
                    <SPLIT distance="75" swimtime="00:01:14.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="125" reactiontime="+79" swimtime="00:00:45.88" resultid="3733" lane="1" heatid="7282" entrytime="00:00:45.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="125" reactiontime="+94" swimtime="00:01:42.20" resultid="3730" lane="7" heatid="6732" entrytime="00:01:40.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.70" />
                    <SPLIT distance="50" swimtime="00:00:46.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Ewa" gender="F" lastname="Białosiewicz" nation="POL" athleteid="3735">
              <RESULTS>
                <RESULT eventid="1290" points="117" reactiontime="+85" swimtime="00:04:15.46" resultid="3737" heatid="6877" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:31.22" />
                    <SPLIT distance="50" swimtime="00:01:02.86" />
                    <SPLIT distance="75" swimtime="00:01:35.45" />
                    <SPLIT distance="100" swimtime="00:02:08.14" />
                    <SPLIT distance="125" swimtime="00:02:40.90" />
                    <SPLIT distance="150" swimtime="00:03:12.94" />
                    <SPLIT distance="175" swimtime="00:03:45.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1058" points="180" swimtime="00:14:34.34" resultid="3736" lane="7" heatid="6714" entrytime="00:14:50.00" />
                <RESULT eventid="1713" points="108" reactiontime="+82" swimtime="00:02:03.37" resultid="3739" lane="1" heatid="7314" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.22" />
                    <SPLIT distance="50" swimtime="00:01:01.31" />
                    <SPLIT distance="75" swimtime="00:01:32.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="176" reactiontime="+97" swimtime="00:07:10.38" resultid="3738" lane="3" heatid="6895" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.63" />
                    <SPLIT distance="50" swimtime="00:00:49.32" />
                    <SPLIT distance="75" swimtime="00:01:15.85" />
                    <SPLIT distance="100" swimtime="00:01:42.46" />
                    <SPLIT distance="125" swimtime="00:02:09.76" />
                    <SPLIT distance="150" swimtime="00:02:36.67" />
                    <SPLIT distance="175" swimtime="00:03:04.00" />
                    <SPLIT distance="200" swimtime="00:03:31.34" />
                    <SPLIT distance="225" swimtime="00:03:58.76" />
                    <SPLIT distance="250" swimtime="00:04:26.24" />
                    <SPLIT distance="275" swimtime="00:04:53.75" />
                    <SPLIT distance="300" swimtime="00:05:21.09" />
                    <SPLIT distance="325" swimtime="00:05:48.62" />
                    <SPLIT distance="350" swimtime="00:06:16.04" />
                    <SPLIT distance="375" swimtime="00:06:43.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-01" firstname="Mirosław" gender="M" lastname="Leszczyński" nation="POL" athleteid="3740">
              <RESULTS>
                <RESULT eventid="1696" points="334" reactiontime="+94" swimtime="00:01:24.88" resultid="3743" lane="4" heatid="7308" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.45" />
                    <SPLIT distance="50" swimtime="00:00:39.97" />
                    <SPLIT distance="75" swimtime="00:01:02.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="316" reactiontime="+95" swimtime="00:03:07.18" resultid="3742" lane="3" heatid="7009" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.10" />
                    <SPLIT distance="50" swimtime="00:00:42.38" />
                    <SPLIT distance="75" swimtime="00:01:05.60" />
                    <SPLIT distance="100" swimtime="00:01:29.72" />
                    <SPLIT distance="125" swimtime="00:01:54.06" />
                    <SPLIT distance="150" swimtime="00:02:18.60" />
                    <SPLIT distance="175" swimtime="00:02:42.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="351" reactiontime="+93" swimtime="00:00:38.53" resultid="3741" lane="4" heatid="6860" entrytime="00:00:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-01" firstname="Bartłomiej" gender="M" lastname="Sieczyński" nation="POL" athleteid="3744">
              <RESULTS>
                <RESULT eventid="1375" points="317" reactiontime="+98" swimtime="00:05:22.53" resultid="3746" lane="3" heatid="6906" entrytime="00:05:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.64" />
                    <SPLIT distance="50" swimtime="00:00:35.77" />
                    <SPLIT distance="75" swimtime="00:00:54.49" />
                    <SPLIT distance="100" swimtime="00:01:14.16" />
                    <SPLIT distance="125" swimtime="00:01:34.12" />
                    <SPLIT distance="150" swimtime="00:01:54.33" />
                    <SPLIT distance="175" swimtime="00:02:14.87" />
                    <SPLIT distance="200" swimtime="00:02:35.47" />
                    <SPLIT distance="225" swimtime="00:02:56.23" />
                    <SPLIT distance="250" swimtime="00:03:17.11" />
                    <SPLIT distance="275" swimtime="00:03:37.93" />
                    <SPLIT distance="300" swimtime="00:03:58.75" />
                    <SPLIT distance="325" swimtime="00:04:19.42" />
                    <SPLIT distance="350" swimtime="00:04:40.53" />
                    <SPLIT distance="375" swimtime="00:05:01.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="295" reactiontime="+86" swimtime="00:01:10.65" resultid="3745" heatid="6836" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.41" />
                    <SPLIT distance="50" swimtime="00:00:33.93" />
                    <SPLIT distance="75" swimtime="00:00:52.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="237" reactiontime="+82" swimtime="00:00:37.06" resultid="3749" lane="7" heatid="7284" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="3748" lane="7" heatid="7061" entrytime="00:02:35.00" />
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="3750" lane="5" heatid="7341" entrytime="00:00:32.00" />
                <RESULT eventid="1462" status="DNS" swimtime="00:00:00.00" resultid="3747" lane="6" heatid="7017" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Waldemar" gender="M" lastname="Rusowicz" nation="POL" athleteid="3751">
              <RESULTS>
                <RESULT eventid="1496" points="100" reactiontime="+90" swimtime="00:00:52.66" resultid="3755" lane="6" heatid="7035" entrytime="00:00:46.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="100" reactiontime="+97" swimtime="00:00:49.44" resultid="3757" lane="7" heatid="7282" entrytime="00:00:46.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="123" reactiontime="+95" swimtime="00:03:49.28" resultid="3756" lane="7" heatid="7073" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.49" />
                    <SPLIT distance="50" swimtime="00:00:52.50" />
                    <SPLIT distance="75" swimtime="00:01:24.87" />
                    <SPLIT distance="100" swimtime="00:01:55.76" />
                    <SPLIT distance="125" swimtime="00:02:26.76" />
                    <SPLIT distance="150" swimtime="00:02:56.83" />
                    <SPLIT distance="175" swimtime="00:03:24.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="207" reactiontime="+94" swimtime="00:00:45.91" resultid="3753" lane="5" heatid="6856" entrytime="00:00:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="187" reactiontime="+91" swimtime="00:01:43.00" resultid="3758" lane="8" heatid="7305" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.38" />
                    <SPLIT distance="50" swimtime="00:00:48.81" />
                    <SPLIT distance="75" swimtime="00:01:16.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="123" reactiontime="+99" swimtime="00:07:21.63" resultid="3754" lane="8" heatid="6901" entrytime="00:07:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.93" />
                    <SPLIT distance="50" swimtime="00:00:47.48" />
                    <SPLIT distance="75" swimtime="00:01:13.71" />
                    <SPLIT distance="100" swimtime="00:01:40.73" />
                    <SPLIT distance="125" swimtime="00:02:08.78" />
                    <SPLIT distance="150" swimtime="00:02:36.74" />
                    <SPLIT distance="175" swimtime="00:03:04.75" />
                    <SPLIT distance="200" swimtime="00:03:33.31" />
                    <SPLIT distance="225" swimtime="00:04:02.57" />
                    <SPLIT distance="250" swimtime="00:04:31.08" />
                    <SPLIT distance="275" swimtime="00:05:00.56" />
                    <SPLIT distance="300" swimtime="00:05:29.79" />
                    <SPLIT distance="325" swimtime="00:05:58.26" />
                    <SPLIT distance="350" swimtime="00:06:26.28" />
                    <SPLIT distance="375" swimtime="00:06:55.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="122" reactiontime="+87" swimtime="00:01:43.11" resultid="3752" lane="4" heatid="6731" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.33" />
                    <SPLIT distance="50" swimtime="00:00:52.23" />
                    <SPLIT distance="75" swimtime="00:01:19.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Janusz" gender="M" lastname="Wasiuk" nation="POL" athleteid="3759">
              <RESULTS>
                <RESULT eventid="1143" status="DNS" swimtime="00:00:00.00" resultid="3760" lane="4" heatid="6748" entrytime="00:33:00.00" />
                <RESULT eventid="1696" status="DNS" swimtime="00:00:00.00" resultid="3765" lane="4" heatid="7303" entrytime="00:01:50.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1341" points="247" reactiontime="+83" swimtime="00:02:32.15" resultid="6980" lane="6" heatid="6985">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:01:02.00" />
                    <SPLIT distance="50" swimtime="00:00:44.59" />
                    <SPLIT distance="75" swimtime="00:01:40.02" />
                    <SPLIT distance="100" swimtime="00:01:22.75" />
                    <SPLIT distance="125" swimtime="00:02:15.63" />
                    <SPLIT distance="150" swimtime="00:02:00.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3729" number="1" reactiontime="+83" />
                    <RELAYPOSITION athleteid="3740" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="3744" number="3" reactiontime="+64" />
                    <RELAYPOSITION athleteid="3725" number="4" reactiontime="+67" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="AZPOZ" name="AZS UAM Poznań" nation="POL">
          <ATHLETES>
            <ATHLETE birthdate="1986-01-01" firstname="Bartosz" gender="M" lastname="Ziemniarski" nation="POL" athleteid="3768">
              <RESULTS>
                <RESULT comment="Rekord Polski " eventid="1205" points="737" reactiontime="+77" swimtime="00:00:52.08" resultid="3769" lane="2" heatid="6846" entrytime="00:00:54.39">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.77" />
                    <SPLIT distance="50" swimtime="00:00:24.72" />
                    <SPLIT distance="75" swimtime="00:00:38.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="719" reactiontime="+74" swimtime="00:00:23.75" resultid="3771" lane="5" heatid="7354" entrytime="00:00:24.39">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="655" reactiontime="+78" swimtime="00:01:58.53" resultid="3770" lane="1" heatid="7066" entrytime="00:02:03.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.68" />
                    <SPLIT distance="50" swimtime="00:00:27.14" />
                    <SPLIT distance="75" swimtime="00:00:41.93" />
                    <SPLIT distance="100" swimtime="00:00:57.10" />
                    <SPLIT distance="125" swimtime="00:01:12.33" />
                    <SPLIT distance="150" swimtime="00:01:27.92" />
                    <SPLIT distance="175" swimtime="00:01:43.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Jakub" gender="M" lastname="Sterczyński" nation="POL" athleteid="3772">
              <RESULTS>
                <RESULT eventid="1798" points="494" reactiontime="+72" swimtime="00:05:08.30" resultid="3775" lane="3" heatid="7364" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.76" />
                    <SPLIT distance="50" swimtime="00:00:30.23" />
                    <SPLIT distance="75" swimtime="00:00:47.30" />
                    <SPLIT distance="100" swimtime="00:01:05.08" />
                    <SPLIT distance="125" swimtime="00:01:25.74" />
                    <SPLIT distance="150" swimtime="00:01:45.37" />
                    <SPLIT distance="175" swimtime="00:02:05.84" />
                    <SPLIT distance="200" swimtime="00:02:25.82" />
                    <SPLIT distance="225" swimtime="00:02:47.03" />
                    <SPLIT distance="250" swimtime="00:03:08.68" />
                    <SPLIT distance="275" swimtime="00:03:30.63" />
                    <SPLIT distance="300" swimtime="00:03:52.89" />
                    <SPLIT distance="325" swimtime="00:04:12.51" />
                    <SPLIT distance="350" swimtime="00:04:31.49" />
                    <SPLIT distance="375" swimtime="00:04:50.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="523" reactiontime="+75" swimtime="00:02:21.75" resultid="3774" lane="3" heatid="7080" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.53" />
                    <SPLIT distance="50" swimtime="00:00:29.56" />
                    <SPLIT distance="75" swimtime="00:00:48.55" />
                    <SPLIT distance="100" swimtime="00:01:05.94" />
                    <SPLIT distance="125" swimtime="00:01:26.09" />
                    <SPLIT distance="150" swimtime="00:01:46.72" />
                    <SPLIT distance="175" swimtime="00:02:04.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="498" swimtime="00:01:04.49" resultid="3773" lane="6" heatid="6745" entrytime="00:01:02.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-01" firstname="Michał" gender="M" lastname="Kamiński" nation="POL" athleteid="3776">
              <RESULTS>
                <RESULT eventid="1109" points="529" swimtime="00:01:03.23" resultid="3777" lane="2" heatid="6745" entrytime="00:01:01.00" />
                <RESULT eventid="1205" points="605" reactiontime="+76" swimtime="00:00:55.60" resultid="3778" lane="6" heatid="6846" entrytime="00:00:54.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.66" />
                    <SPLIT distance="50" swimtime="00:00:26.85" />
                    <SPLIT distance="75" swimtime="00:00:41.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-01" firstname="Jan" gender="M" lastname="Bręczewski" nation="POL" athleteid="3780">
              <RESULTS>
                <RESULT eventid="1645" points="507" reactiontime="+73" swimtime="00:00:28.79" resultid="3782" lane="4" heatid="7293" entrytime="00:00:27.01">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="567" reactiontime="+72" swimtime="00:00:25.71" resultid="3783" lane="8" heatid="7354" entrytime="00:00:25.01">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-01" firstname="Juliusz" gender="M" lastname="Żebrowski" nation="POL" athleteid="3784">
              <RESULTS>
                <RESULT eventid="1411" points="522" reactiontime="+66" swimtime="00:02:38.28" resultid="3787" lane="6" heatid="7011" entrytime="00:02:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.76" />
                    <SPLIT distance="50" swimtime="00:00:34.35" />
                    <SPLIT distance="75" swimtime="00:00:54.26" />
                    <SPLIT distance="100" swimtime="00:01:14.95" />
                    <SPLIT distance="125" swimtime="00:01:35.82" />
                    <SPLIT distance="150" swimtime="00:01:57.36" />
                    <SPLIT distance="175" swimtime="00:02:17.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="570" reactiontime="+67" swimtime="00:01:11.04" resultid="3788" heatid="7311" entrytime="00:01:12.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.02" />
                    <SPLIT distance="50" swimtime="00:00:32.84" />
                    <SPLIT distance="75" swimtime="00:00:51.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="462" reactiontime="+66" swimtime="00:01:06.16" resultid="3785" lane="8" heatid="6742" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.59" />
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                    <SPLIT distance="75" swimtime="00:00:49.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="543" reactiontime="+65" swimtime="00:00:26.07" resultid="3789" lane="7" heatid="7352" entrytime="00:00:26.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.84" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="07" eventid="1239" reactiontime="+66" status="DSQ" swimtime="00:00:31.83" resultid="3786" lane="4" heatid="6865" entrytime="00:00:32.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-01" firstname="Piotr" gender="M" lastname="Kowalik" nation="POL" athleteid="3790">
              <RESULTS>
                <RESULT eventid="1764" points="674" reactiontime="+66" swimtime="00:00:24.26" resultid="7491" lane="1" heatid="7354">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="762" reactiontime="+64" swimtime="00:00:25.13" resultid="3792" lane="3" heatid="7294" entrytime="00:00:25.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="695" reactiontime="+67" swimtime="00:00:56.89" resultid="3791" lane="3" heatid="7023" entrytime="00:00:56.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.43" />
                    <SPLIT distance="50" swimtime="00:00:25.40" />
                    <SPLIT distance="75" swimtime="00:00:40.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="96" agemin="80" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1177" points="680" reactiontime="+76" swimtime="00:01:38.64" resultid="3793" lane="3" heatid="6810" bonus="yes" entrytime="00:01:41.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.28" />
                    <SPLIT distance="50" swimtime="00:00:25.21" />
                    <SPLIT distance="75" swimtime="00:00:37.70" />
                    <SPLIT distance="100" swimtime="00:00:51.34" />
                    <SPLIT distance="125" swimtime="00:01:03.37" />
                    <SPLIT distance="150" swimtime="00:01:19.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3776" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="3772" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="3790" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="3768" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1341" points="675" reactiontime="+61" swimtime="00:01:48.84" resultid="3794" lane="3" heatid="6988" entrytime="00:01:53.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.86" />
                    <SPLIT distance="50" swimtime="00:00:27.97" />
                    <SPLIT distance="75" swimtime="00:00:41.87" />
                    <SPLIT distance="100" swimtime="00:00:58.99" />
                    <SPLIT distance="125" swimtime="00:01:11.02" />
                    <SPLIT distance="150" swimtime="00:01:25.69" />
                    <SPLIT distance="175" swimtime="00:01:36.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3790" number="1" reactiontime="+61" />
                    <RELAYPOSITION athleteid="3784" number="2" reactiontime="+12" />
                    <RELAYPOSITION athleteid="3776" number="3" reactiontime="+28" />
                    <RELAYPOSITION athleteid="3768" number="4" reactiontime="+11" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="319" agemin="280" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1615" status="DNS" swimtime="00:00:00.00" resultid="6664" lane="6" heatid="7441" entrytime="00:04:21.70">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4085" number="1" />
                    <RELAYPOSITION athleteid="4091" number="2" />
                    <RELAYPOSITION athleteid="4114" number="3" />
                    <RELAYPOSITION athleteid="4122" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1815" status="DNS" swimtime="00:00:00.00" resultid="6665" lane="4" heatid="7502" entrytime="00:05:11.80">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4085" number="1" />
                    <RELAYPOSITION athleteid="4091" number="2" />
                    <RELAYPOSITION athleteid="4114" number="3" />
                    <RELAYPOSITION athleteid="4122" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="AZKRA" name="AZS WSZIB Kraków" nation="POL">
          <CONTACT name="Palmowska" />
          <ATHLETES>
            <ATHLETE birthdate="1985-01-01" firstname="Paulina" gender="F" lastname="Palmowska" nation="POL" athleteid="3803">
              <RESULTS>
                <RESULT eventid="1290" points="448" reactiontime="+70" swimtime="00:02:43.65" resultid="3805" lane="5" heatid="6879" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.25" />
                    <SPLIT distance="50" swimtime="00:00:37.89" />
                    <SPLIT distance="75" swimtime="00:00:58.08" />
                    <SPLIT distance="100" swimtime="00:01:18.86" />
                    <SPLIT distance="125" swimtime="00:01:40.28" />
                    <SPLIT distance="150" swimtime="00:02:02.02" />
                    <SPLIT distance="175" swimtime="00:02:23.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="486" reactiontime="+67" swimtime="00:01:14.70" resultid="3807" lane="3" heatid="7317" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.50" />
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                    <SPLIT distance="75" swimtime="00:00:55.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="530" reactiontime="+66" swimtime="00:00:34.17" resultid="3806" lane="3" heatid="7031" entrytime="00:00:33.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="435" reactiontime="+68" swimtime="00:01:17.58" resultid="3804" lane="5" heatid="6729" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.78" />
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                    <SPLIT distance="75" swimtime="00:00:58.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="461" reactiontime="+69" swimtime="00:00:31.02" resultid="3808" lane="2" heatid="7335" entrytime="00:00:29.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Kamil" gender="M" lastname="Latuszek" nation="POL" athleteid="3809">
              <RESULTS>
                <RESULT eventid="1564" points="325" reactiontime="+75" swimtime="00:02:29.70" resultid="3811" lane="7" heatid="7064" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.54" />
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                    <SPLIT distance="75" swimtime="00:00:51.82" />
                    <SPLIT distance="100" swimtime="00:01:10.90" />
                    <SPLIT distance="125" swimtime="00:01:30.01" />
                    <SPLIT distance="150" swimtime="00:01:49.80" />
                    <SPLIT distance="175" swimtime="00:02:10.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="557" reactiontime="+73" swimtime="00:00:25.85" resultid="3812" lane="1" heatid="7353" entrytime="00:00:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="508" reactiontime="+76" swimtime="00:00:58.94" resultid="3810" lane="3" heatid="6844" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.84" />
                    <SPLIT distance="50" swimtime="00:00:27.21" />
                    <SPLIT distance="75" swimtime="00:00:42.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Konrad" gender="M" lastname="Latuszek" nation="POL" athleteid="3813">
              <RESULTS>
                <RESULT eventid="1239" points="543" reactiontime="+77" swimtime="00:00:33.30" resultid="3815" lane="4" heatid="6862" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="495" reactiontime="+75" swimtime="00:01:14.47" resultid="3819" lane="6" heatid="7310" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.77" />
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                    <SPLIT distance="75" swimtime="00:00:54.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="458" reactiontime="+82" swimtime="00:01:06.34" resultid="3814" lane="3" heatid="6743" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.20" />
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                    <SPLIT distance="75" swimtime="00:00:49.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" status="DNS" swimtime="00:00:00.00" resultid="3817" lane="1" heatid="7080" entrytime="00:02:25.00" />
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="3818" lane="3" heatid="7291" entrytime="00:00:29.00" />
                <RESULT comment="K 3" eventid="1411" reactiontime="+77" status="DSQ" swimtime="00:00:00.00" resultid="3816" lane="4" heatid="7010" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.54" />
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                    <SPLIT distance="75" swimtime="00:00:57.28" />
                    <SPLIT distance="100" swimtime="00:01:18.60" />
                    <SPLIT distance="125" swimtime="00:01:39.90" />
                    <SPLIT distance="150" swimtime="00:02:01.22" />
                    <SPLIT distance="175" swimtime="00:02:22.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KOOLS" name="Kormoran Olsztyn" nation="POL">
          <CONTACT name="Goździejewska" />
          <ATHLETES>
            <ATHLETE birthdate="1967-01-01" firstname="Anna" gender="F" lastname="Goździejewska" nation="POL" athleteid="3821">
              <RESULTS>
                <RESULT eventid="1781" points="275" reactiontime="+87" swimtime="00:06:54.03" resultid="3827" lane="2" heatid="7356" entrytime="00:06:48.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.06" />
                    <SPLIT distance="50" swimtime="00:00:47.51" />
                    <SPLIT distance="75" swimtime="00:01:13.49" />
                    <SPLIT distance="100" swimtime="00:01:41.36" />
                    <SPLIT distance="125" swimtime="00:02:08.10" />
                    <SPLIT distance="150" swimtime="00:02:35.34" />
                    <SPLIT distance="175" swimtime="00:03:01.71" />
                    <SPLIT distance="200" swimtime="00:03:27.52" />
                    <SPLIT distance="225" swimtime="00:03:55.20" />
                    <SPLIT distance="250" swimtime="00:04:22.79" />
                    <SPLIT distance="275" swimtime="00:04:50.87" />
                    <SPLIT distance="300" swimtime="00:05:18.99" />
                    <SPLIT distance="325" swimtime="00:05:42.73" />
                    <SPLIT distance="350" swimtime="00:06:08.06" />
                    <SPLIT distance="375" swimtime="00:06:31.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="314" reactiontime="+88" swimtime="00:02:48.86" resultid="3825" lane="7" heatid="7052" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.66" />
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                    <SPLIT distance="75" swimtime="00:00:58.32" />
                    <SPLIT distance="100" swimtime="00:01:19.46" />
                    <SPLIT distance="125" swimtime="00:01:41.34" />
                    <SPLIT distance="150" swimtime="00:02:03.83" />
                    <SPLIT distance="175" swimtime="00:02:26.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1409" points="306" reactiontime="+84" swimtime="00:03:28.06" resultid="3824" lane="2" heatid="7000" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.89" />
                    <SPLIT distance="50" swimtime="00:00:47.51" />
                    <SPLIT distance="75" swimtime="00:01:13.69" />
                    <SPLIT distance="100" swimtime="00:01:40.03" />
                    <SPLIT distance="125" swimtime="00:02:06.64" />
                    <SPLIT distance="150" swimtime="00:02:33.81" />
                    <SPLIT distance="175" swimtime="00:03:01.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="318" reactiontime="+84" swimtime="00:05:53.85" resultid="3823" lane="1" heatid="6897" entrytime="00:05:49.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.04" />
                    <SPLIT distance="50" swimtime="00:00:39.02" />
                    <SPLIT distance="75" swimtime="00:01:00.15" />
                    <SPLIT distance="100" swimtime="00:01:21.73" />
                    <SPLIT distance="125" swimtime="00:01:43.87" />
                    <SPLIT distance="150" swimtime="00:02:06.45" />
                    <SPLIT distance="175" swimtime="00:02:28.58" />
                    <SPLIT distance="200" swimtime="00:02:51.54" />
                    <SPLIT distance="225" swimtime="00:03:13.94" />
                    <SPLIT distance="250" swimtime="00:03:37.02" />
                    <SPLIT distance="275" swimtime="00:04:00.12" />
                    <SPLIT distance="300" swimtime="00:04:23.04" />
                    <SPLIT distance="325" swimtime="00:04:46.16" />
                    <SPLIT distance="350" swimtime="00:05:08.96" />
                    <SPLIT distance="375" swimtime="00:05:31.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1126" points="334" swimtime="00:22:37.86" resultid="3822" lane="5" heatid="6747" entrytime="00:22:50.00" />
                <RESULT eventid="1679" points="299" reactiontime="+84" swimtime="00:01:37.29" resultid="3826" lane="3" heatid="7299" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.32" />
                    <SPLIT distance="50" swimtime="00:00:46.10" />
                    <SPLIT distance="75" swimtime="00:01:11.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KOSZA" name="Koszalin" nation="POL">
          <CONTACT name="Michałkowski" />
          <ATHLETES>
            <ATHLETE birthdate="1951-01-01" firstname="Andrzej" gender="M" lastname="Michałkowski" nation="POL" athleteid="3829">
              <RESULTS>
                <RESULT eventid="1239" points="245" reactiontime="+104" swimtime="00:00:43.38" resultid="3832" lane="6" heatid="6858" entrytime="00:00:41.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="216" reactiontime="+110" swimtime="00:01:38.07" resultid="3835" lane="6" heatid="7305" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.89" />
                    <SPLIT distance="50" swimtime="00:00:45.91" />
                    <SPLIT distance="75" swimtime="00:01:11.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="102" reactiontime="+110" swimtime="00:01:49.37" resultid="3830" lane="8" heatid="6731" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.66" />
                    <SPLIT distance="50" swimtime="00:00:56.83" />
                    <SPLIT distance="75" swimtime="00:01:24.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="148" reactiontime="+103" swimtime="00:01:28.90" resultid="3831" lane="5" heatid="6831" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.56" />
                    <SPLIT distance="50" swimtime="00:00:40.65" />
                    <SPLIT distance="75" swimtime="00:01:04.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="178" reactiontime="+116" swimtime="00:03:46.35" resultid="3833" lane="8" heatid="7005" entrytime="00:03:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.60" />
                    <SPLIT distance="50" swimtime="00:00:48.23" />
                    <SPLIT distance="75" swimtime="00:01:15.92" />
                    <SPLIT distance="100" swimtime="00:01:44.63" />
                    <SPLIT distance="125" swimtime="00:02:13.69" />
                    <SPLIT distance="150" swimtime="00:02:41.90" />
                    <SPLIT distance="175" swimtime="00:03:16.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="170" reactiontime="+106" swimtime="00:00:38.34" resultid="3836" lane="5" heatid="7337" entrytime="00:00:38.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="3834" lane="5" heatid="7055" entrytime="00:03:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-01" firstname="Marek" gender="M" lastname="Michałkowski" nation="POL" athleteid="3837">
              <RESULTS>
                <RESULT eventid="1696" points="684" reactiontime="+62" swimtime="00:01:06.85" resultid="3842" lane="3" heatid="7311" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.30" />
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                    <SPLIT distance="75" swimtime="00:00:49.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="709" reactiontime="+65" swimtime="00:00:30.47" resultid="3840" lane="6" heatid="6866" entrytime="00:00:31.26">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="619" reactiontime="+65" swimtime="00:00:55.19" resultid="3839" lane="8" heatid="6846" entrytime="00:00:57.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.46" />
                    <SPLIT distance="50" swimtime="00:00:26.52" />
                    <SPLIT distance="75" swimtime="00:00:41.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="544" swimtime="00:01:02.65" resultid="3838" heatid="6745" entrytime="00:01:04.00" />
                <RESULT eventid="1496" points="434" reactiontime="+84" swimtime="00:00:32.31" resultid="3841" lane="6" heatid="7043" entrytime="00:00:29.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="621" reactiontime="+65" swimtime="00:00:24.94" resultid="3843" lane="3" heatid="7352" entrytime="00:00:26.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LEWAR" name="Legia Warszawa" nation="POL">
          <CONTACT name="Drzewiński" />
          <ATHLETES>
            <ATHLETE birthdate="1981-01-01" firstname="Marcin" gender="M" lastname="Wilczęga" nation="POL" athleteid="3845">
              <RESULTS>
                <RESULT eventid="1109" points="409" reactiontime="+69" swimtime="00:01:08.90" resultid="3846" lane="6" heatid="6742" entrytime="00:01:09.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.61" />
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                    <SPLIT distance="75" swimtime="00:00:51.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="532" reactiontime="+67" swimtime="00:00:26.25" resultid="3847" lane="5" heatid="7352" entrytime="00:00:26.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-01" firstname="Maciej" gender="M" lastname="Bień" nation="POL" athleteid="3848">
              <RESULTS>
                <RESULT eventid="1239" points="408" reactiontime="+85" swimtime="00:00:36.62" resultid="3850" heatid="6864" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="273" reactiontime="+91" swimtime="00:01:18.83" resultid="3849" lane="5" heatid="6737" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.55" />
                    <SPLIT distance="50" swimtime="00:00:38.20" />
                    <SPLIT distance="75" swimtime="00:01:00.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" status="DNS" swimtime="00:00:00.00" resultid="3852" lane="2" heatid="7009" entrytime="00:03:06.00" />
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="3853" lane="8" heatid="7062" entrytime="00:02:30.00" />
                <RESULT eventid="1696" status="DNS" swimtime="00:00:00.00" resultid="3854" lane="3" heatid="7308" entrytime="00:01:25.00" />
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="3855" lane="2" heatid="7345" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-01-01" firstname="Piotr" gender="M" lastname="Fuliński" nation="POL" athleteid="3856">
              <RESULTS>
                <RESULT eventid="1764" points="518" reactiontime="+94" swimtime="00:00:26.48" resultid="3857" heatid="7353" entrytime="00:00:26.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-01-01" firstname="Maciej" gender="M" lastname="Grzelak" nation="POL" athleteid="3858">
              <RESULTS>
                <RESULT eventid="1598" points="218" reactiontime="+77" swimtime="00:03:09.78" resultid="3863" heatid="7076" entrytime="00:03:06.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.19" />
                    <SPLIT distance="50" swimtime="00:00:34.55" />
                    <SPLIT distance="75" swimtime="00:01:03.15" />
                    <SPLIT distance="100" swimtime="00:01:32.27" />
                    <SPLIT distance="125" swimtime="00:01:58.70" />
                    <SPLIT distance="150" swimtime="00:02:26.06" />
                    <SPLIT distance="175" swimtime="00:02:48.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="254" reactiontime="+85" swimtime="00:01:19.54" resultid="3862" lane="5" heatid="7019" entrytime="00:01:18.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.30" />
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                    <SPLIT distance="75" swimtime="00:00:55.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="253" reactiontime="+68" swimtime="00:01:20.80" resultid="3859" lane="5" heatid="6736" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.98" />
                    <SPLIT distance="50" swimtime="00:00:38.11" />
                    <SPLIT distance="75" swimtime="00:01:01.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="343" reactiontime="+76" swimtime="00:00:38.82" resultid="3861" lane="1" heatid="6862" entrytime="00:00:37.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="201" reactiontime="+97" swimtime="00:06:56.11" resultid="3865" lane="7" heatid="7359" entrytime="00:07:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.04" />
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                    <SPLIT distance="75" swimtime="00:00:59.20" />
                    <SPLIT distance="100" swimtime="00:01:25.12" />
                    <SPLIT distance="125" swimtime="00:01:55.94" />
                    <SPLIT distance="150" swimtime="00:02:27.65" />
                    <SPLIT distance="175" swimtime="00:02:58.00" />
                    <SPLIT distance="200" swimtime="00:03:28.40" />
                    <SPLIT distance="225" swimtime="00:03:56.85" />
                    <SPLIT distance="250" swimtime="00:04:25.40" />
                    <SPLIT distance="275" swimtime="00:04:53.68" />
                    <SPLIT distance="300" swimtime="00:05:22.87" />
                    <SPLIT distance="325" swimtime="00:05:46.25" />
                    <SPLIT distance="350" swimtime="00:06:10.68" />
                    <SPLIT distance="375" swimtime="00:06:34.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="259" reactiontime="+86" swimtime="00:01:13.77" resultid="3860" lane="2" heatid="6840" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.04" />
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                    <SPLIT distance="75" swimtime="00:00:53.72" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="04" eventid="1696" reactiontime="+42" status="DSQ" swimtime="00:00:00.00" resultid="3864" lane="4" heatid="7306" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.63" />
                    <SPLIT distance="50" swimtime="00:00:42.06" />
                    <SPLIT distance="75" swimtime="00:01:05.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Krzesimir" gender="M" lastname="Sieczych" nation="POL" athleteid="3866">
              <RESULTS>
                <RESULT eventid="1205" points="426" reactiontime="+72" swimtime="00:01:02.53" resultid="3868" lane="1" heatid="6845" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.76" />
                    <SPLIT distance="50" swimtime="00:00:29.38" />
                    <SPLIT distance="75" swimtime="00:00:45.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="474" reactiontime="+79" swimtime="00:00:27.29" resultid="3870" lane="8" heatid="7353" entrytime="00:00:26.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="326" reactiontime="+75" swimtime="00:01:14.29" resultid="3867" lane="2" heatid="6742" entrytime="00:01:09.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.04" />
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                    <SPLIT distance="75" swimtime="00:00:56.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="422" reactiontime="+71" swimtime="00:00:30.60" resultid="3869" lane="8" heatid="7292" entrytime="00:00:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-01" firstname="Łukasz" gender="M" lastname="Drzewiński" nation="POL" athleteid="3871">
              <RESULTS>
                <RESULT eventid="1462" points="649" reactiontime="+75" swimtime="00:00:58.20" resultid="3874" lane="5" heatid="7023" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.31" />
                    <SPLIT distance="50" swimtime="00:00:27.09" />
                    <SPLIT distance="75" swimtime="00:00:42.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="560" reactiontime="+77" swimtime="00:02:15.91" resultid="3873" lane="5" heatid="6874" entrytime="00:02:16.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.82" />
                    <SPLIT distance="50" swimtime="00:00:28.29" />
                    <SPLIT distance="75" swimtime="00:00:44.97" />
                    <SPLIT distance="100" swimtime="00:01:02.34" />
                    <SPLIT distance="125" swimtime="00:01:19.98" />
                    <SPLIT distance="150" swimtime="00:01:38.21" />
                    <SPLIT distance="175" swimtime="00:01:56.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="567" reactiontime="+74" swimtime="00:01:01.77" resultid="3872" lane="4" heatid="6744" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.21" />
                    <SPLIT distance="50" swimtime="00:00:28.62" />
                    <SPLIT distance="75" swimtime="00:00:46.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="3875" lane="5" heatid="7066" entrytime="00:01:59.00" />
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="3876" lane="2" heatid="7293" entrytime="00:00:27.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1341" points="444" reactiontime="+74" swimtime="00:02:05.14" resultid="3878" lane="6" heatid="6988" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.15" />
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                    <SPLIT distance="75" swimtime="00:00:46.62" />
                    <SPLIT distance="100" swimtime="00:01:06.16" />
                    <SPLIT distance="125" swimtime="00:01:20.75" />
                    <SPLIT distance="150" swimtime="00:01:39.47" />
                    <SPLIT distance="175" swimtime="00:01:51.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3871" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="3848" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="3858" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="3856" number="4" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1177" points="558" reactiontime="+86" swimtime="00:01:45.40" resultid="3877" lane="5" heatid="6810" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.91" />
                    <SPLIT distance="50" swimtime="00:00:26.29" />
                    <SPLIT distance="75" swimtime="00:00:39.28" />
                    <SPLIT distance="100" swimtime="00:00:53.29" />
                    <SPLIT distance="125" swimtime="00:01:05.50" />
                    <SPLIT distance="150" swimtime="00:01:19.02" />
                    <SPLIT distance="175" swimtime="00:01:30.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3856" number="1" reactiontime="+86" />
                    <RELAYPOSITION athleteid="3866" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="3845" number="3" reactiontime="+17" />
                    <RELAYPOSITION athleteid="3871" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="OCOST" name="Oceanik Ostrzeszów" nation="POL">
          <CONTACT name="Burghardt" />
          <ATHLETES>
            <ATHLETE birthdate="1986-01-01" firstname="Nina" gender="F" lastname="Burghardt" nation="POL" athleteid="3887">
              <RESULTS>
                <RESULT eventid="1479" points="593" reactiontime="+68" swimtime="00:00:32.93" resultid="3889" lane="4" heatid="7031" entrytime="00:00:33.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="547" reactiontime="+72" swimtime="00:00:37.06" resultid="3888" lane="3" heatid="6853" entrytime="00:00:37.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="478" reactiontime="+75" swimtime="00:00:32.56" resultid="3890" lane="7" heatid="7280" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="521" reactiontime="+72" swimtime="00:00:29.78" resultid="3891" lane="6" heatid="7335" entrytime="00:00:29.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="POZNA" name="Poznań" nation="POL">
          <CONTACT name="g" />
          <ATHLETES>
            <ATHLETE birthdate="1968-09-07" firstname="Radosław" gender="M" lastname="Kwiek" nation="POL" athleteid="2698">
              <RESULTS>
                <RESULT eventid="1143" points="245" swimtime="00:23:15.97" resultid="2699" lane="1" heatid="6751" entrytime="00:22:30.00" entrycourse="SCM" />
                <RESULT eventid="1375" points="281" reactiontime="+100" swimtime="00:05:35.74" resultid="2701" lane="2" heatid="6906" entrytime="00:05:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.64" />
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                    <SPLIT distance="75" swimtime="00:00:53.45" />
                    <SPLIT distance="100" swimtime="00:01:12.56" />
                    <SPLIT distance="125" swimtime="00:01:32.79" />
                    <SPLIT distance="150" swimtime="00:01:54.23" />
                    <SPLIT distance="175" swimtime="00:02:15.78" />
                    <SPLIT distance="200" swimtime="00:02:37.38" />
                    <SPLIT distance="225" swimtime="00:02:59.19" />
                    <SPLIT distance="250" swimtime="00:03:21.32" />
                    <SPLIT distance="275" swimtime="00:03:43.50" />
                    <SPLIT distance="300" swimtime="00:04:05.87" />
                    <SPLIT distance="325" swimtime="00:04:28.66" />
                    <SPLIT distance="350" swimtime="00:04:51.28" />
                    <SPLIT distance="375" swimtime="00:05:13.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="306" reactiontime="+90" swimtime="00:02:32.73" resultid="2702" heatid="7061" entrytime="00:02:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.86" />
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                    <SPLIT distance="75" swimtime="00:00:51.99" />
                    <SPLIT distance="100" swimtime="00:01:11.39" />
                    <SPLIT distance="125" swimtime="00:01:31.15" />
                    <SPLIT distance="150" swimtime="00:01:51.77" />
                    <SPLIT distance="175" swimtime="00:02:13.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="327" reactiontime="+101" swimtime="00:01:08.23" resultid="2700" lane="2" heatid="6834" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.09" />
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                    <SPLIT distance="75" swimtime="00:00:49.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="2703" lane="6" heatid="7344" entrytime="00:00:30.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1974-01-01" firstname="Marcin" gender="M" lastname="Odziemski" nation="POL" athleteid="3900">
              <RESULTS>
                <RESULT eventid="1205" points="452" reactiontime="+81" swimtime="00:01:01.27" resultid="3901" lane="7" heatid="6844" entrytime="00:00:59.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.44" />
                    <SPLIT distance="50" swimtime="00:00:28.07" />
                    <SPLIT distance="75" swimtime="00:00:43.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="428" reactiontime="+81" swimtime="00:02:16.55" resultid="3903" lane="2" heatid="7064" entrytime="00:02:15.35">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.68" />
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                    <SPLIT distance="75" swimtime="00:00:47.50" />
                    <SPLIT distance="100" swimtime="00:01:04.23" />
                    <SPLIT distance="125" swimtime="00:01:21.42" />
                    <SPLIT distance="150" swimtime="00:01:39.48" />
                    <SPLIT distance="175" swimtime="00:01:57.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" status="DNS" swimtime="00:00:00.00" resultid="3902" heatid="6909" entrytime="00:04:45.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-01" firstname="Mateusz" gender="M" lastname="Powąska" nation="POL" athleteid="3904">
              <RESULTS>
                <RESULT eventid="1645" points="379" reactiontime="+69" swimtime="00:00:31.72" resultid="3906" lane="7" heatid="7291" entrytime="00:00:29.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="419" reactiontime="+70" swimtime="00:01:02.83" resultid="3905" lane="2" heatid="6844" entrytime="00:00:59.35">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.03" />
                    <SPLIT distance="50" swimtime="00:00:29.73" />
                    <SPLIT distance="75" swimtime="00:00:46.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="3907" lane="5" heatid="7349" entrytime="00:00:27.51" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Magdalena" gender="F" lastname="Tomczyk" nation="POL" athleteid="4081">
              <RESULTS>
                <RESULT eventid="1409" status="DNS" swimtime="00:00:00.00" resultid="4082" lane="6" heatid="6997" />
                <RESULT eventid="1679" status="DNS" swimtime="00:00:00.00" resultid="4083" lane="5" heatid="7295" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-01" firstname="Zygmunt" gender="M" lastname="Pawlaczek" nation="POL" athleteid="4502">
              <RESULTS>
                <RESULT eventid="1764" points="224" reactiontime="+107" swimtime="00:00:34.99" resultid="6213" heatid="7336" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="148" reactiontime="+116" swimtime="00:06:55.39" resultid="4505" lane="4" heatid="6899" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.95" />
                    <SPLIT distance="50" swimtime="00:00:41.54" />
                    <SPLIT distance="75" swimtime="00:01:05.57" />
                    <SPLIT distance="100" swimtime="00:01:30.46" />
                    <SPLIT distance="125" swimtime="00:01:55.92" />
                    <SPLIT distance="150" swimtime="00:02:23.20" />
                    <SPLIT distance="175" swimtime="00:02:50.00" />
                    <SPLIT distance="200" swimtime="00:03:17.44" />
                    <SPLIT distance="225" swimtime="00:03:44.33" />
                    <SPLIT distance="250" swimtime="00:04:11.60" />
                    <SPLIT distance="275" swimtime="00:04:39.00" />
                    <SPLIT distance="300" swimtime="00:05:06.90" />
                    <SPLIT distance="325" swimtime="00:05:34.44" />
                    <SPLIT distance="350" swimtime="00:06:02.16" />
                    <SPLIT distance="375" swimtime="00:06:30.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="186" reactiontime="+103" swimtime="00:01:22.28" resultid="4504" lane="3" heatid="6832" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.10" />
                    <SPLIT distance="50" swimtime="00:00:37.14" />
                    <SPLIT distance="75" swimtime="00:00:59.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="149" reactiontime="+117" swimtime="00:01:36.37" resultid="4503" lane="8" heatid="6732" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.86" />
                    <SPLIT distance="50" swimtime="00:00:46.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="162" reactiontime="+93" swimtime="00:00:44.88" resultid="6211" lane="1" heatid="7036" entrytime="00:00:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" status="DNS" swimtime="00:00:00.00" resultid="6212" lane="3" heatid="7304" entrytime="00:01:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1941-01-01" firstname="Zbigniew" gender="M" lastname="Radecki" nation="POL" athleteid="4506">
              <RESULTS>
                <RESULT eventid="1696" points="137" reactiontime="+79" swimtime="00:01:54.02" resultid="4509" lane="8" heatid="7303" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.07" />
                    <SPLIT distance="50" swimtime="00:00:53.11" />
                    <SPLIT distance="75" swimtime="00:01:22.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="132" reactiontime="+91" swimtime="00:04:10.25" resultid="4508" lane="7" heatid="7003" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.70" />
                    <SPLIT distance="50" swimtime="00:00:55.79" />
                    <SPLIT distance="75" swimtime="00:01:26.80" />
                    <SPLIT distance="100" swimtime="00:01:59.05" />
                    <SPLIT distance="125" swimtime="00:02:32.21" />
                    <SPLIT distance="150" swimtime="00:03:05.62" />
                    <SPLIT distance="175" swimtime="00:03:38.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="165" reactiontime="+90" swimtime="00:00:49.50" resultid="4507" lane="2" heatid="6854" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-01" firstname="Barbara" gender="F" lastname="Prange" nation="POL" athleteid="4510">
              <RESULTS>
                <RESULT comment="K 8 K 14" eventid="1222" reactiontime="+134" status="DSQ" swimtime="00:01:04.13" resultid="4511" lane="5" heatid="6847">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="RACIB" name="Racibórz" nation="POL">
          <CONTACT name="Piechula" />
          <ATHLETES>
            <ATHLETE birthdate="1957-01-01" firstname="Adolf" gender="M" lastname="Piechula" nation="POL" athleteid="3909">
              <RESULTS>
                <RESULT eventid="1273" points="235" reactiontime="+89" swimtime="00:03:01.48" resultid="3912" lane="3" heatid="6872" entrytime="00:03:05.67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.95" />
                    <SPLIT distance="50" swimtime="00:00:38.72" />
                    <SPLIT distance="75" swimtime="00:01:01.84" />
                    <SPLIT distance="100" swimtime="00:01:26.23" />
                    <SPLIT distance="125" swimtime="00:01:50.17" />
                    <SPLIT distance="150" swimtime="00:02:14.16" />
                    <SPLIT distance="175" swimtime="00:02:38.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="243" reactiontime="+83" swimtime="00:01:20.66" resultid="3913" lane="8" heatid="7019" entrytime="00:01:22.56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.74" />
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                    <SPLIT distance="75" swimtime="00:00:56.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="281" reactiontime="+83" swimtime="00:02:54.39" resultid="3914" lane="6" heatid="7076" entrytime="00:03:03.45">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.70" />
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                    <SPLIT distance="75" swimtime="00:00:59.87" />
                    <SPLIT distance="100" swimtime="00:01:21.90" />
                    <SPLIT distance="125" swimtime="00:01:48.26" />
                    <SPLIT distance="150" swimtime="00:02:14.22" />
                    <SPLIT distance="175" swimtime="00:02:35.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="312" reactiontime="+73" swimtime="00:01:26.83" resultid="3915" lane="7" heatid="7308" entrytime="00:01:25.67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.17" />
                    <SPLIT distance="50" swimtime="00:00:39.69" />
                    <SPLIT distance="75" swimtime="00:01:03.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="248" reactiontime="+93" swimtime="00:06:27.66" resultid="3916" lane="3" heatid="7361" entrytime="00:06:31.65">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.03" />
                    <SPLIT distance="50" swimtime="00:00:41.58" />
                    <SPLIT distance="75" swimtime="00:01:06.04" />
                    <SPLIT distance="100" swimtime="00:01:31.63" />
                    <SPLIT distance="125" swimtime="00:01:55.94" />
                    <SPLIT distance="150" swimtime="00:02:20.54" />
                    <SPLIT distance="175" swimtime="00:02:45.84" />
                    <SPLIT distance="200" swimtime="00:03:10.17" />
                    <SPLIT distance="225" swimtime="00:03:37.13" />
                    <SPLIT distance="250" swimtime="00:04:04.59" />
                    <SPLIT distance="275" swimtime="00:04:31.77" />
                    <SPLIT distance="300" swimtime="00:04:59.71" />
                    <SPLIT distance="325" swimtime="00:05:22.37" />
                    <SPLIT distance="350" swimtime="00:05:44.81" />
                    <SPLIT distance="375" swimtime="00:06:07.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="372" reactiontime="+78" swimtime="00:00:37.77" resultid="3911" lane="6" heatid="6861" entrytime="00:00:37.68">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="277" reactiontime="+75" swimtime="00:01:18.44" resultid="3910" lane="6" heatid="6738" entrytime="00:01:17.45">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.67" />
                    <SPLIT distance="50" swimtime="00:00:35.67" />
                    <SPLIT distance="75" swimtime="00:00:59.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="UMPOZ" name="UMKSN Poznań" nation="POL">
          <CONTACT name="Jakubowski" />
          <ATHLETES>
            <ATHLETE birthdate="1993-01-01" firstname="Sandra" gender="F" lastname="Michałowska" nation="POL" athleteid="3918">
              <RESULTS>
                <RESULT eventid="1713" points="379" reactiontime="+67" status="EXH" swimtime="00:01:21.14" resultid="4992" lane="3" heatid="7316" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.55" />
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                    <SPLIT distance="75" swimtime="00:00:59.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="428" reactiontime="+72" status="EXH" swimtime="00:00:36.70" resultid="4991" lane="3" heatid="7030" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="321" reactiontime="+81" status="EXH" swimtime="00:01:25.81" resultid="4990" lane="4" heatid="6728" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.85" />
                    <SPLIT distance="50" swimtime="00:00:38.55" />
                    <SPLIT distance="75" swimtime="00:01:06.67" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="04" eventid="1187" reactiontime="+62" status="DSQ" swimtime="00:01:10.69" resultid="4989" lane="5" heatid="6827" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.32" />
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                    <SPLIT distance="75" swimtime="00:00:51.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="466" reactiontime="+95" status="EXH" swimtime="00:00:30.91" resultid="6705" lane="3" heatid="7334" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="487" reactiontime="+83" swimtime="00:00:30.45" resultid="3919" lane="4" heatid="7044" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Bartosz" gender="M" lastname="Wróbel" nation="POL" athleteid="3920">
              <RESULTS>
                <RESULT eventid="1239" points="491" reactiontime="+75" status="EXH" swimtime="00:00:34.44" resultid="4994" lane="3" heatid="6864" entrytime="00:00:34.87">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="445" reactiontime="+73" status="EXH" swimtime="00:01:17.15" resultid="4995" lane="7" heatid="7310" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.77" />
                    <SPLIT distance="50" swimtime="00:00:36.70" />
                    <SPLIT distance="75" swimtime="00:00:57.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="324" reactiontime="+75" status="EXH" swimtime="00:00:35.62" resultid="4996" lane="7" heatid="7039" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="333" reactiontime="+93" status="EXH" swimtime="00:01:13.79" resultid="4993" lane="8" heatid="6740" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.79" />
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                    <SPLIT distance="75" swimtime="00:00:56.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="416" reactiontime="+71" status="EXH" swimtime="00:00:28.49" resultid="6706" lane="3" heatid="7345" entrytime="00:00:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1530" points="432" reactiontime="+73" swimtime="00:00:28.14" resultid="3921" lane="4" heatid="7047" entrytime="00:00:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Jan" gender="M" lastname="Kaptur" nation="POL" athleteid="3922">
              <RESULTS>
                <RESULT comment="Z 2" eventid="1109" reactiontime="+117" status="DSQ" swimtime="00:00:00.00" resultid="4997" lane="6" heatid="6730">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.38" />
                    <SPLIT distance="50" swimtime="00:00:46.61" />
                    <SPLIT distance="75" swimtime="00:01:17.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="178" reactiontime="+80" status="EXH" swimtime="00:01:23.63" resultid="4998" lane="1" heatid="6832" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.09" />
                    <SPLIT distance="50" swimtime="00:00:38.74" />
                    <SPLIT distance="75" swimtime="00:01:01.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="136" reactiontime="+72" status="EXH" swimtime="00:01:41.99" resultid="4999" heatid="7320" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.15" />
                    <SPLIT distance="50" swimtime="00:00:47.43" />
                    <SPLIT distance="75" swimtime="00:01:15.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="136" status="EXH" swimtime="00:00:47.57" resultid="5000" heatid="7032">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1530" points="184" reactiontime="+92" swimtime="00:00:37.38" resultid="3923" lane="4" heatid="7045">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Kacper" gender="M" lastname="Nowicki" nation="POL" athleteid="3924">
              <RESULTS>
                <RESULT eventid="1205" points="182" reactiontime="+98" status="EXH" swimtime="00:01:22.88" resultid="5001" lane="3" heatid="6831" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.54" />
                    <SPLIT distance="50" swimtime="00:00:39.44" />
                    <SPLIT distance="75" swimtime="00:01:01.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="164" reactiontime="+88" status="EXH" swimtime="00:00:44.62" resultid="5002" lane="1" heatid="7032">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="138" reactiontime="+89" status="EXH" swimtime="00:00:44.43" resultid="5003" lane="4" heatid="7281" entrytime="00:00:48.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.84" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="04" eventid="1109" reactiontime="+67" status="DSQ" swimtime="00:00:00.00" resultid="6232" lane="5" heatid="6730">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.21" />
                    <SPLIT distance="50" swimtime="00:00:44.42" />
                    <SPLIT distance="75" swimtime="00:01:14.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1530" points="186" reactiontime="+101" swimtime="00:00:37.26" resultid="3925" lane="2" heatid="7046">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Weronika" gender="F" lastname="Nowicka" nation="POL" athleteid="3926">
              <RESULTS>
                <RESULT eventid="1641" points="131" status="EXH" swimtime="00:00:50.12" resultid="5006" lane="8" heatid="7277" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="173" reactiontime="+67" status="EXH" swimtime="00:00:49.63" resultid="5005" lane="4" heatid="7024">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="196" reactiontime="+67" status="EXH" swimtime="00:01:30.90" resultid="5004" lane="6" heatid="6823" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.15" />
                    <SPLIT distance="50" swimtime="00:00:41.77" />
                    <SPLIT distance="75" swimtime="00:01:07.32" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="04" eventid="1092" status="DSQ" swimtime="00:00:00.00" resultid="6233" lane="6" heatid="6723">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.94" />
                    <SPLIT distance="50" swimtime="00:00:52.73" />
                    <SPLIT distance="75" swimtime="00:01:23.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="207" reactiontime="+79" swimtime="00:00:40.52" resultid="3927" lane="7" heatid="7044">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Wanessa" gender="F" lastname="Stoinska" nation="POL" athleteid="3928">
              <RESULTS>
                <RESULT eventid="1187" points="207" reactiontime="+125" status="EXH" swimtime="00:01:29.28" resultid="5007" lane="1" heatid="6823" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.98" />
                    <SPLIT distance="50" swimtime="00:00:42.40" />
                    <SPLIT distance="75" swimtime="00:01:06.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="175" reactiontime="+82" status="EXH" swimtime="00:00:49.41" resultid="5008" lane="7" heatid="7025">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="114" reactiontime="+117" status="EXH" swimtime="00:00:52.39" resultid="5009" lane="5" heatid="7276" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="210" reactiontime="+114" swimtime="00:00:40.28" resultid="3929" lane="2" heatid="7044">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Sara" gender="F" lastname="Plewczyńska" nation="POL" athleteid="3930">
              <RESULTS>
                <RESULT eventid="1479" points="134" reactiontime="+79" status="EXH" swimtime="00:00:54.03" resultid="5010" lane="1" heatid="7025">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="107" swimtime="00:00:50.42" resultid="3931" lane="5" heatid="7044">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WIOST" name="Wieloboista Ostrów Wlkp" nation="POL">
          <CONTACT name="k" />
          <ATHLETES>
            <ATHLETE birthdate="1965-01-01" firstname="Bogusław" gender="M" lastname="Wawrzyniak" nation="POL" athleteid="3933">
              <RESULTS>
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="3940" lane="8" heatid="7342" entrytime="00:00:32.00" />
                <RESULT eventid="1462" status="DNS" swimtime="00:00:00.00" resultid="3937" lane="8" heatid="7017" entrytime="00:01:35.00" />
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="3939" lane="2" heatid="7284" entrytime="00:00:37.00" />
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="3938" lane="3" heatid="7058" entrytime="00:02:45.00" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="3936" lane="7" heatid="6871" entrytime="00:03:30.00" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="3935" lane="1" heatid="6836" entrytime="00:01:11.00" />
                <RESULT eventid="1143" status="DNS" swimtime="00:00:00.00" resultid="3934" lane="6" heatid="6750" entrytime="00:24:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-01-01" firstname="Krzysztof" gender="M" lastname="Kaźmierowski" nation="POL" athleteid="4888">
              <RESULTS>
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="4894" heatid="7339" entrytime="00:00:35.00" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="4889" lane="8" heatid="6855" entrytime="00:00:55.00" />
                <RESULT eventid="1307" status="DNS" swimtime="00:00:00.00" resultid="4890" lane="2" heatid="6881" entrytime="00:04:30.00" />
                <RESULT eventid="1496" status="DNS" swimtime="00:00:00.00" resultid="4891" lane="5" heatid="7033" entrytime="00:00:55.00" />
                <RESULT eventid="1730" status="DNS" swimtime="00:00:00.00" resultid="4893" lane="4" heatid="7318" entrytime="00:02:10.00" />
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="4892" lane="4" heatid="7054" entrytime="00:03:50.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="FLGDY" name="WKS Flota Gdynia" nation="POL">
          <CONTACT name="Kuźniak" />
          <ATHLETES>
            <ATHLETE birthdate="1931-01-01" firstname="Zbigniew" gender="M" lastname="Zajączkowski" nation="POL" athleteid="3942">
              <RESULTS>
                <RESULT comment="Rekord Polski " eventid="1205" points="47" reactiontime="+111" swimtime="00:02:10.34" resultid="3943" lane="8" heatid="6831" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.16" />
                    <SPLIT distance="75" swimtime="00:01:36.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="61" reactiontime="+93" swimtime="00:00:54.04" resultid="3944" lane="5" heatid="7336" entrytime="00:00:49.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1934-01-01" firstname="Bogdan" gender="M" lastname="Ciundziewicki" nation="POL" athleteid="3945">
              <RESULTS>
                <RESULT eventid="1696" points="168" swimtime="00:01:46.58" resultid="3948" lane="5" heatid="7304" entrytime="00:01:41.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.20" />
                    <SPLIT distance="50" swimtime="00:00:49.78" />
                    <SPLIT distance="75" swimtime="00:01:18.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="205" reactiontime="+90" swimtime="00:00:46.04" resultid="3946" lane="4" heatid="6856" entrytime="00:00:44.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" status="DNS" swimtime="00:00:00.00" resultid="3947" heatid="7005" entrytime="00:03:41.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Czesław" gender="M" lastname="Mikołajczyk" nation="POL" athleteid="3949">
              <RESULTS>
                <RESULT eventid="1696" points="225" reactiontime="+98" swimtime="00:01:36.79" resultid="3953" lane="3" heatid="7305" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.53" />
                    <SPLIT distance="50" swimtime="00:00:46.47" />
                    <SPLIT distance="75" swimtime="00:01:11.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="257" reactiontime="+101" swimtime="00:00:42.72" resultid="3951" heatid="6858" entrytime="00:00:42.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="150" reactiontime="+99" swimtime="00:07:38.08" resultid="3954" lane="2" heatid="7359" entrytime="00:07:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.43" />
                    <SPLIT distance="50" swimtime="00:00:51.71" />
                    <SPLIT distance="75" swimtime="00:01:21.63" />
                    <SPLIT distance="100" swimtime="00:01:52.54" />
                    <SPLIT distance="125" swimtime="00:02:23.65" />
                    <SPLIT distance="150" swimtime="00:02:53.47" />
                    <SPLIT distance="175" swimtime="00:03:26.99" />
                    <SPLIT distance="200" swimtime="00:03:57.74" />
                    <SPLIT distance="225" swimtime="00:04:29.10" />
                    <SPLIT distance="250" swimtime="00:04:59.61" />
                    <SPLIT distance="275" swimtime="00:05:28.71" />
                    <SPLIT distance="300" swimtime="00:05:58.42" />
                    <SPLIT distance="350" swimtime="00:07:38.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="206" reactiontime="+110" swimtime="00:03:35.72" resultid="3952" lane="2" heatid="7005" entrytime="00:03:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.21" />
                    <SPLIT distance="50" swimtime="00:00:48.94" />
                    <SPLIT distance="75" swimtime="00:01:16.23" />
                    <SPLIT distance="100" swimtime="00:01:43.88" />
                    <SPLIT distance="125" swimtime="00:02:11.43" />
                    <SPLIT distance="150" swimtime="00:02:39.50" />
                    <SPLIT distance="175" swimtime="00:03:08.00" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Z 2" eventid="1109" reactiontime="+104" status="DSQ" swimtime="00:01:32.61" resultid="3950" heatid="6734" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.23" />
                    <SPLIT distance="50" swimtime="00:00:47.21" />
                    <SPLIT distance="75" swimtime="00:01:10.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Witosława" gender="F" lastname="Olechnicka" nation="POL" athleteid="3955">
              <RESULTS>
                <RESULT eventid="1445" points="143" reactiontime="+97" swimtime="00:01:48.23" resultid="3957" heatid="7013" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.34" />
                    <SPLIT distance="50" swimtime="00:00:51.63" />
                    <SPLIT distance="75" swimtime="00:01:20.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="187" reactiontime="+97" swimtime="00:00:44.51" resultid="3958" lane="4" heatid="7276" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="239" reactiontime="+86" swimtime="00:01:25.11" resultid="3956" lane="5" heatid="6824" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.52" />
                    <SPLIT distance="50" swimtime="00:00:39.77" />
                    <SPLIT distance="75" swimtime="00:01:02.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="198" reactiontime="+72" swimtime="00:01:40.82" resultid="3959" lane="8" heatid="7315" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.01" />
                    <SPLIT distance="50" swimtime="00:00:48.31" />
                    <SPLIT distance="75" swimtime="00:01:14.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Jola" gender="F" lastname="Dołżyńska" nation="POL" athleteid="3960">
              <RESULTS>
                <RESULT eventid="1409" points="153" reactiontime="+102" swimtime="00:04:22.13" resultid="3962" lane="2" heatid="6998" entrytime="00:04:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.49" />
                    <SPLIT distance="50" swimtime="00:01:00.83" />
                    <SPLIT distance="75" swimtime="00:01:34.56" />
                    <SPLIT distance="100" swimtime="00:02:08.85" />
                    <SPLIT distance="125" swimtime="00:02:43.01" />
                    <SPLIT distance="150" swimtime="00:03:16.93" />
                    <SPLIT distance="175" swimtime="00:03:50.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="132" reactiontime="+91" swimtime="00:04:05.77" resultid="3961" lane="8" heatid="6877" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.28" />
                    <SPLIT distance="50" swimtime="00:00:56.81" />
                    <SPLIT distance="75" swimtime="00:01:26.92" />
                    <SPLIT distance="100" swimtime="00:01:58.24" />
                    <SPLIT distance="125" swimtime="00:02:30.49" />
                    <SPLIT distance="150" swimtime="00:03:02.47" />
                    <SPLIT distance="175" swimtime="00:03:35.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-01-01" firstname="Ewa" gender="F" lastname="Mierwald" nation="POL" athleteid="3963">
              <RESULTS>
                <RESULT eventid="1222" points="227" reactiontime="+106" swimtime="00:00:49.67" resultid="3965" lane="2" heatid="6850" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="204" reactiontime="+115" swimtime="00:01:50.54" resultid="3968" lane="7" heatid="7298" entrytime="00:01:47.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.74" />
                    <SPLIT distance="50" swimtime="00:00:52.90" />
                    <SPLIT distance="75" swimtime="00:01:21.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1581" points="176" reactiontime="+109" swimtime="00:03:49.16" resultid="3967" lane="1" heatid="7068" entrytime="00:03:54.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.77" />
                    <SPLIT distance="50" swimtime="00:00:52.67" />
                    <SPLIT distance="75" swimtime="00:01:22.13" />
                    <SPLIT distance="100" swimtime="00:01:52.00" />
                    <SPLIT distance="125" swimtime="00:02:22.54" />
                    <SPLIT distance="150" swimtime="00:02:53.20" />
                    <SPLIT distance="175" swimtime="00:03:20.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="194" reactiontime="+86" swimtime="00:00:47.77" resultid="3966" lane="2" heatid="7027" entrytime="00:00:47.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="183" reactiontime="+115" swimtime="00:01:43.50" resultid="3964" lane="8" heatid="6725" entrytime="00:01:48.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.50" />
                    <SPLIT distance="50" swimtime="00:00:49.05" />
                    <SPLIT distance="75" swimtime="00:01:17.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-01" firstname="Karina" gender="F" lastname="Marszałek" nation="POL" athleteid="3969">
              <RESULTS>
                <RESULT eventid="1256" points="122" reactiontime="+133" swimtime="00:04:09.87" resultid="3972" lane="7" heatid="6868" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.70" />
                    <SPLIT distance="50" swimtime="00:00:53.79" />
                    <SPLIT distance="75" swimtime="00:01:24.33" />
                    <SPLIT distance="100" swimtime="00:01:55.65" />
                    <SPLIT distance="125" swimtime="00:02:31.16" />
                    <SPLIT distance="150" swimtime="00:03:04.14" />
                    <SPLIT distance="175" swimtime="00:03:38.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1581" points="192" reactiontime="+105" swimtime="00:03:42.52" resultid="3974" lane="5" heatid="7068" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.81" />
                    <SPLIT distance="50" swimtime="00:00:54.09" />
                    <SPLIT distance="75" swimtime="00:02:21.95" />
                    <SPLIT distance="100" swimtime="00:01:53.63" />
                    <SPLIT distance="125" swimtime="00:03:18.28" />
                    <SPLIT distance="150" swimtime="00:02:50.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1445" points="129" reactiontime="+99" swimtime="00:01:51.85" resultid="3973" lane="2" heatid="7013" entrytime="00:01:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.16" />
                    <SPLIT distance="50" swimtime="00:00:53.25" />
                    <SPLIT distance="75" swimtime="00:01:23.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1781" points="196" reactiontime="+120" swimtime="00:07:43.11" resultid="3975" heatid="7356" entrytime="00:07:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.44" />
                    <SPLIT distance="50" swimtime="00:00:54.13" />
                    <SPLIT distance="75" swimtime="00:01:23.35" />
                    <SPLIT distance="100" swimtime="00:01:56.39" />
                    <SPLIT distance="125" swimtime="00:02:28.14" />
                    <SPLIT distance="150" swimtime="00:02:57.56" />
                    <SPLIT distance="175" swimtime="00:03:27.23" />
                    <SPLIT distance="200" swimtime="00:03:56.55" />
                    <SPLIT distance="225" swimtime="00:04:26.90" />
                    <SPLIT distance="250" swimtime="00:04:57.38" />
                    <SPLIT distance="275" swimtime="00:05:26.28" />
                    <SPLIT distance="300" swimtime="00:05:57.30" />
                    <SPLIT distance="325" swimtime="00:06:24.84" />
                    <SPLIT distance="350" swimtime="00:06:52.35" />
                    <SPLIT distance="375" swimtime="00:07:19.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="203" reactiontime="+107" swimtime="00:01:40.01" resultid="3970" lane="4" heatid="6725" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.11" />
                    <SPLIT distance="50" swimtime="00:00:48.13" />
                    <SPLIT distance="75" swimtime="00:01:15.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="250" reactiontime="+107" swimtime="00:00:48.07" resultid="3971" lane="8" heatid="6851" entrytime="00:00:48.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WOTCZ" name="WOPR Tczew" nation="POL">
          <CONTACT name="o" />
          <ATHLETES>
            <ATHLETE birthdate="1987-01-01" firstname="Aleksandra" gender="F" lastname="Hebel" nation="POL" athleteid="3977">
              <RESULTS>
                <RESULT eventid="1747" points="344" reactiontime="+94" swimtime="00:00:34.19" resultid="3981" lane="4" heatid="7333" entrytime="00:00:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="324" reactiontime="+91" swimtime="00:01:16.99" resultid="3978" lane="6" heatid="6826" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.36" />
                    <SPLIT distance="50" swimtime="00:00:36.97" />
                    <SPLIT distance="75" swimtime="00:00:57.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="266" reactiontime="+109" swimtime="00:02:58.49" resultid="3980" lane="1" heatid="7051" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.03" />
                    <SPLIT distance="50" swimtime="00:00:38.85" />
                    <SPLIT distance="75" swimtime="00:01:00.60" />
                    <SPLIT distance="100" swimtime="00:01:23.19" />
                    <SPLIT distance="125" swimtime="00:01:46.45" />
                    <SPLIT distance="150" swimtime="00:02:10.95" />
                    <SPLIT distance="175" swimtime="00:02:35.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="274" reactiontime="+66" swimtime="00:00:42.60" resultid="3979" lane="7" heatid="7029" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Kamila" gender="F" lastname="Ormianin" nation="POL" athleteid="4628">
              <RESULTS>
                <RESULT eventid="1058" points="455" swimtime="00:10:42.25" resultid="4629" lane="3" heatid="6715" entrytime="00:11:00.00" />
                <RESULT eventid="1547" points="518" reactiontime="+74" swimtime="00:02:22.93" resultid="4632" lane="4" heatid="7053" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.47" />
                    <SPLIT distance="50" swimtime="00:00:32.84" />
                    <SPLIT distance="75" swimtime="00:00:50.59" />
                    <SPLIT distance="100" swimtime="00:01:08.75" />
                    <SPLIT distance="125" swimtime="00:01:27.51" />
                    <SPLIT distance="150" swimtime="00:01:46.59" />
                    <SPLIT distance="175" swimtime="00:02:05.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="484" reactiontime="+80" swimtime="00:05:07.47" resultid="4631" lane="7" heatid="6898" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.16" />
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                    <SPLIT distance="75" swimtime="00:00:54.13" />
                    <SPLIT distance="100" swimtime="00:01:13.92" />
                    <SPLIT distance="125" swimtime="00:01:33.00" />
                    <SPLIT distance="150" swimtime="00:01:52.43" />
                    <SPLIT distance="175" swimtime="00:02:12.32" />
                    <SPLIT distance="200" swimtime="00:02:31.97" />
                    <SPLIT distance="225" swimtime="00:02:51.25" />
                    <SPLIT distance="250" swimtime="00:03:10.61" />
                    <SPLIT distance="275" swimtime="00:03:30.13" />
                    <SPLIT distance="300" swimtime="00:03:49.86" />
                    <SPLIT distance="325" swimtime="00:04:09.46" />
                    <SPLIT distance="350" swimtime="00:04:28.97" />
                    <SPLIT distance="375" swimtime="00:04:48.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="489" reactiontime="+71" swimtime="00:01:07.08" resultid="4630" lane="2" heatid="6828" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.05" />
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                    <SPLIT distance="75" swimtime="00:00:49.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="479" reactiontime="+72" swimtime="00:00:30.63" resultid="4633" lane="1" heatid="7335" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ALWAR" name="AZS Almamer Warszawa" nation="POL">
          <CONTACT name="Sołtyk" />
          <ATHLETES>
            <ATHLETE birthdate="1974-01-01" firstname="Judyta" gender="F" lastname="Sołtyk" nation="POL" athleteid="3983">
              <RESULTS>
                <RESULT eventid="1058" points="405" swimtime="00:11:07.48" resultid="3984" lane="4" heatid="6715" entrytime="00:10:50.00" />
                <RESULT eventid="1358" points="427" reactiontime="+84" swimtime="00:05:20.52" resultid="3985" lane="2" heatid="6898" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.09" />
                    <SPLIT distance="50" swimtime="00:00:36.09" />
                    <SPLIT distance="75" swimtime="00:00:55.43" />
                    <SPLIT distance="100" swimtime="00:01:15.27" />
                    <SPLIT distance="125" swimtime="00:01:35.00" />
                    <SPLIT distance="150" swimtime="00:01:55.03" />
                    <SPLIT distance="175" swimtime="00:02:15.10" />
                    <SPLIT distance="200" swimtime="00:02:35.37" />
                    <SPLIT distance="225" swimtime="00:02:55.79" />
                    <SPLIT distance="250" swimtime="00:03:16.72" />
                    <SPLIT distance="275" swimtime="00:03:37.32" />
                    <SPLIT distance="300" swimtime="00:03:58.28" />
                    <SPLIT distance="325" swimtime="00:04:19.21" />
                    <SPLIT distance="350" swimtime="00:04:40.19" />
                    <SPLIT distance="375" swimtime="00:05:00.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" status="DNS" swimtime="00:00:00.00" resultid="3986" heatid="7053" entrytime="00:02:32.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="BIALY" name="Białystok" nation="POL">
          <CONTACT name="Dziekoński" />
          <ATHLETES>
            <ATHLETE birthdate="1943-01-01" firstname="Edward" gender="M" lastname="Dziekoński" nation="POL" athleteid="3988">
              <RESULTS>
                <RESULT eventid="1462" status="DNS" swimtime="00:00:00.00" resultid="3992" lane="2" heatid="7016" entrytime="00:01:46.00" />
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="3994" lane="2" heatid="7282" entrytime="00:00:43.00" />
                <RESULT eventid="1496" status="DNS" swimtime="00:00:00.00" resultid="3993" lane="1" heatid="7035" entrytime="00:00:47.00" />
                <RESULT eventid="1375" status="DNS" swimtime="00:00:00.00" resultid="3991" lane="4" heatid="6900" entrytime="00:07:12.00" />
                <RESULT eventid="1307" status="DNS" swimtime="00:00:00.00" resultid="3990" lane="2" heatid="6882" entrytime="00:03:49.00" />
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="3989" lane="5" heatid="6717" entrytime="00:14:50.00" />
                <RESULT eventid="1730" status="DNS" swimtime="00:00:00.00" resultid="3995" lane="1" heatid="7320" entrytime="00:01:47.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DEINO" name="Delfin Inowrocław" nation="POL">
          <CONTACT name="Lewandowski" />
          <ATHLETES>
            <ATHLETE birthdate="1937-01-01" firstname="Zygmunt" gender="M" lastname="Lewandowski" nation="POL" athleteid="3997">
              <RESULTS>
                <RESULT eventid="1143" points="144" swimtime="00:27:46.72" resultid="3998" lane="8" heatid="6749" entrytime="00:31:00.00" />
                <RESULT eventid="1564" points="144" reactiontime="+106" swimtime="00:03:16.17" resultid="4000" lane="2" heatid="7055" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.24" />
                    <SPLIT distance="50" swimtime="00:00:43.41" />
                    <SPLIT distance="75" swimtime="00:01:07.42" />
                    <SPLIT distance="100" swimtime="00:01:32.85" />
                    <SPLIT distance="125" swimtime="00:01:58.47" />
                    <SPLIT distance="150" swimtime="00:02:25.03" />
                    <SPLIT distance="175" swimtime="00:02:51.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="146" reactiontime="+97" swimtime="00:06:57.14" resultid="3999" lane="2" heatid="6900" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.30" />
                    <SPLIT distance="50" swimtime="00:00:47.14" />
                    <SPLIT distance="75" swimtime="00:01:13.05" />
                    <SPLIT distance="100" swimtime="00:01:39.38" />
                    <SPLIT distance="125" swimtime="00:02:05.87" />
                    <SPLIT distance="150" swimtime="00:02:32.75" />
                    <SPLIT distance="175" swimtime="00:02:59.43" />
                    <SPLIT distance="200" swimtime="00:03:27.02" />
                    <SPLIT distance="225" swimtime="00:03:53.47" />
                    <SPLIT distance="250" swimtime="00:04:20.14" />
                    <SPLIT distance="275" swimtime="00:04:46.94" />
                    <SPLIT distance="300" swimtime="00:05:13.65" />
                    <SPLIT distance="325" swimtime="00:05:39.73" />
                    <SPLIT distance="350" swimtime="00:06:06.14" />
                    <SPLIT distance="375" swimtime="00:06:32.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="104" swimtime="00:00:48.71" resultid="4001" lane="3" heatid="7281" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="HEKAI" name="Helyopolis Kair" nation="POL" region="WIE">
          <CONTACT name="Makay" />
          <ATHLETES>
            <ATHLETE birthdate="1950-01-01" firstname="Marek" gender="M" lastname="Makay" nation="POL" athleteid="4003">
              <RESULTS>
                <RESULT comment="Rekord Polski " eventid="1075" points="290" swimtime="00:11:32.37" resultid="4004" lane="1" heatid="6719" entrytime="00:12:20.00" />
                <RESULT eventid="1375" points="278" swimtime="00:05:37.20" resultid="4006" lane="3" heatid="6904" entrytime="00:05:48.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.68" />
                    <SPLIT distance="50" swimtime="00:00:38.28" />
                    <SPLIT distance="75" swimtime="00:00:58.89" />
                    <SPLIT distance="100" swimtime="00:01:19.61" />
                    <SPLIT distance="125" swimtime="00:01:41.25" />
                    <SPLIT distance="150" swimtime="00:02:02.80" />
                    <SPLIT distance="175" swimtime="00:02:25.00" />
                    <SPLIT distance="200" swimtime="00:02:46.74" />
                    <SPLIT distance="225" swimtime="00:03:08.10" />
                    <SPLIT distance="250" swimtime="00:03:29.87" />
                    <SPLIT distance="275" swimtime="00:03:51.43" />
                    <SPLIT distance="300" swimtime="00:04:13.23" />
                    <SPLIT distance="325" swimtime="00:04:34.64" />
                    <SPLIT distance="350" swimtime="00:04:56.34" />
                    <SPLIT distance="375" swimtime="00:05:17.34" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1564" points="293" reactiontime="+110" swimtime="00:02:34.91" resultid="4008" lane="6" heatid="7058" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.24" />
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                    <SPLIT distance="75" swimtime="00:00:55.04" />
                    <SPLIT distance="100" swimtime="00:01:14.51" />
                    <SPLIT distance="125" swimtime="00:01:34.57" />
                    <SPLIT distance="150" swimtime="00:01:55.30" />
                    <SPLIT distance="175" swimtime="00:02:15.40" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1730" points="249" reactiontime="+66" swimtime="00:01:23.48" resultid="4009" lane="8" heatid="7322" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.03" />
                    <SPLIT distance="50" swimtime="00:00:40.83" />
                    <SPLIT distance="75" swimtime="00:01:02.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="303" reactiontime="+121" swimtime="00:01:10.02" resultid="4005" lane="8" heatid="6836" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.82" />
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                    <SPLIT distance="75" swimtime="00:00:51.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="240" reactiontime="+70" swimtime="00:00:39.33" resultid="4007" heatid="7037" entrytime="00:00:39.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="309" reactiontime="+95" swimtime="00:00:31.45" resultid="4010" lane="6" heatid="7341" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KIELC" name="Kielce" nation="POL">
          <CONTACT name="Zembala" />
          <ATHLETES>
            <ATHLETE birthdate="1971-01-01" firstname="Tomasz" gender="M" lastname="Zembala" nation="POL" athleteid="4012">
              <RESULTS>
                <RESULT eventid="1375" points="264" reactiontime="+107" swimtime="00:05:42.90" resultid="4015" lane="1" heatid="6904" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.36" />
                    <SPLIT distance="50" swimtime="00:00:38.72" />
                    <SPLIT distance="75" swimtime="00:00:59.36" />
                    <SPLIT distance="100" swimtime="00:01:20.20" />
                    <SPLIT distance="125" swimtime="00:01:41.72" />
                    <SPLIT distance="150" swimtime="00:02:03.48" />
                    <SPLIT distance="175" swimtime="00:02:25.26" />
                    <SPLIT distance="200" swimtime="00:02:47.22" />
                    <SPLIT distance="225" swimtime="00:03:08.53" />
                    <SPLIT distance="250" swimtime="00:03:30.37" />
                    <SPLIT distance="275" swimtime="00:03:52.75" />
                    <SPLIT distance="300" swimtime="00:04:15.61" />
                    <SPLIT distance="325" swimtime="00:04:37.76" />
                    <SPLIT distance="350" swimtime="00:05:00.32" />
                    <SPLIT distance="375" swimtime="00:05:21.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="243" swimtime="00:12:14.10" resultid="4013" lane="5" heatid="6720" entrytime="00:12:00.00" />
                <RESULT eventid="1462" points="151" reactiontime="+108" swimtime="00:01:34.63" resultid="4016" lane="1" heatid="7019" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.91" />
                    <SPLIT distance="50" swimtime="00:00:43.21" />
                    <SPLIT distance="75" swimtime="00:01:09.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="207" reactiontime="+105" swimtime="00:00:38.77" resultid="4018" lane="2" heatid="7285" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="299" reactiontime="+100" swimtime="00:00:31.80" resultid="4019" lane="8" heatid="7343" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" status="DNS" swimtime="00:00:00.00" resultid="4017" heatid="7074" entrytime="00:03:30.00" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="4014" lane="4" heatid="6870" entrytime="00:03:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KOLOB" name="Kołobrzeg" nation="POL">
          <CONTACT name="Rogiński" />
          <ATHLETES>
            <ATHLETE birthdate="1971-01-01" firstname="Mariusz" gender="M" lastname="Rogiński" nation="POL" athleteid="4021">
              <RESULTS>
                <RESULT eventid="1645" points="334" reactiontime="+79" swimtime="00:00:33.06" resultid="4023" lane="1" heatid="7289" entrytime="00:00:31.28">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="371" reactiontime="+76" swimtime="00:00:29.59" resultid="4024" lane="2" heatid="7346" entrytime="00:00:28.54">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="4022" lane="4" heatid="6839" entrytime="00:01:06.45" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Jacek" gender="M" lastname="Dziarek" nation="POL" athleteid="4025">
              <RESULTS>
                <RESULT eventid="1564" points="297" reactiontime="+108" swimtime="00:02:34.22" resultid="4029" lane="5" heatid="7060" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.61" />
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                    <SPLIT distance="75" swimtime="00:00:52.90" />
                    <SPLIT distance="100" swimtime="00:01:12.22" />
                    <SPLIT distance="125" swimtime="00:01:32.01" />
                    <SPLIT distance="150" swimtime="00:01:52.78" />
                    <SPLIT distance="175" swimtime="00:02:13.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="278" swimtime="00:22:18.78" resultid="4026" lane="6" heatid="6751" entrytime="00:22:30.00" />
                <RESULT eventid="1764" points="335" reactiontime="+109" swimtime="00:00:30.61" resultid="4031" lane="6" heatid="7343" entrytime="00:00:30.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="326" reactiontime="+112" swimtime="00:01:08.30" resultid="4027" lane="7" heatid="6838" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.66" />
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                    <SPLIT distance="75" swimtime="00:00:51.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="278" reactiontime="+110" swimtime="00:05:36.90" resultid="4028" lane="4" heatid="6905" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.87" />
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                    <SPLIT distance="75" swimtime="00:00:56.90" />
                    <SPLIT distance="100" swimtime="00:01:16.92" />
                    <SPLIT distance="125" swimtime="00:01:38.34" />
                    <SPLIT distance="150" swimtime="00:01:59.98" />
                    <SPLIT distance="175" swimtime="00:02:21.75" />
                    <SPLIT distance="200" swimtime="00:02:43.24" />
                    <SPLIT distance="225" swimtime="00:03:05.31" />
                    <SPLIT distance="250" swimtime="00:03:27.33" />
                    <SPLIT distance="275" swimtime="00:03:49.23" />
                    <SPLIT distance="300" swimtime="00:04:11.29" />
                    <SPLIT distance="325" swimtime="00:04:33.23" />
                    <SPLIT distance="350" swimtime="00:04:54.48" />
                    <SPLIT distance="375" swimtime="00:05:15.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="4030" lane="6" heatid="7284" entrytime="00:00:37.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Jakub" gender="M" lastname="Jankowski" nation="POL" athleteid="4032">
              <RESULTS>
                <RESULT eventid="1075" points="244" swimtime="00:12:13.75" resultid="4033" lane="4" heatid="6720" entrytime="00:11:58.40" />
                <RESULT eventid="1375" points="271" reactiontime="+129" swimtime="00:05:40.00" resultid="4035" lane="6" heatid="6906" entrytime="00:05:30.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.94" />
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                    <SPLIT distance="75" swimtime="00:00:54.68" />
                    <SPLIT distance="100" swimtime="00:01:14.77" />
                    <SPLIT distance="125" swimtime="00:01:35.89" />
                    <SPLIT distance="150" swimtime="00:01:57.30" />
                    <SPLIT distance="175" swimtime="00:02:19.14" />
                    <SPLIT distance="200" swimtime="00:02:40.84" />
                    <SPLIT distance="225" swimtime="00:03:03.12" />
                    <SPLIT distance="250" swimtime="00:03:25.46" />
                    <SPLIT distance="275" swimtime="00:03:48.14" />
                    <SPLIT distance="300" swimtime="00:04:10.47" />
                    <SPLIT distance="325" swimtime="00:04:33.37" />
                    <SPLIT distance="350" swimtime="00:04:56.38" />
                    <SPLIT distance="375" swimtime="00:05:19.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="311" reactiontime="+126" swimtime="00:02:31.94" resultid="4036" lane="4" heatid="7060" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.03" />
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                    <SPLIT distance="75" swimtime="00:00:51.08" />
                    <SPLIT distance="100" swimtime="00:01:10.11" />
                    <SPLIT distance="125" swimtime="00:01:29.86" />
                    <SPLIT distance="150" swimtime="00:01:50.36" />
                    <SPLIT distance="175" swimtime="00:02:11.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="365" reactiontime="+111" swimtime="00:01:05.78" resultid="4034" lane="8" heatid="6840" entrytime="00:01:06.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.79" />
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                    <SPLIT distance="75" swimtime="00:00:48.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="4037" lane="7" heatid="7345" entrytime="00:00:29.30" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KRIVB" name="Krivbassmasters" nation="UKR">
          <CONTACT name="Sklyar" />
          <ATHLETES>
            <ATHLETE birthdate="1968-01-01" firstname="Konstantin" gender="M" lastname="Sklyar" nation="UKR" athleteid="4039">
              <RESULTS>
                <RESULT eventid="1375" points="403" reactiontime="+89" swimtime="00:04:57.81" resultid="4041" lane="2" heatid="6907" entrytime="00:05:10.31">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.99" />
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                    <SPLIT distance="75" swimtime="00:00:51.94" />
                    <SPLIT distance="100" swimtime="00:01:10.08" />
                    <SPLIT distance="125" swimtime="00:01:28.74" />
                    <SPLIT distance="150" swimtime="00:01:47.71" />
                    <SPLIT distance="175" swimtime="00:02:06.39" />
                    <SPLIT distance="200" swimtime="00:02:25.55" />
                    <SPLIT distance="225" swimtime="00:02:44.61" />
                    <SPLIT distance="250" swimtime="00:03:03.83" />
                    <SPLIT distance="275" swimtime="00:03:23.00" />
                    <SPLIT distance="300" swimtime="00:03:42.55" />
                    <SPLIT distance="325" swimtime="00:04:01.67" />
                    <SPLIT distance="350" swimtime="00:04:21.20" />
                    <SPLIT distance="375" swimtime="00:04:39.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="380" swimtime="00:10:32.75" resultid="4040" lane="5" heatid="6721" entrytime="00:10:59.34" />
                <RESULT eventid="1798" points="324" reactiontime="+74" swimtime="00:05:54.93" resultid="4043" lane="6" heatid="7363" entrytime="00:06:07.67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.52" />
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                    <SPLIT distance="75" swimtime="00:00:58.85" />
                    <SPLIT distance="100" swimtime="00:01:20.51" />
                    <SPLIT distance="125" swimtime="00:01:45.23" />
                    <SPLIT distance="150" swimtime="00:02:09.20" />
                    <SPLIT distance="175" swimtime="00:02:32.41" />
                    <SPLIT distance="200" swimtime="00:02:56.07" />
                    <SPLIT distance="225" swimtime="00:03:21.14" />
                    <SPLIT distance="250" swimtime="00:03:45.84" />
                    <SPLIT distance="275" swimtime="00:04:10.70" />
                    <SPLIT distance="300" swimtime="00:04:35.54" />
                    <SPLIT distance="325" swimtime="00:04:56.38" />
                    <SPLIT distance="350" swimtime="00:05:16.44" />
                    <SPLIT distance="375" swimtime="00:05:35.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="405" reactiontime="+91" swimtime="00:02:19.15" resultid="4042" lane="5" heatid="7062" entrytime="00:02:23.15">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.37" />
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                    <SPLIT distance="75" swimtime="00:00:49.74" />
                    <SPLIT distance="100" swimtime="00:01:07.76" />
                    <SPLIT distance="125" swimtime="00:01:25.51" />
                    <SPLIT distance="150" swimtime="00:01:43.77" />
                    <SPLIT distance="175" swimtime="00:02:02.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LUBLI" name="Lublin" nation="POL">
          <CONTACT name="Dobrowolski" />
          <ATHLETES>
            <ATHLETE birthdate="1984-01-01" firstname="Wojciech" gender="M" lastname="Dobrowolski" nation="POL" athleteid="4045">
              <RESULTS>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="4046" lane="5" heatid="6839" entrytime="00:01:06.84" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOCZE" name="MOSiR Częstochowa" nation="POL">
          <CONTACT name="Stachurski" />
          <ATHLETES>
            <ATHLETE birthdate="1969-01-01" firstname="Ireneusz" gender="M" lastname="Stachurski" nation="POL" athleteid="4048">
              <RESULTS>
                <RESULT eventid="1730" points="150" reactiontime="+90" swimtime="00:01:38.82" resultid="4053" heatid="7321" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.09" />
                    <SPLIT distance="50" swimtime="00:00:46.25" />
                    <SPLIT distance="75" swimtime="00:01:13.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="149" reactiontime="+89" swimtime="00:03:34.73" resultid="4050" lane="3" heatid="6882" entrytime="00:03:44.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.54" />
                    <SPLIT distance="50" swimtime="00:00:48.38" />
                    <SPLIT distance="75" swimtime="00:01:16.77" />
                    <SPLIT distance="100" swimtime="00:01:44.52" />
                    <SPLIT distance="125" swimtime="00:02:12.37" />
                    <SPLIT distance="150" swimtime="00:02:40.40" />
                    <SPLIT distance="175" swimtime="00:03:08.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="188" reactiontime="+117" swimtime="00:06:23.89" resultid="4051" lane="5" heatid="6901" entrytime="00:06:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.25" />
                    <SPLIT distance="50" swimtime="00:00:42.50" />
                    <SPLIT distance="75" swimtime="00:01:05.55" />
                    <SPLIT distance="100" swimtime="00:01:29.82" />
                    <SPLIT distance="125" swimtime="00:01:54.40" />
                    <SPLIT distance="150" swimtime="00:02:18.98" />
                    <SPLIT distance="175" swimtime="00:02:43.57" />
                    <SPLIT distance="200" swimtime="00:03:08.27" />
                    <SPLIT distance="225" swimtime="00:03:33.31" />
                    <SPLIT distance="250" swimtime="00:03:58.01" />
                    <SPLIT distance="275" swimtime="00:04:23.20" />
                    <SPLIT distance="300" swimtime="00:04:48.12" />
                    <SPLIT distance="325" swimtime="00:05:12.68" />
                    <SPLIT distance="350" swimtime="00:05:37.15" />
                    <SPLIT distance="375" swimtime="00:06:01.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" status="DNS" swimtime="00:00:00.00" resultid="4049" lane="5" heatid="6748" />
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="4052" lane="6" heatid="7056" entrytime="00:03:05.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MOOST" name="MOSiR Ostrowiec Świętokrzyski" nation="POL">
          <CONTACT name="Różalski" />
          <ATHLETES>
            <ATHLETE birthdate="1945-01-01" firstname="Józef" gender="M" lastname="Różalski" nation="POL" athleteid="4055">
              <RESULTS>
                <RESULT eventid="1764" points="313" reactiontime="+88" swimtime="00:00:31.33" resultid="4062" lane="1" heatid="7341" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="204" reactiontime="+87" swimtime="00:01:26.78" resultid="4056" lane="3" heatid="6734" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.24" />
                    <SPLIT distance="50" swimtime="00:00:41.50" />
                    <SPLIT distance="75" swimtime="00:01:07.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="269" reactiontime="+93" swimtime="00:01:12.81" resultid="4057" lane="1" heatid="6834" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.94" />
                    <SPLIT distance="50" swimtime="00:00:34.89" />
                    <SPLIT distance="75" swimtime="00:00:53.27" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1645" points="313" reactiontime="+87" swimtime="00:00:33.79" resultid="4061" heatid="7287" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="166" reactiontime="+97" swimtime="00:01:31.53" resultid="4059" lane="7" heatid="7018" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.54" />
                    <SPLIT distance="50" swimtime="00:00:43.10" />
                    <SPLIT distance="75" swimtime="00:01:09.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="173" swimtime="00:03:24.71" resultid="4060" lane="7" heatid="7074" entrytime="00:03:30.00" />
                <RESULT eventid="1273" points="118" reactiontime="+96" swimtime="00:03:48.20" resultid="4058" lane="5" heatid="6870" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.72" />
                    <SPLIT distance="50" swimtime="00:00:47.74" />
                    <SPLIT distance="75" swimtime="00:01:16.23" />
                    <SPLIT distance="100" swimtime="00:01:46.06" />
                    <SPLIT distance="125" swimtime="00:02:16.46" />
                    <SPLIT distance="150" swimtime="00:02:48.32" />
                    <SPLIT distance="175" swimtime="00:03:19.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="OLSTR" name="Olimpic Strawczyn" nation="POL">
          <CONTACT name="Śliwiński" />
          <ATHLETES>
            <ATHLETE birthdate="1952-01-01" firstname="Janusz" gender="M" lastname="Lipski" nation="POL" athleteid="4064">
              <RESULTS>
                <RESULT comment="Rekord Polski " eventid="1075" points="283" swimtime="00:11:38.14" resultid="4065" lane="4" heatid="6718" entrytime="00:12:30.20" />
                <RESULT eventid="1375" points="279" reactiontime="+113" swimtime="00:05:36.77" resultid="4067" heatid="6904" entrytime="00:05:52.16">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.60" />
                    <SPLIT distance="50" swimtime="00:00:37.85" />
                    <SPLIT distance="75" swimtime="00:00:58.61" />
                    <SPLIT distance="100" swimtime="00:01:19.60" />
                    <SPLIT distance="125" swimtime="00:01:41.08" />
                    <SPLIT distance="150" swimtime="00:02:02.63" />
                    <SPLIT distance="175" swimtime="00:02:24.30" />
                    <SPLIT distance="200" swimtime="00:02:46.05" />
                    <SPLIT distance="225" swimtime="00:03:07.37" />
                    <SPLIT distance="250" swimtime="00:03:29.19" />
                    <SPLIT distance="275" swimtime="00:03:50.23" />
                    <SPLIT distance="300" swimtime="00:04:11.78" />
                    <SPLIT distance="325" swimtime="00:04:33.66" />
                    <SPLIT distance="350" swimtime="00:04:55.35" />
                    <SPLIT distance="375" swimtime="00:05:16.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="261" reactiontime="+104" swimtime="00:02:41.06" resultid="4068" lane="4" heatid="7057" entrytime="00:02:50.15">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.39" />
                    <SPLIT distance="50" swimtime="00:00:36.60" />
                    <SPLIT distance="75" swimtime="00:00:56.79" />
                    <SPLIT distance="100" swimtime="00:01:17.69" />
                    <SPLIT distance="125" swimtime="00:01:38.83" />
                    <SPLIT distance="150" swimtime="00:02:00.59" />
                    <SPLIT distance="175" swimtime="00:02:21.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="282" reactiontime="+99" swimtime="00:01:11.70" resultid="4066" lane="2" heatid="6835" entrytime="00:01:12.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.25" />
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                    <SPLIT distance="75" swimtime="00:00:53.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" status="DNS" swimtime="00:00:00.00" resultid="4069" lane="4" heatid="7359" entrytime="00:07:24.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-01" firstname="Rafał" gender="M" lastname="Śliwiński" nation="POL" athleteid="4070">
              <RESULTS>
                <RESULT eventid="1273" points="115" reactiontime="+92" swimtime="00:03:49.79" resultid="4072" lane="1" heatid="6869">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.74" />
                    <SPLIT distance="50" swimtime="00:00:51.36" />
                    <SPLIT distance="75" swimtime="00:01:21.04" />
                    <SPLIT distance="100" swimtime="00:01:51.48" />
                    <SPLIT distance="125" swimtime="00:02:22.15" />
                    <SPLIT distance="150" swimtime="00:02:52.26" />
                    <SPLIT distance="175" swimtime="00:03:21.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="187" reactiontime="+89" swimtime="00:02:59.95" resultid="4073" lane="5" heatid="7056" entrytime="00:03:02.55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.86" />
                    <SPLIT distance="50" swimtime="00:00:37.87" />
                    <SPLIT distance="75" swimtime="00:00:59.10" />
                    <SPLIT distance="100" swimtime="00:01:21.99" />
                    <SPLIT distance="125" swimtime="00:01:45.46" />
                    <SPLIT distance="150" swimtime="00:02:10.46" />
                    <SPLIT distance="175" swimtime="00:02:36.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="183" reactiontime="+84" swimtime="00:01:30.03" resultid="4071" lane="5" heatid="6734" entrytime="00:01:28.55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.09" />
                    <SPLIT distance="50" swimtime="00:00:42.64" />
                    <SPLIT distance="75" swimtime="00:01:08.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="4075" lane="7" heatid="7342" entrytime="00:00:31.50" />
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="4074" heatid="7286" entrytime="00:00:34.60" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="OSWIE" name="Oświęcim" nation="POL">
          <CONTACT name="Dorywalski" />
          <ATHLETES>
            <ATHLETE birthdate="1961-01-01" firstname="Tomasz" gender="M" lastname="Dorywalski" nation="POL" athleteid="4077">
              <RESULTS>
                <RESULT eventid="1307" points="294" reactiontime="+64" swimtime="00:02:51.34" resultid="4078" lane="1" heatid="6885" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.80" />
                    <SPLIT distance="50" swimtime="00:00:38.82" />
                    <SPLIT distance="75" swimtime="00:00:59.41" />
                    <SPLIT distance="100" swimtime="00:01:20.65" />
                    <SPLIT distance="125" swimtime="00:01:42.46" />
                    <SPLIT distance="150" swimtime="00:02:05.02" />
                    <SPLIT distance="175" swimtime="00:02:28.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="319" reactiontime="+67" swimtime="00:00:35.79" resultid="4079" lane="8" heatid="7038" entrytime="00:00:36.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="309" reactiontime="+65" swimtime="00:01:17.68" resultid="4080" lane="8" heatid="7324" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.27" />
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                    <SPLIT distance="75" swimtime="00:00:57.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="STSZC" name="Szczecineckie Towarzystwo Pływackie Masters" nation="POL">
          <CONTACT name="Ludwiczak" />
          <ATHLETES>
            <ATHLETE birthdate="1937-01-01" firstname="Irena" gender="F" lastname="Filipowska" nation="POL" athleteid="4085">
              <RESULTS>
                <RESULT eventid="1222" points="41" swimtime="00:01:27.66" resultid="4086" lane="7" heatid="6848" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:42.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="24" reactiontime="+120" swimtime="00:07:09.01" resultid="4087" lane="5" heatid="6875" entrytime="00:07:24.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:47.92" />
                    <SPLIT distance="50" swimtime="00:01:41.15" />
                    <SPLIT distance="75" swimtime="00:02:36.90" />
                    <SPLIT distance="100" swimtime="00:03:31.57" />
                    <SPLIT distance="125" swimtime="00:04:27.82" />
                    <SPLIT distance="150" swimtime="00:05:22.96" />
                    <SPLIT distance="175" swimtime="00:06:19.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="26" swimtime="00:03:16.72" resultid="4089" lane="4" heatid="7312" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:44.71" />
                    <SPLIT distance="75" swimtime="00:02:23.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="14" swimtime="00:01:38.90" resultid="4090" lane="7" heatid="7328" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:46.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="31" reactiontime="+104" swimtime="00:01:27.48" resultid="4088" lane="2" heatid="7025" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:41.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-01-01" firstname="Krystyna" gender="F" lastname="Witkowska" nation="POL" athleteid="4091">
              <RESULTS>
                <RESULT eventid="1187" points="36" reactiontime="+121" swimtime="00:02:38.97" resultid="4092" lane="7" heatid="6822" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.10" />
                    <SPLIT distance="50" swimtime="00:01:14.43" />
                    <SPLIT distance="75" swimtime="00:01:56.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="38" reactiontime="+120" swimtime="00:05:39.41" resultid="4095" lane="5" heatid="7048" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.65" />
                    <SPLIT distance="50" swimtime="00:01:13.95" />
                    <SPLIT distance="75" swimtime="00:01:56.53" />
                    <SPLIT distance="100" swimtime="00:02:42.16" />
                    <SPLIT distance="125" swimtime="00:03:26.20" />
                    <SPLIT distance="150" swimtime="00:04:12.61" />
                    <SPLIT distance="175" swimtime="00:04:57.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="40" reactiontime="+111" swimtime="00:01:09.91" resultid="4097" lane="1" heatid="7328" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="34" reactiontime="+123" swimtime="00:01:32.87" resultid="4093" heatid="6848" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:42.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="22" reactiontime="+96" swimtime="00:01:37.94" resultid="4094" lane="6" heatid="7025" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:44.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="23" reactiontime="+89" swimtime="00:03:24.41" resultid="4096" lane="3" heatid="7312" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:45.36" />
                    <SPLIT distance="50" swimtime="00:01:41.28" />
                    <SPLIT distance="75" swimtime="00:02:33.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Barbara" gender="F" lastname="Jaczewska" nation="POL" athleteid="4098">
              <RESULTS>
                <RESULT eventid="1747" points="272" reactiontime="+97" swimtime="00:00:36.97" resultid="4105" lane="7" heatid="7332" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="259" reactiontime="+98" swimtime="00:01:22.93" resultid="4100" lane="5" heatid="6825" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.76" />
                    <SPLIT distance="50" swimtime="00:00:39.51" />
                    <SPLIT distance="75" swimtime="00:01:01.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="200" reactiontime="+95" swimtime="00:01:40.40" resultid="4099" lane="3" heatid="6725" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.05" />
                    <SPLIT distance="50" swimtime="00:00:46.25" />
                    <SPLIT distance="75" swimtime="00:01:16.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="198" reactiontime="+101" swimtime="00:06:54.00" resultid="4101" lane="5" heatid="6896" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.26" />
                    <SPLIT distance="50" swimtime="00:00:42.55" />
                    <SPLIT distance="75" swimtime="00:01:06.09" />
                    <SPLIT distance="100" swimtime="00:01:30.40" />
                    <SPLIT distance="125" swimtime="00:01:55.46" />
                    <SPLIT distance="150" swimtime="00:02:21.44" />
                    <SPLIT distance="175" swimtime="00:02:47.87" />
                    <SPLIT distance="200" swimtime="00:03:14.97" />
                    <SPLIT distance="225" swimtime="00:03:41.58" />
                    <SPLIT distance="250" swimtime="00:04:09.09" />
                    <SPLIT distance="275" swimtime="00:04:36.65" />
                    <SPLIT distance="300" swimtime="00:05:04.40" />
                    <SPLIT distance="325" swimtime="00:05:32.01" />
                    <SPLIT distance="350" swimtime="00:05:59.44" />
                    <SPLIT distance="375" swimtime="00:06:27.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="180" reactiontime="+69" swimtime="00:00:48.98" resultid="4102" heatid="7027" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1581" points="175" reactiontime="+100" swimtime="00:03:49.57" resultid="4103" lane="6" heatid="7069" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.90" />
                    <SPLIT distance="50" swimtime="00:00:52.46" />
                    <SPLIT distance="75" swimtime="00:01:22.18" />
                    <SPLIT distance="100" swimtime="00:01:51.73" />
                    <SPLIT distance="125" swimtime="00:02:25.41" />
                    <SPLIT distance="150" swimtime="00:02:58.51" />
                    <SPLIT distance="175" swimtime="00:03:24.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="188" reactiontime="+100" swimtime="00:01:53.57" resultid="4104" heatid="7297" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.34" />
                    <SPLIT distance="50" swimtime="00:00:54.63" />
                    <SPLIT distance="75" swimtime="00:01:23.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1933-01-01" firstname="Zbigniew" gender="M" lastname="Ludwiczak" nation="POL" athleteid="4106">
              <RESULTS>
                <RESULT eventid="1730" points="63" reactiontime="+100" swimtime="00:02:11.61" resultid="4113" heatid="7319" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.22" />
                    <SPLIT distance="50" swimtime="00:01:03.46" />
                    <SPLIT distance="75" swimtime="00:01:38.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="74" swimtime="00:18:10.49" resultid="4107" lane="4" heatid="6716" entrytime="00:18:02.00" />
                <RESULT eventid="1307" points="70" reactiontime="+94" swimtime="00:04:35.55" resultid="4108" lane="7" heatid="6881" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:33.49" />
                    <SPLIT distance="50" swimtime="00:01:06.56" />
                    <SPLIT distance="75" swimtime="00:01:40.37" />
                    <SPLIT distance="100" swimtime="00:02:15.42" />
                    <SPLIT distance="125" swimtime="00:02:51.55" />
                    <SPLIT distance="150" swimtime="00:03:27.85" />
                    <SPLIT distance="175" swimtime="00:04:02.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="82" swimtime="00:08:25.89" resultid="4109" lane="3" heatid="6899" entrytime="00:08:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.78" />
                    <SPLIT distance="50" swimtime="00:00:57.05" />
                    <SPLIT distance="75" swimtime="00:01:27.78" />
                    <SPLIT distance="100" swimtime="00:01:59.59" />
                    <SPLIT distance="125" swimtime="00:02:31.53" />
                    <SPLIT distance="150" swimtime="00:03:03.24" />
                    <SPLIT distance="175" swimtime="00:03:35.66" />
                    <SPLIT distance="200" swimtime="00:04:08.21" />
                    <SPLIT distance="225" swimtime="00:04:40.33" />
                    <SPLIT distance="250" swimtime="00:05:11.89" />
                    <SPLIT distance="275" swimtime="00:05:44.55" />
                    <SPLIT distance="300" swimtime="00:06:17.16" />
                    <SPLIT distance="325" swimtime="00:06:50.31" />
                    <SPLIT distance="350" swimtime="00:07:22.85" />
                    <SPLIT distance="375" swimtime="00:07:54.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="74" reactiontime="+89" swimtime="00:00:58.04" resultid="4110" lane="6" heatid="7033" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="76" swimtime="00:04:02.34" resultid="4111" lane="3" heatid="7054" entrytime="00:04:06.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.39" />
                    <SPLIT distance="50" swimtime="00:00:55.79" />
                    <SPLIT distance="75" swimtime="00:01:26.39" />
                    <SPLIT distance="100" swimtime="00:01:57.62" />
                    <SPLIT distance="125" swimtime="00:02:29.30" />
                    <SPLIT distance="150" swimtime="00:03:01.01" />
                    <SPLIT distance="175" swimtime="00:03:32.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="100" swimtime="00:02:06.78" resultid="4112" lane="5" heatid="7302" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.50" />
                    <SPLIT distance="50" swimtime="00:01:02.13" />
                    <SPLIT distance="75" swimtime="00:01:34.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-01-01" firstname="Ryszard" gender="M" lastname="Szwedowicz" nation="POL" athleteid="4114">
              <RESULTS>
                <RESULT eventid="1205" points="60" reactiontime="+122" swimtime="00:01:59.79" resultid="4116" lane="4" heatid="6830" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.72" />
                    <SPLIT distance="50" swimtime="00:00:53.13" />
                    <SPLIT distance="75" swimtime="00:01:25.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="46" reactiontime="+116" swimtime="00:04:45.75" resultid="4119" lane="2" heatid="7054" entrytime="00:04:46.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.29" />
                    <SPLIT distance="50" swimtime="00:00:55.43" />
                    <SPLIT distance="75" swimtime="00:01:29.68" />
                    <SPLIT distance="100" swimtime="00:02:08.47" />
                    <SPLIT distance="125" swimtime="00:02:46.73" />
                    <SPLIT distance="150" swimtime="00:03:28.10" />
                    <SPLIT distance="175" swimtime="00:04:07.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="84" reactiontime="+117" swimtime="00:02:13.99" resultid="4121" lane="6" heatid="7302" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.91" />
                    <SPLIT distance="50" swimtime="00:01:02.99" />
                    <SPLIT distance="75" swimtime="00:01:37.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="96" reactiontime="+126" swimtime="00:00:59.23" resultid="4117" lane="3" heatid="6854" entrytime="00:00:57.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.27" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Z 2" eventid="1109" reactiontime="+104" status="DSQ" swimtime="00:00:00.00" resultid="4115" lane="3" heatid="6730" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.49" />
                    <SPLIT distance="50" swimtime="00:01:09.56" />
                    <SPLIT distance="75" swimtime="00:01:49.06" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K 8" eventid="1411" reactiontime="+99" status="DSQ" swimtime="00:05:04.53" resultid="4118" lane="5" heatid="7002" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.53" />
                    <SPLIT distance="50" swimtime="00:01:01.83" />
                    <SPLIT distance="75" swimtime="00:01:37.98" />
                    <SPLIT distance="100" swimtime="00:02:17.88" />
                    <SPLIT distance="125" swimtime="00:03:00.71" />
                    <SPLIT distance="150" swimtime="00:03:43.03" />
                    <SPLIT distance="175" swimtime="00:04:25.66" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="M 10" eventid="1645" reactiontime="+118" status="DSQ" swimtime="00:00:00.00" resultid="4120" lane="7" heatid="7281" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:33.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-01-01" firstname="Ryszard" gender="M" lastname="Przelicki" nation="POL" athleteid="4122">
              <RESULTS>
                <RESULT eventid="1764" points="83" reactiontime="+112" swimtime="00:00:48.70" resultid="4126" lane="4" heatid="7336" entrytime="00:00:47.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="56" reactiontime="+129" swimtime="00:02:02.57" resultid="4123" lane="3" heatid="6830" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.20" />
                    <SPLIT distance="50" swimtime="00:00:53.76" />
                    <SPLIT distance="75" swimtime="00:01:25.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="4125" heatid="7281" entrytime="00:01:18.00" />
                <RESULT comment="K 8" eventid="1239" reactiontime="+141" status="DSQ" swimtime="00:01:09.23" resultid="4124" lane="1" heatid="6854" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-01-01" firstname="Mariusz" gender="M" lastname="Świąder" nation="POL" athleteid="4127">
              <RESULTS>
                <RESULT eventid="1564" points="286" reactiontime="+84" swimtime="00:02:36.18" resultid="4131" lane="4" heatid="7061" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.42" />
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                    <SPLIT distance="75" swimtime="00:00:51.38" />
                    <SPLIT distance="100" swimtime="00:01:10.91" />
                    <SPLIT distance="125" swimtime="00:01:30.97" />
                    <SPLIT distance="150" swimtime="00:01:52.12" />
                    <SPLIT distance="175" swimtime="00:02:14.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="243" reactiontime="+74" swimtime="00:00:39.18" resultid="4130" lane="1" heatid="7039" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="366" reactiontime="+82" swimtime="00:01:05.72" resultid="4129" heatid="6839" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.55" />
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                    <SPLIT distance="75" swimtime="00:00:47.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="264" reactiontime="+85" swimtime="00:01:19.69" resultid="4128" lane="1" heatid="6739" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.71" />
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                    <SPLIT distance="75" swimtime="00:00:58.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="339" reactiontime="+83" swimtime="00:00:32.91" resultid="4132" lane="6" heatid="7289" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="401" reactiontime="+81" swimtime="00:00:28.84" resultid="4133" lane="8" heatid="7346" entrytime="00:00:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="319" agemin="280" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1815" swimtime="00:05:12.12" resultid="7498" lane="3" heatid="7502">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:42.59" />
                    <SPLIT distance="50" swimtime="00:01:30.13" />
                    <SPLIT distance="75" swimtime="00:02:15.88" />
                    <SPLIT distance="100" swimtime="00:03:03.65" />
                    <SPLIT distance="125" swimtime="00:03:35.84" />
                    <SPLIT distance="150" swimtime="00:04:22.63" />
                    <SPLIT distance="175" swimtime="00:04:45.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4085" number="1" />
                    <RELAYPOSITION athleteid="4091" number="2" reactiontime="+107" />
                    <RELAYPOSITION athleteid="4114" number="3" reactiontime="+72" />
                    <RELAYPOSITION athleteid="4122" number="4" reactiontime="+115" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1615" swimtime="00:04:16.47" resultid="7267" lane="1" heatid="7441">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:43.29" />
                    <SPLIT distance="50" swimtime="00:01:30.37" />
                    <SPLIT distance="75" swimtime="00:02:03.32" />
                    <SPLIT distance="100" swimtime="00:02:40.40" />
                    <SPLIT distance="125" swimtime="00:03:03.15" />
                    <SPLIT distance="150" swimtime="00:03:29.61" />
                    <SPLIT distance="175" swimtime="00:03:51.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4085" number="1" />
                    <RELAYPOSITION athleteid="4091" number="2" reactiontime="+63" />
                    <RELAYPOSITION athleteid="4122" number="3" reactiontime="+27" />
                    <RELAYPOSITION athleteid="4114" number="4" reactiontime="+76" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SRODA" name="Środa Wlkp" nation="POL">
          <CONTACT name="Hańczyk" />
          <ATHLETES>
            <ATHLETE birthdate="1965-01-01" firstname="Jacek" gender="M" lastname="Hańczyk" nation="POL" athleteid="4135">
              <RESULTS>
                <RESULT eventid="1143" points="243" swimtime="00:23:20.91" resultid="4136" lane="8" heatid="6751" entrytime="00:23:15.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="JAROS" name="Jarosław" nation="POL">
          <CONTACT name="Jaroń" />
          <ATHLETES>
            <ATHLETE birthdate="1971-01-01" firstname="Tomasz" gender="M" lastname="Jaroń" nation="POL" athleteid="4138">
              <RESULTS>
                <RESULT eventid="1696" points="319" reactiontime="+70" swimtime="00:01:26.16" resultid="4144" lane="3" heatid="7306" entrytime="00:01:30.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.67" />
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                    <SPLIT distance="75" swimtime="00:01:03.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="178" reactiontime="+74" swimtime="00:03:19.01" resultid="4140" lane="5" heatid="6871" entrytime="00:03:22.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.84" />
                    <SPLIT distance="50" swimtime="00:00:40.06" />
                    <SPLIT distance="75" swimtime="00:01:03.07" />
                    <SPLIT distance="100" swimtime="00:01:27.85" />
                    <SPLIT distance="125" swimtime="00:01:54.39" />
                    <SPLIT distance="150" swimtime="00:02:22.68" />
                    <SPLIT distance="175" swimtime="00:02:51.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="295" reactiontime="+74" swimtime="00:03:11.52" resultid="4142" lane="3" heatid="7007" entrytime="00:03:15.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.14" />
                    <SPLIT distance="50" swimtime="00:00:41.90" />
                    <SPLIT distance="75" swimtime="00:01:05.59" />
                    <SPLIT distance="100" swimtime="00:01:30.19" />
                    <SPLIT distance="125" swimtime="00:01:55.42" />
                    <SPLIT distance="150" swimtime="00:02:20.36" />
                    <SPLIT distance="175" swimtime="00:02:45.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="223" reactiontime="+67" swimtime="00:06:41.67" resultid="4145" lane="6" heatid="7361" entrytime="00:06:45.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.80" />
                    <SPLIT distance="50" swimtime="00:00:39.41" />
                    <SPLIT distance="75" swimtime="00:01:03.12" />
                    <SPLIT distance="100" swimtime="00:01:28.89" />
                    <SPLIT distance="125" swimtime="00:01:58.61" />
                    <SPLIT distance="150" swimtime="00:02:26.23" />
                    <SPLIT distance="175" swimtime="00:02:53.82" />
                    <SPLIT distance="200" swimtime="00:03:22.33" />
                    <SPLIT distance="225" swimtime="00:03:48.82" />
                    <SPLIT distance="250" swimtime="00:04:15.77" />
                    <SPLIT distance="275" swimtime="00:04:42.46" />
                    <SPLIT distance="300" swimtime="00:05:10.00" />
                    <SPLIT distance="325" swimtime="00:05:32.83" />
                    <SPLIT distance="350" swimtime="00:05:55.38" />
                    <SPLIT distance="375" swimtime="00:06:18.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="261" reactiontime="+65" swimtime="00:05:44.34" resultid="4141" lane="7" heatid="6905" entrytime="00:05:45.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.63" />
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                    <SPLIT distance="75" swimtime="00:00:55.32" />
                    <SPLIT distance="100" swimtime="00:01:16.15" />
                    <SPLIT distance="125" swimtime="00:01:36.82" />
                    <SPLIT distance="150" swimtime="00:01:58.18" />
                    <SPLIT distance="175" swimtime="00:02:19.73" />
                    <SPLIT distance="200" swimtime="00:02:42.30" />
                    <SPLIT distance="225" swimtime="00:03:04.75" />
                    <SPLIT distance="250" swimtime="00:03:27.38" />
                    <SPLIT distance="275" swimtime="00:03:50.47" />
                    <SPLIT distance="300" swimtime="00:04:13.69" />
                    <SPLIT distance="325" swimtime="00:04:36.61" />
                    <SPLIT distance="350" swimtime="00:05:00.09" />
                    <SPLIT distance="375" swimtime="00:05:23.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="225" swimtime="00:12:33.90" resultid="4139" lane="3" heatid="6719" entrytime="00:12:15.10" />
                <RESULT eventid="1564" points="236" reactiontime="+73" swimtime="00:02:46.40" resultid="4143" lane="4" heatid="7058" entrytime="00:02:42.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.89" />
                    <SPLIT distance="50" swimtime="00:00:34.41" />
                    <SPLIT distance="75" swimtime="00:00:54.60" />
                    <SPLIT distance="100" swimtime="00:01:15.87" />
                    <SPLIT distance="125" swimtime="00:01:38.08" />
                    <SPLIT distance="150" swimtime="00:02:00.77" />
                    <SPLIT distance="175" swimtime="00:02:24.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WALBR" name="Wałbrzych" nation="POL">
          <CONTACT name="Maciejewski" />
          <ATHLETES>
            <ATHLETE birthdate="1981-01-01" firstname="Robert" gender="M" lastname="Maciejewski" nation="POL" athleteid="4147">
              <RESULTS>
                <RESULT eventid="1307" status="DNS" swimtime="00:00:00.00" resultid="4148" lane="4" heatid="6880" />
                <RESULT eventid="1411" status="DNS" swimtime="00:00:00.00" resultid="4149" lane="6" heatid="7002" />
                <RESULT eventid="1696" status="DNS" swimtime="00:00:00.00" resultid="4150" lane="3" heatid="7301" />
                <RESULT eventid="1730" status="DNS" swimtime="00:00:00.00" resultid="4151" lane="6" heatid="7318" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WOKUT" name="WOPR Kutno" nation="POL">
          <CONTACT name="From" />
          <ATHLETES>
            <ATHLETE birthdate="1932-01-01" firstname="Kazimierz" gender="M" lastname="From" nation="POL" athleteid="4153">
              <RESULTS>
                <RESULT eventid="1205" points="50" reactiontime="+121" swimtime="00:02:07.33" resultid="4155" lane="5" heatid="6829">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.17" />
                    <SPLIT distance="50" swimtime="00:00:58.09" />
                    <SPLIT distance="75" swimtime="00:01:32.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="54" reactiontime="+117" swimtime="00:00:55.99" resultid="4160" lane="8" heatid="7336">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="39" reactiontime="+122" swimtime="00:05:03.12" resultid="4158" lane="7" heatid="7054">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.04" />
                    <SPLIT distance="50" swimtime="00:01:02.43" />
                    <SPLIT distance="75" swimtime="00:01:38.71" />
                    <SPLIT distance="100" swimtime="00:02:17.69" />
                    <SPLIT distance="125" swimtime="00:02:58.49" />
                    <SPLIT distance="150" swimtime="00:03:40.97" />
                    <SPLIT distance="175" swimtime="00:04:25.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="29" reactiontime="+89" swimtime="00:06:09.98" resultid="4156" lane="3" heatid="6880">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:38.25" />
                    <SPLIT distance="50" swimtime="00:01:20.65" />
                    <SPLIT distance="75" swimtime="00:02:06.24" />
                    <SPLIT distance="100" swimtime="00:02:55.93" />
                    <SPLIT distance="125" swimtime="00:03:46.97" />
                    <SPLIT distance="150" swimtime="00:04:37.25" />
                    <SPLIT distance="175" swimtime="00:05:25.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="31" reactiontime="+97" swimtime="00:02:46.17" resultid="4159" lane="1" heatid="7318">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:36.47" />
                    <SPLIT distance="50" swimtime="00:01:17.11" />
                    <SPLIT distance="75" swimtime="00:02:01.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="37" reactiontime="+86" swimtime="00:01:13.26" resultid="4157" lane="7" heatid="7032">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:35.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" status="DNS" swimtime="00:00:00.00" resultid="4154" lane="3" heatid="6748" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WOZGI" name="WOPR Zgiersko-Łęczycki" nation="POL">
          <CONTACT name="Niedźwiedź" />
          <ATHLETES>
            <ATHLETE birthdate="1962-01-01" firstname="Ewa" gender="F" lastname="Stępień" nation="POL" athleteid="4162">
              <RESULTS>
                <RESULT eventid="1679" points="319" reactiontime="+78" swimtime="00:01:35.20" resultid="4167" lane="8" heatid="7300" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.07" />
                    <SPLIT distance="50" swimtime="00:00:45.40" />
                    <SPLIT distance="75" swimtime="00:01:09.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1581" points="254" reactiontime="+76" swimtime="00:03:22.75" resultid="4166" lane="3" heatid="7069" entrytime="00:03:16.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.07" />
                    <SPLIT distance="50" swimtime="00:00:43.38" />
                    <SPLIT distance="75" swimtime="00:01:10.34" />
                    <SPLIT distance="100" swimtime="00:01:37.81" />
                    <SPLIT distance="125" swimtime="00:02:05.53" />
                    <SPLIT distance="150" swimtime="00:02:32.76" />
                    <SPLIT distance="175" swimtime="00:02:59.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="321" reactiontime="+74" swimtime="00:00:34.99" resultid="4168" lane="6" heatid="7333" entrytime="00:00:33.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="361" reactiontime="+79" swimtime="00:00:42.55" resultid="4164" lane="7" heatid="6852" entrytime="00:00:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="229" reactiontime="+79" swimtime="00:06:34.51" resultid="4165" lane="7" heatid="6896" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.18" />
                    <SPLIT distance="50" swimtime="00:00:42.95" />
                    <SPLIT distance="75" swimtime="00:01:06.43" />
                    <SPLIT distance="100" swimtime="00:01:30.95" />
                    <SPLIT distance="125" swimtime="00:01:56.05" />
                    <SPLIT distance="150" swimtime="00:02:22.27" />
                    <SPLIT distance="175" swimtime="00:02:47.77" />
                    <SPLIT distance="200" swimtime="00:03:13.54" />
                    <SPLIT distance="225" swimtime="00:03:39.55" />
                    <SPLIT distance="250" swimtime="00:04:05.39" />
                    <SPLIT distance="275" swimtime="00:04:31.89" />
                    <SPLIT distance="300" swimtime="00:04:57.67" />
                    <SPLIT distance="325" swimtime="00:05:22.99" />
                    <SPLIT distance="350" swimtime="00:05:48.06" />
                    <SPLIT distance="375" swimtime="00:06:12.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="292" reactiontime="+77" swimtime="00:01:28.54" resultid="4163" lane="5" heatid="6727" entrytime="00:01:25.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.32" />
                    <SPLIT distance="50" swimtime="00:00:41.75" />
                    <SPLIT distance="75" swimtime="00:01:06.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-01" firstname="Urszula" gender="F" lastname="Mróz" nation="POL" athleteid="4169">
              <RESULTS>
                <RESULT eventid="1479" points="371" reactiontime="+72" swimtime="00:00:38.50" resultid="4173" lane="6" heatid="7030" entrytime="00:00:38.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="342" reactiontime="+86" swimtime="00:00:34.25" resultid="4175" lane="2" heatid="7333" entrytime="00:00:33.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="299" reactiontime="+90" swimtime="00:00:38.07" resultid="4174" heatid="7279" entrytime="00:00:36.25">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="268" reactiontime="+75" swimtime="00:03:14.07" resultid="4172" lane="6" heatid="6878" entrytime="00:03:15.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.70" />
                    <SPLIT distance="50" swimtime="00:00:44.57" />
                    <SPLIT distance="75" swimtime="00:01:08.00" />
                    <SPLIT distance="100" swimtime="00:01:32.71" />
                    <SPLIT distance="125" swimtime="00:01:57.93" />
                    <SPLIT distance="150" swimtime="00:02:23.65" />
                    <SPLIT distance="175" swimtime="00:02:49.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="284" reactiontime="+101" swimtime="00:01:20.40" resultid="4171" heatid="6826" entrytime="00:01:16.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.17" />
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                    <SPLIT distance="75" swimtime="00:01:00.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="297" reactiontime="+95" swimtime="00:01:28.05" resultid="4170" lane="3" heatid="6727" entrytime="00:01:25.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.03" />
                    <SPLIT distance="50" swimtime="00:00:39.33" />
                    <SPLIT distance="75" swimtime="00:01:06.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Mirosława" gender="F" lastname="Rajtar" nation="POL" athleteid="4176">
              <RESULTS>
                <RESULT eventid="1641" points="213" reactiontime="+94" swimtime="00:00:42.60" resultid="4182" lane="8" heatid="7278" entrytime="00:00:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1581" points="219" reactiontime="+93" swimtime="00:03:32.90" resultid="4181" heatid="7069" entrytime="00:03:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.78" />
                    <SPLIT distance="50" swimtime="00:00:45.27" />
                    <SPLIT distance="75" swimtime="00:01:11.91" />
                    <SPLIT distance="100" swimtime="00:01:39.44" />
                    <SPLIT distance="125" swimtime="00:02:10.52" />
                    <SPLIT distance="150" swimtime="00:02:42.60" />
                    <SPLIT distance="175" swimtime="00:03:08.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="245" reactiontime="+72" swimtime="00:00:44.22" resultid="4180" lane="5" heatid="7027" entrytime="00:00:46.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="272" reactiontime="+90" swimtime="00:01:21.59" resultid="4178" lane="1" heatid="6825" entrytime="00:01:22.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.91" />
                    <SPLIT distance="50" swimtime="00:00:37.89" />
                    <SPLIT distance="75" swimtime="00:00:59.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="238" reactiontime="+97" swimtime="00:01:34.76" resultid="4177" lane="1" heatid="6726" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.34" />
                    <SPLIT distance="50" swimtime="00:00:42.74" />
                    <SPLIT distance="75" swimtime="00:01:11.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="207" reactiontime="+92" swimtime="00:06:47.75" resultid="4179" lane="6" heatid="6895" entrytime="00:07:10.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.57" />
                    <SPLIT distance="50" swimtime="00:00:41.73" />
                    <SPLIT distance="75" swimtime="00:01:05.78" />
                    <SPLIT distance="100" swimtime="00:01:30.48" />
                    <SPLIT distance="125" swimtime="00:01:56.50" />
                    <SPLIT distance="150" swimtime="00:02:22.75" />
                    <SPLIT distance="175" swimtime="00:02:49.40" />
                    <SPLIT distance="200" swimtime="00:03:15.91" />
                    <SPLIT distance="225" swimtime="00:03:43.08" />
                    <SPLIT distance="250" swimtime="00:04:09.87" />
                    <SPLIT distance="275" swimtime="00:04:36.95" />
                    <SPLIT distance="300" swimtime="00:05:04.15" />
                    <SPLIT distance="325" swimtime="00:05:30.47" />
                    <SPLIT distance="350" swimtime="00:05:57.34" />
                    <SPLIT distance="375" swimtime="00:06:23.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="261" reactiontime="+96" swimtime="00:00:37.50" resultid="4183" lane="7" heatid="7331" entrytime="00:00:37.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Bogdan" gender="M" lastname="Wąsik" nation="POL" athleteid="4184">
              <RESULTS>
                <RESULT eventid="1239" points="333" reactiontime="+94" swimtime="00:00:39.21" resultid="4186" lane="7" heatid="6860" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="297" reactiontime="+90" swimtime="00:03:10.99" resultid="4188" lane="8" heatid="7008" entrytime="00:03:14.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.78" />
                    <SPLIT distance="50" swimtime="00:00:43.14" />
                    <SPLIT distance="75" swimtime="00:01:06.66" />
                    <SPLIT distance="100" swimtime="00:01:30.72" />
                    <SPLIT distance="125" swimtime="00:01:55.41" />
                    <SPLIT distance="150" swimtime="00:02:21.00" />
                    <SPLIT distance="175" swimtime="00:02:46.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="323" reactiontime="+94" swimtime="00:01:25.78" resultid="4190" lane="8" heatid="7308" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.94" />
                    <SPLIT distance="50" swimtime="00:00:41.21" />
                    <SPLIT distance="75" swimtime="00:01:03.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="199" reactiontime="+104" swimtime="00:06:57.53" resultid="4191" lane="7" heatid="7360" entrytime="00:07:17.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.32" />
                    <SPLIT distance="50" swimtime="00:00:44.86" />
                    <SPLIT distance="75" swimtime="00:01:09.90" />
                    <SPLIT distance="100" swimtime="00:01:36.03" />
                    <SPLIT distance="125" swimtime="00:02:03.37" />
                    <SPLIT distance="150" swimtime="00:02:31.62" />
                    <SPLIT distance="175" swimtime="00:02:59.80" />
                    <SPLIT distance="200" swimtime="00:03:27.88" />
                    <SPLIT distance="225" swimtime="00:03:53.47" />
                    <SPLIT distance="250" swimtime="00:04:18.76" />
                    <SPLIT distance="275" swimtime="00:04:44.07" />
                    <SPLIT distance="300" swimtime="00:05:11.30" />
                    <SPLIT distance="350" swimtime="00:06:57.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="165" reactiontime="+81" swimtime="00:03:27.50" resultid="4187" lane="5" heatid="6883" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.93" />
                    <SPLIT distance="50" swimtime="00:00:48.32" />
                    <SPLIT distance="75" swimtime="00:01:13.20" />
                    <SPLIT distance="100" swimtime="00:01:39.69" />
                    <SPLIT distance="125" swimtime="00:02:06.78" />
                    <SPLIT distance="150" swimtime="00:02:33.87" />
                    <SPLIT distance="175" swimtime="00:03:01.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="198" reactiontime="+96" swimtime="00:03:15.75" resultid="4189" lane="8" heatid="7075" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.53" />
                    <SPLIT distance="50" swimtime="00:00:40.84" />
                    <SPLIT distance="75" swimtime="00:01:06.30" />
                    <SPLIT distance="100" swimtime="00:01:32.66" />
                    <SPLIT distance="125" swimtime="00:01:57.49" />
                    <SPLIT distance="150" swimtime="00:02:22.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="203" reactiontime="+92" swimtime="00:01:27.01" resultid="4185" lane="8" heatid="6735" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.81" />
                    <SPLIT distance="50" swimtime="00:00:40.26" />
                    <SPLIT distance="75" swimtime="00:01:03.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="Roman" gender="M" lastname="Wiczel" nation="POL" athleteid="4192">
              <RESULTS>
                <RESULT eventid="1696" points="286" reactiontime="+88" swimtime="00:01:29.40" resultid="4195" heatid="7307" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.05" />
                    <SPLIT distance="50" swimtime="00:00:41.62" />
                    <SPLIT distance="75" swimtime="00:01:04.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="263" reactiontime="+91" swimtime="00:03:18.95" resultid="4194" heatid="7006" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.25" />
                    <SPLIT distance="50" swimtime="00:00:44.72" />
                    <SPLIT distance="75" swimtime="00:01:10.00" />
                    <SPLIT distance="100" swimtime="00:01:35.86" />
                    <SPLIT distance="125" swimtime="00:02:02.21" />
                    <SPLIT distance="150" swimtime="00:02:28.66" />
                    <SPLIT distance="175" swimtime="00:02:54.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="340" reactiontime="+85" swimtime="00:00:38.92" resultid="4193" lane="4" heatid="6859" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1922-01-01" firstname="Kazimierz" gender="M" lastname="Mrówczyński" nation="POL" athleteid="4196">
              <RESULTS>
                <RESULT eventid="1764" points="72" reactiontime="+92" swimtime="00:00:50.93" resultid="4201" lane="6" heatid="7336" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="45" reactiontime="+113" swimtime="00:04:47.93" resultid="4200" lane="5" heatid="7054" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.99" />
                    <SPLIT distance="50" swimtime="00:01:01.22" />
                    <SPLIT distance="75" swimtime="00:01:37.78" />
                    <SPLIT distance="100" swimtime="00:02:15.91" />
                    <SPLIT distance="125" swimtime="00:02:54.72" />
                    <SPLIT distance="150" swimtime="00:03:33.82" />
                    <SPLIT distance="175" swimtime="00:04:12.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="45" reactiontime="+87" swimtime="00:10:18.65" resultid="4199" lane="5" heatid="6899" entrytime="00:10:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.63" />
                    <SPLIT distance="50" swimtime="00:01:03.40" />
                    <SPLIT distance="75" swimtime="00:01:40.41" />
                    <SPLIT distance="100" swimtime="00:02:18.86" />
                    <SPLIT distance="125" swimtime="00:02:58.18" />
                    <SPLIT distance="150" swimtime="00:03:38.01" />
                    <SPLIT distance="175" swimtime="00:04:17.83" />
                    <SPLIT distance="200" swimtime="00:04:57.84" />
                    <SPLIT distance="225" swimtime="00:05:38.42" />
                    <SPLIT distance="250" swimtime="00:06:18.77" />
                    <SPLIT distance="275" swimtime="00:06:58.84" />
                    <SPLIT distance="300" swimtime="00:07:39.09" />
                    <SPLIT distance="325" swimtime="00:08:18.69" />
                    <SPLIT distance="350" swimtime="00:08:59.09" />
                    <SPLIT distance="375" swimtime="00:09:39.45" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1075" points="47" swimtime="00:21:06.69" resultid="4197" lane="3" heatid="6716" entrytime="00:21:00.00" />
                <RESULT eventid="1205" points="47" reactiontime="+128" swimtime="00:02:10.21" resultid="4198" lane="5" heatid="6830" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.05" />
                    <SPLIT distance="50" swimtime="00:00:59.21" />
                    <SPLIT distance="75" swimtime="00:00:47.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Włodzimierz" gender="M" lastname="Przytulski" nation="POL" athleteid="4202">
              <RESULTS>
                <RESULT eventid="1462" points="269" reactiontime="+85" swimtime="00:01:18.03" resultid="4206" lane="8" heatid="7020" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.51" />
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                    <SPLIT distance="75" swimtime="00:00:55.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="342" reactiontime="+90" swimtime="00:01:07.27" resultid="4204" lane="3" heatid="6838" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.20" />
                    <SPLIT distance="50" swimtime="00:00:31.93" />
                    <SPLIT distance="75" swimtime="00:00:49.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="355" reactiontime="+79" swimtime="00:00:32.41" resultid="4208" lane="1" heatid="7288" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="277" reactiontime="+74" swimtime="00:01:18.43" resultid="4203" heatid="6738" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.24" />
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                    <SPLIT distance="75" swimtime="00:01:00.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="4205" heatid="6872" entrytime="00:03:15.00" />
                <RESULT eventid="1496" status="DNS" swimtime="00:00:00.00" resultid="4207" lane="3" heatid="7037" entrytime="00:00:37.00" />
                <RESULT eventid="1730" status="DNS" swimtime="00:00:00.00" resultid="4209" lane="3" heatid="7322" entrytime="00:01:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Mateusz" gender="M" lastname="Sass" nation="POL" athleteid="4210">
              <RESULTS>
                <RESULT eventid="1798" points="449" reactiontime="+74" swimtime="00:05:18.43" resultid="4216" lane="1" heatid="7364" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.61" />
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                    <SPLIT distance="75" swimtime="00:00:48.21" />
                    <SPLIT distance="100" swimtime="00:01:07.40" />
                    <SPLIT distance="125" swimtime="00:01:29.07" />
                    <SPLIT distance="150" swimtime="00:01:50.05" />
                    <SPLIT distance="175" swimtime="00:02:11.08" />
                    <SPLIT distance="200" swimtime="00:02:32.37" />
                    <SPLIT distance="225" swimtime="00:02:54.75" />
                    <SPLIT distance="250" swimtime="00:03:17.38" />
                    <SPLIT distance="275" swimtime="00:03:39.90" />
                    <SPLIT distance="300" swimtime="00:04:02.79" />
                    <SPLIT distance="325" swimtime="00:04:22.65" />
                    <SPLIT distance="350" swimtime="00:04:41.56" />
                    <SPLIT distance="375" swimtime="00:05:00.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="480" reactiontime="+78" swimtime="00:02:25.82" resultid="4214" lane="4" heatid="7079" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.30" />
                    <SPLIT distance="50" swimtime="00:00:29.48" />
                    <SPLIT distance="75" swimtime="00:00:48.95" />
                    <SPLIT distance="100" swimtime="00:01:07.70" />
                    <SPLIT distance="125" swimtime="00:01:28.90" />
                    <SPLIT distance="150" swimtime="00:01:50.09" />
                    <SPLIT distance="175" swimtime="00:02:08.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="357" reactiontime="+84" swimtime="00:02:37.90" resultid="4212" lane="6" heatid="6873" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.98" />
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                    <SPLIT distance="75" swimtime="00:00:49.17" />
                    <SPLIT distance="100" swimtime="00:01:08.38" />
                    <SPLIT distance="125" swimtime="00:01:29.29" />
                    <SPLIT distance="150" swimtime="00:01:50.93" />
                    <SPLIT distance="175" swimtime="00:02:14.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="479" swimtime="00:01:05.33" resultid="4211" lane="7" heatid="6745" entrytime="00:01:04.00" />
                <RESULT eventid="1645" points="502" reactiontime="+117" swimtime="00:00:28.88" resultid="4215" lane="5" heatid="7293" entrytime="00:00:27.49">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" status="DNS" swimtime="00:00:00.00" resultid="4213" lane="6" heatid="7019" entrytime="00:01:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-01" firstname="Tomasz" gender="M" lastname="Niedźwiedź" nation="POL" athleteid="4217">
              <RESULTS>
                <RESULT eventid="1798" points="188" reactiontime="+93" swimtime="00:07:05.37" resultid="4223" lane="8" heatid="7360" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.98" />
                    <SPLIT distance="50" swimtime="00:00:47.73" />
                    <SPLIT distance="75" swimtime="00:01:14.43" />
                    <SPLIT distance="100" swimtime="00:01:41.48" />
                    <SPLIT distance="125" swimtime="00:02:10.60" />
                    <SPLIT distance="150" swimtime="00:02:38.75" />
                    <SPLIT distance="175" swimtime="00:03:07.25" />
                    <SPLIT distance="200" swimtime="00:03:35.24" />
                    <SPLIT distance="225" swimtime="00:04:03.35" />
                    <SPLIT distance="250" swimtime="00:04:31.40" />
                    <SPLIT distance="275" swimtime="00:05:00.43" />
                    <SPLIT distance="300" swimtime="00:05:29.20" />
                    <SPLIT distance="325" swimtime="00:05:54.54" />
                    <SPLIT distance="350" swimtime="00:06:18.96" />
                    <SPLIT distance="375" swimtime="00:06:42.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="177" reactiontime="+92" swimtime="00:03:23.32" resultid="4221" lane="1" heatid="7074" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.53" />
                    <SPLIT distance="50" swimtime="00:00:43.48" />
                    <SPLIT distance="75" swimtime="00:01:11.79" />
                    <SPLIT distance="100" swimtime="00:01:40.69" />
                    <SPLIT distance="125" swimtime="00:02:08.74" />
                    <SPLIT distance="150" swimtime="00:02:36.66" />
                    <SPLIT distance="175" swimtime="00:03:00.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="132" reactiontime="+101" swimtime="00:03:39.86" resultid="4219" lane="3" heatid="6870" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.92" />
                    <SPLIT distance="50" swimtime="00:00:49.15" />
                    <SPLIT distance="75" swimtime="00:01:16.46" />
                    <SPLIT distance="100" swimtime="00:01:45.24" />
                    <SPLIT distance="125" swimtime="00:02:14.49" />
                    <SPLIT distance="150" swimtime="00:02:43.74" />
                    <SPLIT distance="175" swimtime="00:03:12.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="190" reactiontime="+96" swimtime="00:01:28.85" resultid="4218" lane="3" heatid="6733" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.21" />
                    <SPLIT distance="50" swimtime="00:00:42.59" />
                    <SPLIT distance="75" swimtime="00:01:08.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" status="DNS" swimtime="00:00:00.00" resultid="4220" lane="3" heatid="7016" entrytime="00:01:40.00" />
                <RESULT eventid="1645" reactiontime="+105" status="DNS" swimtime="00:00:00.00" resultid="4222" lane="7" heatid="7283" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Tadeusz" gender="M" lastname="Obiedziński" nation="POL" athleteid="4224">
              <RESULTS>
                <RESULT eventid="1696" points="257" reactiontime="+100" swimtime="00:01:32.54" resultid="4228" lane="8" heatid="7306" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.42" />
                    <SPLIT distance="50" swimtime="00:00:42.44" />
                    <SPLIT distance="75" swimtime="00:01:07.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="306" reactiontime="+93" swimtime="00:00:40.30" resultid="4226" lane="3" heatid="6857" entrytime="00:00:42.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="188" reactiontime="+100" swimtime="00:01:29.21" resultid="4225" lane="2" heatid="6733" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.35" />
                    <SPLIT distance="50" swimtime="00:00:41.32" />
                    <SPLIT distance="75" swimtime="00:01:05.73" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K 11" eventid="1411" reactiontime="+113" status="DSQ" swimtime="00:00:00.00" resultid="4227" lane="8" heatid="7006" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.84" />
                    <SPLIT distance="50" swimtime="00:00:46.87" />
                    <SPLIT distance="75" swimtime="00:01:13.96" />
                    <SPLIT distance="100" swimtime="00:01:41.23" />
                    <SPLIT distance="125" swimtime="00:02:09.10" />
                    <SPLIT distance="150" swimtime="00:02:37.42" />
                    <SPLIT distance="175" swimtime="00:03:05.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Krzysztof" gender="M" lastname="Bednarek" nation="POL" athleteid="5426">
              <RESULTS>
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="5427" lane="1" heatid="6732" entrytime="00:01:40.00" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="5428" lane="7" heatid="6834" entrytime="00:01:18.00" />
                <RESULT eventid="1375" status="DNS" swimtime="00:00:00.00" resultid="5429" lane="7" heatid="6902" entrytime="00:06:20.00" />
                <RESULT eventid="1598" status="DNS" swimtime="00:00:00.00" resultid="5430" lane="2" heatid="7074" entrytime="00:03:20.00" />
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="5431" lane="1" heatid="7284" entrytime="00:00:37.00" />
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="5432" lane="5" heatid="7340" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="BIWAR" name="UKS G-8 Bielany" nation="POL">
          <CONTACT name="Obukowicz Marcin" phone="601 066 343" />
          <ATHLETES>
            <ATHLETE birthdate="1990-06-24" firstname="Michał" gender="M" lastname="Choiński" nation="POL" athleteid="4232">
              <RESULTS>
                <RESULT eventid="1730" points="509" reactiontime="+70" swimtime="00:01:05.80" resultid="4236" lane="4" heatid="7326" entrytime="00:00:59.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.73" />
                    <SPLIT distance="50" swimtime="00:00:30.81" />
                    <SPLIT distance="75" swimtime="00:00:48.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="574" reactiontime="+73" swimtime="00:00:29.43" resultid="4234" lane="4" heatid="7043" entrytime="00:00:27.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="638" reactiontime="+68" swimtime="00:00:26.67" resultid="4235" lane="5" heatid="7294" entrytime="00:00:25.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="574" reactiontime="+71" swimtime="00:00:56.59" resultid="4233" lane="3" heatid="6846" entrytime="00:00:54.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.82" />
                    <SPLIT distance="50" swimtime="00:00:27.54" />
                    <SPLIT distance="75" swimtime="00:00:42.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DEINO" name="Delfin Inowrocław" nation="POL" region="KUJ">
          <CONTACT state="KUJ" />
          <ATHLETES>
            <ATHLETE birthdate="1965-07-15" firstname="Jarosław" gender="M" lastname="Molenda" nation="POL" license="S01202200044" athleteid="4238">
              <RESULTS>
                <RESULT eventid="1239" points="375" reactiontime="+81" swimtime="00:00:37.68" resultid="4239" lane="4" heatid="6861" entrytime="00:00:37.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-10-21" firstname="Wiesław" gender="M" lastname="Chabecki" nation="POL" license="S01202200045" athleteid="4240">
              <RESULTS>
                <RESULT eventid="1496" points="137" reactiontime="+89" swimtime="00:00:47.36" resultid="4241" lane="5" heatid="7034" entrytime="00:00:48.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="192" reactiontime="+110" swimtime="00:00:36.88" resultid="4242" heatid="7338" entrytime="00:00:37.48">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-01-28" firstname="Krzysztof" gender="M" lastname="Derkowski" nation="POL" license="S01202200043" athleteid="4243">
              <RESULTS>
                <RESULT eventid="1645" points="236" reactiontime="+76" swimtime="00:00:37.11" resultid="4247" lane="5" heatid="7284" entrytime="00:00:36.92">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="272" reactiontime="+80" swimtime="00:00:32.84" resultid="4248" lane="1" heatid="7340" entrytime="00:00:33.66">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="222" reactiontime="+84" swimtime="00:01:17.64" resultid="4245" heatid="6834" entrytime="00:01:18.09">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.73" />
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                    <SPLIT distance="75" swimtime="00:00:55.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="252" reactiontime="+84" swimtime="00:00:43.01" resultid="4246" lane="6" heatid="6857" entrytime="00:00:42.92">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="177" reactiontime="+82" swimtime="00:01:31.01" resultid="4244" lane="5" heatid="6733" entrytime="00:01:31.02">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.34" />
                    <SPLIT distance="50" swimtime="00:00:41.77" />
                    <SPLIT distance="75" swimtime="00:01:08.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-08-07" firstname="Tomasz" gender="M" lastname="Glubiak" nation="POL" license="S01202200046" athleteid="4249">
              <RESULTS>
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="4250" lane="2" heatid="7340" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1177" status="DNS" swimtime="00:00:00.00" resultid="4251" lane="1" heatid="6808" entrytime="00:02:16.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4249" number="1" />
                    <RELAYPOSITION athleteid="4240" number="2" />
                    <RELAYPOSITION athleteid="4243" number="3" />
                    <RELAYPOSITION athleteid="4238" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1341" points="222" reactiontime="+74" swimtime="00:02:37.62" resultid="4252" heatid="6986" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.48" />
                    <SPLIT distance="50" swimtime="00:00:48.22" />
                    <SPLIT distance="75" swimtime="00:01:05.56" />
                    <SPLIT distance="100" swimtime="00:01:26.54" />
                    <SPLIT distance="125" swimtime="00:01:44.10" />
                    <SPLIT distance="150" swimtime="00:02:03.99" />
                    <SPLIT distance="175" swimtime="00:02:19.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4240" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="4238" number="2" reactiontime="+52" />
                    <RELAYPOSITION athleteid="4243" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="4249" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1177" points="262" reactiontime="+97" swimtime="00:02:15.46" resultid="6668" lane="5" heatid="6807">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.83" />
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                    <SPLIT distance="75" swimtime="00:00:52.22" />
                    <SPLIT distance="100" swimtime="00:01:11.51" />
                    <SPLIT distance="125" swimtime="00:01:27.94" />
                    <SPLIT distance="150" swimtime="00:01:45.84" />
                    <SPLIT distance="175" swimtime="00:01:59.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4249" number="1" reactiontime="+97" />
                    <RELAYPOSITION athleteid="4240" number="2" reactiontime="+69" />
                    <RELAYPOSITION athleteid="4243" number="3" reactiontime="+42" />
                    <RELAYPOSITION athleteid="4238" number="4" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="UCWAR" name="UCSiR Warszawa" nation="POL" region="MAZ">
          <CONTACT city="Warszawa" name="Michał Nowak" />
          <ATHLETES>
            <ATHLETE birthdate="1985-05-26" firstname="Urszula" gender="F" lastname="Bielawska" nation="POL" athleteid="4261">
              <RESULTS>
                <RESULT eventid="1679" points="278" reactiontime="+96" swimtime="00:01:39.66" resultid="4267" lane="2" heatid="7298" entrytime="00:01:44.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.21" />
                    <SPLIT distance="50" swimtime="00:00:47.45" />
                    <SPLIT distance="75" swimtime="00:01:13.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1058" points="285" swimtime="00:12:30.48" resultid="4262" lane="4" heatid="6714" entrytime="00:12:30.00" />
                <RESULT eventid="1222" points="301" reactiontime="+83" swimtime="00:00:45.21" resultid="4263" lane="5" heatid="6851" entrytime="00:00:44.88">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="344" reactiontime="+84" swimtime="00:02:43.79" resultid="4266" heatid="7052" entrytime="00:02:46.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.82" />
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                    <SPLIT distance="75" swimtime="00:00:58.20" />
                    <SPLIT distance="100" swimtime="00:01:18.87" />
                    <SPLIT distance="125" swimtime="00:01:40.40" />
                    <SPLIT distance="150" swimtime="00:02:02.84" />
                    <SPLIT distance="175" swimtime="00:02:23.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="389" reactiontime="+85" swimtime="00:00:32.81" resultid="4268" lane="8" heatid="7334" entrytime="00:00:32.61">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="234" reactiontime="+90" swimtime="00:00:44.88" resultid="4265" lane="1" heatid="7028" entrytime="00:00:43.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="328" reactiontime="+92" swimtime="00:05:50.15" resultid="4264" lane="5" heatid="6897" entrytime="00:05:46.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.25" />
                    <SPLIT distance="50" swimtime="00:00:38.11" />
                    <SPLIT distance="75" swimtime="00:00:58.69" />
                    <SPLIT distance="100" swimtime="00:01:19.93" />
                    <SPLIT distance="125" swimtime="00:01:41.53" />
                    <SPLIT distance="150" swimtime="00:02:03.80" />
                    <SPLIT distance="175" swimtime="00:02:25.71" />
                    <SPLIT distance="200" swimtime="00:02:47.91" />
                    <SPLIT distance="225" swimtime="00:03:10.62" />
                    <SPLIT distance="250" swimtime="00:03:33.03" />
                    <SPLIT distance="275" swimtime="00:03:55.79" />
                    <SPLIT distance="300" swimtime="00:04:18.83" />
                    <SPLIT distance="325" swimtime="00:04:42.24" />
                    <SPLIT distance="350" swimtime="00:05:05.83" />
                    <SPLIT distance="375" swimtime="00:05:28.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-09-16" firstname="Monika" gender="F" lastname="Kuryłowicz" nation="POL" athleteid="4269">
              <RESULTS>
                <RESULT comment="Rekord Polski " eventid="1126" points="207" swimtime="00:26:32.27" resultid="4270" heatid="6747" entrytime="00:27:00.00" />
                <RESULT eventid="1547" points="230" reactiontime="+88" swimtime="00:03:07.15" resultid="4273" lane="3" heatid="7050" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.60" />
                    <SPLIT distance="50" swimtime="00:00:41.99" />
                    <SPLIT distance="75" swimtime="00:01:05.55" />
                    <SPLIT distance="100" swimtime="00:01:29.85" />
                    <SPLIT distance="125" swimtime="00:01:54.55" />
                    <SPLIT distance="150" swimtime="00:02:19.49" />
                    <SPLIT distance="175" swimtime="00:02:44.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="228" reactiontime="+90" swimtime="00:06:34.95" resultid="4272" lane="8" heatid="6896" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.98" />
                    <SPLIT distance="50" swimtime="00:00:43.28" />
                    <SPLIT distance="75" swimtime="00:01:07.80" />
                    <SPLIT distance="100" swimtime="00:01:32.24" />
                    <SPLIT distance="125" swimtime="00:01:57.89" />
                    <SPLIT distance="150" swimtime="00:02:23.14" />
                    <SPLIT distance="175" swimtime="00:02:49.34" />
                    <SPLIT distance="200" swimtime="00:03:15.00" />
                    <SPLIT distance="225" swimtime="00:03:41.05" />
                    <SPLIT distance="250" swimtime="00:04:06.61" />
                    <SPLIT distance="275" swimtime="00:04:33.00" />
                    <SPLIT distance="300" swimtime="00:04:58.51" />
                    <SPLIT distance="325" swimtime="00:05:24.62" />
                    <SPLIT distance="350" swimtime="00:05:49.62" />
                    <SPLIT distance="375" swimtime="00:06:13.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="269" reactiontime="+81" swimtime="00:00:37.10" resultid="4274" lane="2" heatid="7331" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="244" reactiontime="+86" swimtime="00:01:24.59" resultid="4271" lane="8" heatid="6825" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.33" />
                    <SPLIT distance="50" swimtime="00:00:39.88" />
                    <SPLIT distance="75" swimtime="00:01:02.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-05-26" firstname="Małgorzata" gender="F" lastname="Kotańska" nation="POL" athleteid="4275">
              <RESULTS>
                <RESULT eventid="1409" points="291" reactiontime="+98" swimtime="00:03:31.48" resultid="4279" lane="7" heatid="7000" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.13" />
                    <SPLIT distance="50" swimtime="00:00:47.37" />
                    <SPLIT distance="75" swimtime="00:01:13.84" />
                    <SPLIT distance="100" swimtime="00:01:41.38" />
                    <SPLIT distance="125" swimtime="00:02:09.12" />
                    <SPLIT distance="150" swimtime="00:02:37.21" />
                    <SPLIT distance="175" swimtime="00:03:04.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="293" reactiontime="+89" swimtime="00:01:37.89" resultid="4281" lane="8" heatid="7299" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.57" />
                    <SPLIT distance="50" swimtime="00:00:46.21" />
                    <SPLIT distance="75" swimtime="00:01:11.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="325" reactiontime="+90" swimtime="00:00:44.06" resultid="4277" lane="8" heatid="6852" entrytime="00:00:44.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="220" reactiontime="+84" swimtime="00:00:45.83" resultid="4280" lane="8" heatid="7028" entrytime="00:00:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="247" reactiontime="+77" swimtime="00:00:38.18" resultid="4282" lane="4" heatid="7330" entrytime="00:00:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="190" swimtime="00:06:59.68" resultid="4278" lane="1" heatid="6895" entrytime="00:07:15.00" />
                <RESULT eventid="1092" points="224" reactiontime="+92" swimtime="00:01:36.81" resultid="4276" lane="3" heatid="6726" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.52" />
                    <SPLIT distance="50" swimtime="00:00:47.22" />
                    <SPLIT distance="75" swimtime="00:01:13.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-04-10" firstname="Andrzej" gender="M" lastname="Rubaszkiewicz" nation="POL" athleteid="4290">
              <RESULTS>
                <RESULT eventid="1764" points="392" reactiontime="+81" swimtime="00:00:29.06" resultid="4297" lane="7" heatid="7346" entrytime="00:00:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="312" reactiontime="+81" swimtime="00:00:33.84" resultid="4296" lane="2" heatid="7287" entrytime="00:00:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="269" reactiontime="+76" swimtime="00:00:37.89" resultid="4294" heatid="7038" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="245" reactiontime="+87" swimtime="00:01:21.65" resultid="4291" lane="4" heatid="6736" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.35" />
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                    <SPLIT distance="75" swimtime="00:01:02.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="344" reactiontime="+70" swimtime="00:01:07.09" resultid="4292" lane="1" heatid="6840" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.40" />
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                    <SPLIT distance="75" swimtime="00:00:49.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="287" reactiontime="+87" swimtime="00:00:41.17" resultid="4293" heatid="6859" entrytime="00:00:40.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" status="DNS" swimtime="00:00:00.00" resultid="4295" lane="7" heatid="7076" entrytime="00:03:06.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-01-23" firstname="Michał" gender="M" lastname="Rybarczyk" nation="POL" athleteid="4298">
              <RESULTS>
                <RESULT eventid="1645" points="335" reactiontime="+83" swimtime="00:00:33.04" resultid="4303" lane="7" heatid="7287" entrytime="00:00:33.99">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="186" reactiontime="+78" swimtime="00:00:42.81" resultid="4301" lane="7" heatid="7036" entrytime="00:00:43.12">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="292" reactiontime="+83" swimtime="00:02:35.04" resultid="4302" lane="1" heatid="7060" entrytime="00:02:39.04">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.02" />
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                    <SPLIT distance="75" swimtime="00:00:54.09" />
                    <SPLIT distance="100" swimtime="00:01:13.60" />
                    <SPLIT distance="125" swimtime="00:01:34.66" />
                    <SPLIT distance="150" swimtime="00:01:55.65" />
                    <SPLIT distance="175" swimtime="00:02:16.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="391" reactiontime="+79" swimtime="00:00:29.09" resultid="4304" lane="1" heatid="7346" entrytime="00:00:28.99">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="365" reactiontime="+82" swimtime="00:01:05.81" resultid="4299" lane="4" heatid="6838" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.62" />
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                    <SPLIT distance="75" swimtime="00:00:48.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" status="DNS" swimtime="00:00:00.00" resultid="4300" lane="2" heatid="6904" entrytime="00:05:49.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1615" status="DNS" swimtime="00:00:00.00" resultid="4305" lane="3" heatid="7442" entrytime="00:02:09.00" />
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" name="UCSiR Warszawa 1" number="2">
              <RESULTS>
                <RESULT eventid="1815" status="DNS" swimtime="00:00:00.00" resultid="4306" lane="2" heatid="7503" entrytime="00:02:28.00" />
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="PIKON" name="UKS Piątka Konstantynów" nation="POL" region="LOD">
          <CONTACT email="tomaszkotus@tlen.pl" name="Kotus" phone="603820602" />
          <ATHLETES>
            <ATHLETE birthdate="1979-09-09" firstname="Marcin" gender="M" lastname="Grabarczyk" nation="POL" athleteid="4309">
              <RESULTS>
                <RESULT eventid="1143" points="337" swimtime="00:20:55.90" resultid="4310" lane="5" heatid="6752" entrytime="00:19:37.77" />
                <RESULT eventid="1598" points="362" reactiontime="+79" swimtime="00:02:40.18" resultid="4314" lane="8" heatid="7078" entrytime="00:02:47.77">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.89" />
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                    <SPLIT distance="75" swimtime="00:00:54.22" />
                    <SPLIT distance="100" swimtime="00:01:13.97" />
                    <SPLIT distance="125" swimtime="00:01:38.10" />
                    <SPLIT distance="150" swimtime="00:02:02.58" />
                    <SPLIT distance="175" swimtime="00:02:22.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="381" reactiontime="+78" swimtime="00:05:03.54" resultid="4312" lane="3" heatid="6908" entrytime="00:04:47.77">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.22" />
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                    <SPLIT distance="75" swimtime="00:00:50.24" />
                    <SPLIT distance="100" swimtime="00:01:08.60" />
                    <SPLIT distance="125" swimtime="00:01:27.04" />
                    <SPLIT distance="150" swimtime="00:01:46.38" />
                    <SPLIT distance="175" swimtime="00:02:05.37" />
                    <SPLIT distance="200" swimtime="00:02:25.07" />
                    <SPLIT distance="225" swimtime="00:02:43.98" />
                    <SPLIT distance="250" swimtime="00:03:04.04" />
                    <SPLIT distance="275" swimtime="00:03:23.77" />
                    <SPLIT distance="300" swimtime="00:03:43.96" />
                    <SPLIT distance="325" swimtime="00:04:04.24" />
                    <SPLIT distance="350" swimtime="00:04:24.40" />
                    <SPLIT distance="375" swimtime="00:04:44.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="199" reactiontime="+85" swimtime="00:03:11.84" resultid="4311" lane="5" heatid="6873" entrytime="00:02:47.77">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.51" />
                    <SPLIT distance="50" swimtime="00:00:34.41" />
                    <SPLIT distance="75" swimtime="00:00:54.03" />
                    <SPLIT distance="100" swimtime="00:01:15.73" />
                    <SPLIT distance="125" swimtime="00:01:42.90" />
                    <SPLIT distance="150" swimtime="00:02:13.24" />
                    <SPLIT distance="175" swimtime="00:02:42.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="378" reactiontime="+79" swimtime="00:00:31.73" resultid="4315" heatid="7291" entrytime="00:00:29.77">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="434" reactiontime="+77" swimtime="00:00:28.09" resultid="4316" heatid="7349" entrytime="00:00:27.77">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" status="DNS" swimtime="00:00:00.00" resultid="4313" lane="3" heatid="7020" entrytime="00:01:13.77" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-09-09" firstname="Jakub" gender="M" lastname="Karczmarczyk" nation="POL" athleteid="4317">
              <RESULTS>
                <RESULT eventid="1696" points="371" reactiontime="+86" swimtime="00:01:21.96" resultid="4322" lane="3" heatid="7310" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.79" />
                    <SPLIT distance="50" swimtime="00:00:37.45" />
                    <SPLIT distance="75" swimtime="00:00:59.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="281" reactiontime="+79" swimtime="00:02:53.94" resultid="4320" lane="2" heatid="6886" entrytime="00:02:38.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.09" />
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                    <SPLIT distance="75" swimtime="00:00:59.42" />
                    <SPLIT distance="100" swimtime="00:01:21.98" />
                    <SPLIT distance="125" swimtime="00:01:45.19" />
                    <SPLIT distance="150" swimtime="00:02:08.84" />
                    <SPLIT distance="175" swimtime="00:02:31.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="378" reactiontime="+70" swimtime="00:00:33.83" resultid="4321" lane="3" heatid="7042" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="337" reactiontime="+89" swimtime="00:01:13.49" resultid="4318" lane="6" heatid="6741" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.26" />
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                    <SPLIT distance="75" swimtime="00:00:54.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="436" reactiontime="+90" swimtime="00:00:28.05" resultid="4323" lane="4" heatid="7349" entrytime="00:00:27.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="270" reactiontime="+91" swimtime="00:01:12.75" resultid="4319" lane="7" heatid="6842" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.15" />
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                    <SPLIT distance="75" swimtime="00:00:52.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-07-07" firstname="Jakub" gender="M" lastname="Gryczyński" nation="POL" athleteid="4324">
              <RESULTS>
                <RESULT eventid="1696" points="331" reactiontime="+85" swimtime="00:01:25.08" resultid="4328" heatid="7309" entrytime="00:01:22.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.87" />
                    <SPLIT distance="50" swimtime="00:00:38.79" />
                    <SPLIT distance="75" swimtime="00:01:01.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="285" reactiontime="+103" swimtime="00:03:13.61" resultid="4327" lane="8" heatid="7009" entrytime="00:03:09.61">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.94" />
                    <SPLIT distance="50" swimtime="00:00:41.78" />
                    <SPLIT distance="75" swimtime="00:01:05.70" />
                    <SPLIT distance="100" swimtime="00:01:29.90" />
                    <SPLIT distance="125" swimtime="00:01:55.18" />
                    <SPLIT distance="150" swimtime="00:02:21.10" />
                    <SPLIT distance="175" swimtime="00:02:48.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="358" reactiontime="+81" swimtime="00:00:38.25" resultid="4326" lane="6" heatid="6860" entrytime="00:00:38.19">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="271" reactiontime="+85" swimtime="00:01:19.03" resultid="4325" lane="3" heatid="6739" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.57" />
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                    <SPLIT distance="75" swimtime="00:00:57.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-06-06" firstname="Wojciech" gender="M" lastname="Zdzieszyński" nation="POL" athleteid="4329">
              <RESULTS>
                <RESULT eventid="1205" points="428" reactiontime="+90" swimtime="00:01:02.39" resultid="4331" heatid="6838" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.95" />
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                    <SPLIT distance="75" swimtime="00:00:45.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="361" reactiontime="+90" swimtime="00:01:11.79" resultid="4330" lane="4" heatid="6739" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.91" />
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                    <SPLIT distance="75" swimtime="00:00:54.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="323" reactiontime="+75" swimtime="00:00:35.63" resultid="4332" lane="1" heatid="7041" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="490" reactiontime="+86" swimtime="00:00:26.99" resultid="4334" lane="1" heatid="7348" entrytime="00:00:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="393" reactiontime="+89" swimtime="00:00:31.32" resultid="4333" heatid="7285" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-09-09" firstname="Witold" gender="M" lastname="Pietrowski" nation="POL" athleteid="4335">
              <RESULTS>
                <RESULT eventid="1645" points="393" reactiontime="+84" swimtime="00:00:31.34" resultid="4338" lane="8" heatid="7286" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="305" reactiontime="+78" swimtime="00:01:09.88" resultid="4336" lane="6" heatid="6837" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.72" />
                    <SPLIT distance="50" swimtime="00:00:31.15" />
                    <SPLIT distance="75" swimtime="00:00:49.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="4337" lane="8" heatid="7058" entrytime="00:02:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-08-08" firstname="Damian" gender="M" lastname="Karkusiński" nation="POL" athleteid="4339">
              <RESULTS>
                <RESULT eventid="1730" points="338" reactiontime="+61" swimtime="00:01:15.39" resultid="4343" lane="6" heatid="7325" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.99" />
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                    <SPLIT distance="75" swimtime="00:00:55.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="278" reactiontime="+65" swimtime="00:02:54.43" resultid="4341" lane="6" heatid="6886" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.68" />
                    <SPLIT distance="50" swimtime="00:00:36.92" />
                    <SPLIT distance="75" swimtime="00:00:57.42" />
                    <SPLIT distance="100" swimtime="00:01:19.08" />
                    <SPLIT distance="125" swimtime="00:01:41.97" />
                    <SPLIT distance="150" swimtime="00:02:05.74" />
                    <SPLIT distance="175" swimtime="00:02:30.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="348" reactiontime="+61" swimtime="00:00:34.76" resultid="4342" lane="2" heatid="7042" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="292" reactiontime="+92" swimtime="00:01:17.04" resultid="4340" heatid="6739" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.84" />
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                    <SPLIT distance="75" swimtime="00:00:57.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="385" reactiontime="+78" swimtime="00:00:29.23" resultid="4344" lane="1" heatid="7351" entrytime="00:00:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-09-09" firstname="Rafał" gender="M" lastname="Trudnos" nation="POL" athleteid="4345">
              <RESULTS>
                <RESULT eventid="1239" points="548" reactiontime="+75" swimtime="00:00:33.20" resultid="4347" lane="5" heatid="6866" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="442" reactiontime="+78" swimtime="00:02:47.33" resultid="4348" lane="1" heatid="7011" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.48" />
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                    <SPLIT distance="75" swimtime="00:00:56.64" />
                    <SPLIT distance="100" swimtime="00:01:17.84" />
                    <SPLIT distance="125" swimtime="00:01:39.55" />
                    <SPLIT distance="150" swimtime="00:02:01.45" />
                    <SPLIT distance="175" swimtime="00:02:24.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="490" reactiontime="+77" swimtime="00:01:14.72" resultid="4350" lane="1" heatid="7311" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.23" />
                    <SPLIT distance="50" swimtime="00:00:34.46" />
                    <SPLIT distance="75" swimtime="00:00:54.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="382" reactiontime="+78" swimtime="00:01:10.48" resultid="4346" lane="3" heatid="6741" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.53" />
                    <SPLIT distance="50" swimtime="00:00:32.42" />
                    <SPLIT distance="75" swimtime="00:00:53.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" status="DNS" swimtime="00:00:00.00" resultid="4349" lane="6" heatid="7079" entrytime="00:02:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-12" firstname="Igor" gender="M" lastname="Olejarczyk" nation="POL" athleteid="4351">
              <RESULTS>
                <RESULT eventid="1645" points="472" reactiontime="+78" swimtime="00:00:29.48" resultid="4354" lane="6" heatid="7288" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="401" reactiontime="+94" swimtime="00:01:03.76" resultid="4352" lane="8" heatid="6844" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.48" />
                    <SPLIT distance="50" swimtime="00:00:28.64" />
                    <SPLIT distance="75" swimtime="00:00:45.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="488" reactiontime="+80" swimtime="00:00:27.02" resultid="4355" lane="2" heatid="7351" entrytime="00:00:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" status="DNS" swimtime="00:00:00.00" resultid="4353" lane="2" heatid="7020" entrytime="00:01:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-03-03" firstname="Marcin" gender="M" lastname="Strąkowski" nation="POL" athleteid="4356">
              <RESULTS>
                <RESULT eventid="1239" points="349" reactiontime="+83" swimtime="00:00:38.60" resultid="4358" lane="2" heatid="6862" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="319" reactiontime="+85" swimtime="00:01:08.82" resultid="4357" lane="5" heatid="6838" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.83" />
                    <SPLIT distance="50" swimtime="00:00:32.16" />
                    <SPLIT distance="75" swimtime="00:00:50.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="401" reactiontime="+78" swimtime="00:00:28.85" resultid="4359" lane="7" heatid="7348" entrytime="00:00:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-04-04" firstname="Łukasz" gender="M" lastname="Raj" nation="POL" athleteid="4360">
              <RESULTS>
                <RESULT eventid="1239" points="321" reactiontime="+89" swimtime="00:00:39.67" resultid="4362" lane="2" heatid="6860" entrytime="00:00:38.19">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="245" reactiontime="+87" swimtime="00:01:21.66" resultid="4361" lane="2" heatid="6739" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.35" />
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                    <SPLIT distance="75" swimtime="00:01:00.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="333" reactiontime="+84" swimtime="00:00:30.69" resultid="4364" lane="6" heatid="7347" entrytime="00:00:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="4363" heatid="7062" entrytime="00:02:29.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-05-05" firstname="Kornel" gender="M" lastname="Pintara" nation="POL" athleteid="4365">
              <RESULTS>
                <RESULT eventid="1564" points="351" reactiontime="+87" swimtime="00:02:25.93" resultid="4366" lane="4" heatid="7063" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.31" />
                    <SPLIT distance="50" swimtime="00:00:30.47" />
                    <SPLIT distance="75" swimtime="00:00:47.01" />
                    <SPLIT distance="100" swimtime="00:01:04.28" />
                    <SPLIT distance="125" swimtime="00:01:22.55" />
                    <SPLIT distance="150" swimtime="00:01:42.88" />
                    <SPLIT distance="175" swimtime="00:02:04.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="411" reactiontime="+81" swimtime="00:00:30.86" resultid="4367" heatid="7290" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="456" reactiontime="+80" swimtime="00:00:27.63" resultid="4368" lane="8" heatid="7347" entrytime="00:00:28.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-03-03" firstname="Arkadiusz" gender="M" lastname="Olkowicz" nation="POL" athleteid="4369">
              <RESULTS>
                <RESULT eventid="1496" points="398" reactiontime="+81" swimtime="00:00:33.25" resultid="4373" lane="5" heatid="7042" entrytime="00:00:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="365" reactiontime="+84" swimtime="00:01:11.57" resultid="4370" lane="4" heatid="6741" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.69" />
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                    <SPLIT distance="75" swimtime="00:00:53.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="340" reactiontime="+78" swimtime="00:05:15.29" resultid="4372" lane="6" heatid="6909" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.98" />
                    <SPLIT distance="50" swimtime="00:00:31.92" />
                    <SPLIT distance="75" swimtime="00:00:49.75" />
                    <SPLIT distance="100" swimtime="00:01:07.95" />
                    <SPLIT distance="125" swimtime="00:01:27.00" />
                    <SPLIT distance="150" swimtime="00:01:46.41" />
                    <SPLIT distance="175" swimtime="00:02:06.68" />
                    <SPLIT distance="200" swimtime="00:02:27.22" />
                    <SPLIT distance="225" swimtime="00:02:47.99" />
                    <SPLIT distance="250" swimtime="00:03:08.86" />
                    <SPLIT distance="275" swimtime="00:03:29.63" />
                    <SPLIT distance="300" swimtime="00:03:51.13" />
                    <SPLIT distance="325" swimtime="00:04:12.49" />
                    <SPLIT distance="350" swimtime="00:04:33.63" />
                    <SPLIT distance="375" swimtime="00:04:54.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="445" reactiontime="+75" swimtime="00:00:27.86" resultid="4375" lane="6" heatid="7351" entrytime="00:00:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="4374" lane="6" heatid="7065" entrytime="00:02:10.00" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="4371" lane="2" heatid="6843" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-14" firstname="Tomasz" gender="M" lastname="Kotus" nation="POL" athleteid="4376">
              <RESULTS>
                <RESULT eventid="1798" points="400" reactiontime="+88" swimtime="00:05:30.91" resultid="4382" lane="8" heatid="7364" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.35" />
                    <SPLIT distance="50" swimtime="00:00:32.08" />
                    <SPLIT distance="75" swimtime="00:00:51.26" />
                    <SPLIT distance="100" swimtime="00:01:11.51" />
                    <SPLIT distance="125" swimtime="00:01:35.23" />
                    <SPLIT distance="150" swimtime="00:01:57.98" />
                    <SPLIT distance="175" swimtime="00:02:20.21" />
                    <SPLIT distance="200" swimtime="00:02:41.71" />
                    <SPLIT distance="225" swimtime="00:03:06.28" />
                    <SPLIT distance="250" swimtime="00:03:30.40" />
                    <SPLIT distance="275" swimtime="00:03:54.42" />
                    <SPLIT distance="300" swimtime="00:04:18.47" />
                    <SPLIT distance="325" swimtime="00:04:37.86" />
                    <SPLIT distance="350" swimtime="00:04:56.53" />
                    <SPLIT distance="375" swimtime="00:05:14.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="351" reactiontime="+88" swimtime="00:02:38.81" resultid="4378" heatid="6873" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.23" />
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                    <SPLIT distance="75" swimtime="00:00:51.62" />
                    <SPLIT distance="100" swimtime="00:01:12.66" />
                    <SPLIT distance="125" swimtime="00:01:33.43" />
                    <SPLIT distance="150" swimtime="00:01:55.30" />
                    <SPLIT distance="175" swimtime="00:02:16.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="396" swimtime="00:10:24.35" resultid="4377" heatid="6722" entrytime="00:10:45.00" />
                <RESULT eventid="1598" points="395" reactiontime="+88" swimtime="00:02:35.68" resultid="4380" lane="8" heatid="7076" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.67" />
                    <SPLIT distance="50" swimtime="00:00:30.04" />
                    <SPLIT distance="75" swimtime="00:00:51.49" />
                    <SPLIT distance="100" swimtime="00:01:12.22" />
                    <SPLIT distance="125" swimtime="00:01:36.63" />
                    <SPLIT distance="150" swimtime="00:02:00.47" />
                    <SPLIT distance="175" swimtime="00:02:18.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="431" reactiontime="+83" swimtime="00:01:06.70" resultid="4379" lane="2" heatid="7022" entrytime="00:01:06.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.59" />
                    <SPLIT distance="50" swimtime="00:00:30.08" />
                    <SPLIT distance="75" swimtime="00:00:47.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="4381" lane="5" heatid="7287" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-04-04" firstname="Joanna" gender="F" lastname="Wilińska Nowak" nation="POL" athleteid="4383">
              <RESULTS>
                <RESULT eventid="1479" points="416" reactiontime="+94" swimtime="00:00:37.04" resultid="4385" lane="1" heatid="7030" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="393" reactiontime="+91" swimtime="00:00:32.71" resultid="4386" heatid="7332" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="381" reactiontime="+94" swimtime="00:01:12.93" resultid="4384" lane="7" heatid="6827" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.48" />
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                    <SPLIT distance="75" swimtime="00:00:53.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-10-17" firstname="Ewa" gender="F" lastname="Kotus" nation="POL" athleteid="4387">
              <RESULTS>
                <RESULT eventid="1409" points="212" reactiontime="+102" swimtime="00:03:55.00" resultid="4391" lane="3" heatid="6999" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.50" />
                    <SPLIT distance="50" swimtime="00:00:52.66" />
                    <SPLIT distance="75" swimtime="00:01:21.95" />
                    <SPLIT distance="100" swimtime="00:01:51.78" />
                    <SPLIT distance="125" swimtime="00:02:22.30" />
                    <SPLIT distance="150" swimtime="00:02:53.04" />
                    <SPLIT distance="175" swimtime="00:03:24.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="193" reactiontime="+73" swimtime="00:03:36.59" resultid="4390" lane="4" heatid="6877" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.83" />
                    <SPLIT distance="50" swimtime="00:00:48.79" />
                    <SPLIT distance="75" swimtime="00:01:15.43" />
                    <SPLIT distance="100" swimtime="00:01:42.48" />
                    <SPLIT distance="125" swimtime="00:02:11.07" />
                    <SPLIT distance="150" swimtime="00:02:39.81" />
                    <SPLIT distance="175" swimtime="00:03:08.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="199" reactiontime="+81" swimtime="00:01:40.66" resultid="4393" lane="3" heatid="7315" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.92" />
                    <SPLIT distance="50" swimtime="00:00:49.46" />
                    <SPLIT distance="75" swimtime="00:01:15.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="171" reactiontime="+120" swimtime="00:01:57.24" resultid="4392" lane="7" heatid="7299" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.04" />
                    <SPLIT distance="50" swimtime="00:00:56.19" />
                    <SPLIT distance="75" swimtime="00:01:26.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="213" reactiontime="+91" swimtime="00:00:50.68" resultid="4389" lane="6" heatid="6850" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="210" reactiontime="+95" swimtime="00:01:38.91" resultid="4388" heatid="6724" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.02" />
                    <SPLIT distance="50" swimtime="00:00:46.08" />
                    <SPLIT distance="75" swimtime="00:01:14.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-05-03" firstname="Justyna" gender="F" lastname="Radzik" nation="POL" athleteid="4394">
              <RESULTS>
                <RESULT eventid="1679" points="188" reactiontime="+111" swimtime="00:01:53.58" resultid="4399" lane="1" heatid="7298" entrytime="00:01:45.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.59" />
                    <SPLIT distance="50" swimtime="00:00:55.46" />
                    <SPLIT distance="75" swimtime="00:01:24.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1409" points="194" reactiontime="+117" swimtime="00:04:01.82" resultid="4397" lane="6" heatid="6999" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.16" />
                    <SPLIT distance="50" swimtime="00:00:53.32" />
                    <SPLIT distance="75" swimtime="00:01:23.64" />
                    <SPLIT distance="100" swimtime="00:01:55.05" />
                    <SPLIT distance="125" swimtime="00:02:26.84" />
                    <SPLIT distance="150" swimtime="00:02:58.87" />
                    <SPLIT distance="175" swimtime="00:03:30.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="151" reactiontime="+109" swimtime="00:03:35.33" resultid="4398" lane="6" heatid="7050" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.48" />
                    <SPLIT distance="50" swimtime="00:00:46.89" />
                    <SPLIT distance="75" swimtime="00:01:13.71" />
                    <SPLIT distance="100" swimtime="00:01:41.95" />
                    <SPLIT distance="125" swimtime="00:02:11.15" />
                    <SPLIT distance="150" swimtime="00:02:40.12" />
                    <SPLIT distance="175" swimtime="00:03:09.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="188" reactiontime="+109" swimtime="00:00:52.90" resultid="4396" lane="4" heatid="6849" entrytime="00:00:52.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="143" reactiontime="+109" swimtime="00:01:52.44" resultid="4395" lane="7" heatid="6724" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.13" />
                    <SPLIT distance="50" swimtime="00:00:57.06" />
                    <SPLIT distance="75" swimtime="00:01:26.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" status="DNS" swimtime="00:00:00.00" resultid="4400" lane="6" heatid="7329" entrytime="00:00:49.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1177" points="447" reactiontime="+84" swimtime="00:01:53.45" resultid="4401" lane="1" heatid="6810" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.24" />
                    <SPLIT distance="50" swimtime="00:00:27.86" />
                    <SPLIT distance="75" swimtime="00:00:41.46" />
                    <SPLIT distance="100" swimtime="00:00:56.44" />
                    <SPLIT distance="125" swimtime="00:01:10.63" />
                    <SPLIT distance="150" swimtime="00:01:26.06" />
                    <SPLIT distance="175" swimtime="00:01:39.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" reactiontime="+84" />
                    <RELAYPOSITION number="2" reactiontime="+60" />
                    <RELAYPOSITION number="3" reactiontime="+81" />
                    <RELAYPOSITION number="4" reactiontime="+64" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1177" points="445" reactiontime="+78" swimtime="00:01:53.63" resultid="4402" heatid="6810" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.55" />
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                    <SPLIT distance="75" swimtime="00:00:42.80" />
                    <SPLIT distance="100" swimtime="00:00:58.62" />
                    <SPLIT distance="125" swimtime="00:01:11.67" />
                    <SPLIT distance="150" swimtime="00:01:25.91" />
                    <SPLIT distance="175" swimtime="00:01:39.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" reactiontime="+78" />
                    <RELAYPOSITION number="2" reactiontime="+58" />
                    <RELAYPOSITION number="3" reactiontime="+54" />
                    <RELAYPOSITION number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1177" points="469" reactiontime="+80" swimtime="00:01:51.62" resultid="4403" lane="5" heatid="6809" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.44" />
                    <SPLIT distance="50" swimtime="00:00:27.67" />
                    <SPLIT distance="75" swimtime="00:00:41.62" />
                    <SPLIT distance="100" swimtime="00:00:57.55" />
                    <SPLIT distance="125" swimtime="00:01:10.21" />
                    <SPLIT distance="150" swimtime="00:01:24.41" />
                    <SPLIT distance="175" swimtime="00:01:37.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" reactiontime="+80" />
                    <RELAYPOSITION number="2" reactiontime="+49" />
                    <RELAYPOSITION number="3" reactiontime="+32" />
                    <RELAYPOSITION number="4" reactiontime="+65" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1341" points="379" reactiontime="+70" swimtime="00:02:11.88" resultid="4404" heatid="6988" entrytime="00:02:04.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.06" />
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                    <SPLIT distance="75" swimtime="00:00:52.38" />
                    <SPLIT distance="100" swimtime="00:01:13.01" />
                    <SPLIT distance="125" swimtime="00:01:27.55" />
                    <SPLIT distance="150" swimtime="00:01:44.96" />
                    <SPLIT distance="175" swimtime="00:01:57.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4317" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="4345" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="4335" number="3" reactiontime="+71" />
                    <RELAYPOSITION athleteid="4329" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1341" points="448" reactiontime="+69" swimtime="00:02:04.73" resultid="4405" lane="8" heatid="6988" entrytime="00:02:04.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.10" />
                    <SPLIT distance="50" swimtime="00:00:34.30" />
                    <SPLIT distance="75" swimtime="00:00:49.26" />
                    <SPLIT distance="100" swimtime="00:01:07.56" />
                    <SPLIT distance="125" swimtime="00:01:21.21" />
                    <SPLIT distance="150" swimtime="00:01:37.65" />
                    <SPLIT distance="175" swimtime="00:01:50.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4339" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="4324" number="2" reactiontime="+38" />
                    <RELAYPOSITION athleteid="4351" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="4365" number="4" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="119" agemin="100" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1815" reactiontime="+69" swimtime="00:02:27.38" resultid="4407" lane="6" heatid="7503" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.24" />
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                    <SPLIT distance="75" swimtime="00:00:58.39" />
                    <SPLIT distance="100" swimtime="00:01:25.71" />
                    <SPLIT distance="125" swimtime="00:01:41.16" />
                    <SPLIT distance="150" swimtime="00:01:59.76" />
                    <SPLIT distance="175" swimtime="00:02:12.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4317" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="4394" number="2" reactiontime="+88" />
                    <RELAYPOSITION athleteid="4383" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="4376" number="4" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1615" reactiontime="+129" swimtime="00:02:17.41" resultid="4408" lane="3" heatid="7441" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.45" />
                    <SPLIT distance="50" swimtime="00:00:43.19" />
                    <SPLIT distance="75" swimtime="00:00:55.97" />
                    <SPLIT distance="100" swimtime="00:01:10.23" />
                    <SPLIT distance="125" swimtime="00:01:28.95" />
                    <SPLIT distance="150" swimtime="00:01:49.48" />
                    <SPLIT distance="175" swimtime="00:02:02.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4394" number="1" reactiontime="+129" />
                    <RELAYPOSITION athleteid="4356" number="2" reactiontime="+13" />
                    <RELAYPOSITION athleteid="4365" number="3" reactiontime="+69" />
                    <RELAYPOSITION athleteid="4387" number="4" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="TRLOD" name="MKS &quot;Trójka&quot; Łódź" nation="POL" region="LOD">
          <CONTACT city="Łódź" name="MKS &quot;Trójka&quot; Łódź" street="Sienkiewicza 46" zip="90-009" />
          <ATHLETES>
            <ATHLETE birthdate="1984-06-08" firstname="Marcin" gender="M" lastname="Babuchowski" nation="POL" athleteid="4411">
              <RESULTS>
                <RESULT comment="Rekord Polski " eventid="1564" points="737" reactiontime="+79" swimtime="00:01:53.94" resultid="4415" lane="4" heatid="7066" entrytime="00:01:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.88" />
                    <SPLIT distance="50" swimtime="00:00:25.85" />
                    <SPLIT distance="75" swimtime="00:00:40.45" />
                    <SPLIT distance="100" swimtime="00:00:55.37" />
                    <SPLIT distance="125" swimtime="00:01:10.38" />
                    <SPLIT distance="150" swimtime="00:01:25.34" />
                    <SPLIT distance="175" swimtime="00:01:40.26" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1645" points="802" reactiontime="+75" swimtime="00:00:24.71" resultid="4416" lane="4" heatid="7294" entrytime="00:00:23.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="734" reactiontime="+74" swimtime="00:00:23.59" resultid="4417" lane="3" heatid="7354" entrytime="00:00:23.97">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.45" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1273" points="758" reactiontime="+80" swimtime="00:02:02.86" resultid="4413" lane="4" heatid="6874" entrytime="00:02:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.61" />
                    <SPLIT distance="50" swimtime="00:00:26.54" />
                    <SPLIT distance="75" swimtime="00:00:41.64" />
                    <SPLIT distance="100" swimtime="00:00:57.34" />
                    <SPLIT distance="125" swimtime="00:01:13.59" />
                    <SPLIT distance="150" swimtime="00:01:30.10" />
                    <SPLIT distance="175" swimtime="00:01:46.81" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1109" points="668" swimtime="00:00:58.50" resultid="4412" lane="4" heatid="6745" entrytime="00:00:56.00" entrycourse="SCM" />
                <RESULT comment="Rekord Polski " eventid="1462" points="779" reactiontime="+77" swimtime="00:00:54.76" resultid="4414" lane="4" heatid="7023" entrytime="00:00:52.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.38" />
                    <SPLIT distance="50" swimtime="00:00:25.13" />
                    <SPLIT distance="75" swimtime="00:00:39.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="STWRO" name="Start Wrocław" nation="POL" region="DOL">
          <CONTACT city="Wrocław" email="wzsstart@post.pl" fax="071 34 372 81" internet="http://www.start.wroclaw.pl" name="Wojewódzkie Zrzeszenie Sportowe Niepełnosprawnych " phone="071 34 302 31" state="DOL" street="Notecka 12" zip="54-128" />
          <ATHLETES>
            <ATHLETE birthdate="1974-04-30" firstname="Sebastian" gender="M" lastname="Szymański" nation="POL" athleteid="4419">
              <RESULTS>
                <RESULT eventid="1764" points="453" reactiontime="+98" swimtime="00:00:27.70" resultid="4424" lane="6" heatid="7349" entrytime="00:00:27.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="442" reactiontime="+86" swimtime="00:00:30.14" resultid="4423" lane="1" heatid="7290" entrytime="00:00:30.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="364" reactiontime="+86" swimtime="00:00:34.26" resultid="4422" lane="2" heatid="7039" entrytime="00:00:34.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="433" reactiontime="+90" swimtime="00:01:02.17" resultid="4420" heatid="6841" entrytime="00:01:03.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.75" />
                    <SPLIT distance="50" swimtime="00:00:28.85" />
                    <SPLIT distance="75" swimtime="00:00:44.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" status="DNS" swimtime="00:00:00.00" resultid="4421" lane="3" heatid="7021" entrytime="00:01:08.90" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MABOL" name="Klub Pływacki Masters Bolesławiec" nation="POL" region="DOL">
          <CONTACT email="sekretarz-masters@o2.pl" name="Satoła Marta" />
          <ATHLETES>
            <ATHLETE birthdate="1948-11-29" firstname="Andrzej" gender="M" lastname="Daszyński" nation="POL" athleteid="4426">
              <RESULTS>
                <RESULT eventid="1462" points="78" reactiontime="+91" swimtime="00:01:57.84" resultid="4430" lane="7" heatid="7016" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.07" />
                    <SPLIT distance="50" swimtime="00:00:53.33" />
                    <SPLIT distance="75" swimtime="00:01:25.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="81" reactiontime="+91" swimtime="00:04:18.20" resultid="4428" heatid="6870" entrytime="00:04:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.03" />
                    <SPLIT distance="50" swimtime="00:00:56.07" />
                    <SPLIT distance="75" swimtime="00:01:28.62" />
                    <SPLIT distance="100" swimtime="00:02:02.40" />
                    <SPLIT distance="125" swimtime="00:02:37.10" />
                    <SPLIT distance="150" swimtime="00:03:12.20" />
                    <SPLIT distance="175" swimtime="00:03:45.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="116" reactiontime="+94" swimtime="00:03:53.89" resultid="4431" lane="3" heatid="7072" entrytime="00:03:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.63" />
                    <SPLIT distance="50" swimtime="00:00:53.91" />
                    <SPLIT distance="75" swimtime="00:01:24.02" />
                    <SPLIT distance="100" swimtime="00:01:51.89" />
                    <SPLIT distance="125" swimtime="00:02:28.73" />
                    <SPLIT distance="150" swimtime="00:03:03.77" />
                    <SPLIT distance="175" swimtime="00:03:31.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="123" reactiontime="+75" swimtime="00:03:48.61" resultid="4429" heatid="6882" entrytime="00:03:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.02" />
                    <SPLIT distance="50" swimtime="00:00:54.85" />
                    <SPLIT distance="75" swimtime="00:01:23.13" />
                    <SPLIT distance="100" swimtime="00:01:52.88" />
                    <SPLIT distance="125" swimtime="00:02:22.31" />
                    <SPLIT distance="150" swimtime="00:02:52.50" />
                    <SPLIT distance="175" swimtime="00:03:21.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="117" swimtime="00:15:35.69" resultid="4427" lane="6" heatid="6717" entrytime="00:15:00.00" />
                <RESULT eventid="1730" points="109" reactiontime="+78" swimtime="00:01:49.71" resultid="4432" lane="4" heatid="7319" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.35" />
                    <SPLIT distance="50" swimtime="00:00:53.96" />
                    <SPLIT distance="75" swimtime="00:01:22.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="114" reactiontime="+93" swimtime="00:08:22.27" resultid="4433" lane="4" heatid="7358" entrytime="00:08:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.02" />
                    <SPLIT distance="50" swimtime="00:00:57.22" />
                    <SPLIT distance="75" swimtime="00:01:32.23" />
                    <SPLIT distance="100" swimtime="00:02:07.58" />
                    <SPLIT distance="125" swimtime="00:02:39.55" />
                    <SPLIT distance="150" swimtime="00:03:10.30" />
                    <SPLIT distance="175" swimtime="00:03:40.63" />
                    <SPLIT distance="200" swimtime="00:04:10.90" />
                    <SPLIT distance="225" swimtime="00:04:46.47" />
                    <SPLIT distance="250" swimtime="00:05:21.35" />
                    <SPLIT distance="275" swimtime="00:05:56.25" />
                    <SPLIT distance="300" swimtime="00:06:32.53" />
                    <SPLIT distance="325" swimtime="00:07:01.41" />
                    <SPLIT distance="350" swimtime="00:07:31.21" />
                    <SPLIT distance="375" swimtime="00:07:58.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="BERLI" name="Berlin" nation="GER">
          <CONTACT name="D" />
          <ATHLETES>
            <ATHLETE birthdate="1967-01-01" firstname="Dariusz" gender="M" lastname="Domanski" nation="GER" athleteid="4483">
              <RESULTS>
                <RESULT eventid="1496" points="402" swimtime="00:00:33.13" resultid="4485" lane="5" heatid="7039" entrytime="00:00:34.50" />
                <RESULT eventid="1205" points="385" reactiontime="+105" swimtime="00:01:04.63" resultid="4484" lane="7" heatid="6841" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.90" />
                    <SPLIT distance="50" swimtime="00:00:31.55" />
                    <SPLIT distance="75" swimtime="00:00:48.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DELOD" name="Delfin Łódź" nation="POL">
          <CONTACT name="k" />
          <ATHLETES>
            <ATHLETE birthdate="1966-01-01" firstname="Piotr" gender="M" lastname="Kapczyński" nation="POL" athleteid="4487">
              <RESULTS>
                <RESULT eventid="1411" points="329" reactiontime="+87" swimtime="00:03:04.59" resultid="4489" lane="1" heatid="7008" entrytime="00:03:10.12">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.14" />
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                    <SPLIT distance="75" swimtime="00:01:04.14" />
                    <SPLIT distance="100" swimtime="00:01:27.48" />
                    <SPLIT distance="125" swimtime="00:01:51.64" />
                    <SPLIT distance="150" swimtime="00:02:16.24" />
                    <SPLIT distance="175" swimtime="00:02:40.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="396" reactiontime="+89" swimtime="00:00:36.99" resultid="4488" lane="1" heatid="6863" entrytime="00:00:36.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="DWTCZ" name="MSP Dwójka Tczew" nation="POL">
          <CONTACT name="g" />
          <ATHLETES>
            <ATHLETE birthdate="1986-01-01" firstname="Andrzej" gender="M" lastname="Gołembiewski" nation="POL" athleteid="4494">
              <RESULTS>
                <RESULT eventid="1075" points="309" swimtime="00:11:17.69" resultid="4495" lane="3" heatid="6721" entrytime="00:10:50.00" />
                <RESULT eventid="1375" points="355" reactiontime="+85" swimtime="00:05:10.60" resultid="4497" lane="8" heatid="6908" entrytime="00:05:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.99" />
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                    <SPLIT distance="75" swimtime="00:00:49.33" />
                    <SPLIT distance="100" swimtime="00:01:07.83" />
                    <SPLIT distance="125" swimtime="00:01:26.43" />
                    <SPLIT distance="150" swimtime="00:01:45.61" />
                    <SPLIT distance="175" swimtime="00:02:04.94" />
                    <SPLIT distance="200" swimtime="00:02:25.06" />
                    <SPLIT distance="225" swimtime="00:02:45.36" />
                    <SPLIT distance="250" swimtime="00:03:05.87" />
                    <SPLIT distance="275" swimtime="00:03:26.88" />
                    <SPLIT distance="300" swimtime="00:03:47.75" />
                    <SPLIT distance="325" swimtime="00:04:08.93" />
                    <SPLIT distance="350" swimtime="00:04:29.89" />
                    <SPLIT distance="375" swimtime="00:04:50.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="394" reactiontime="+91" swimtime="00:02:53.82" resultid="4498" heatid="7010" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.37" />
                    <SPLIT distance="50" swimtime="00:00:38.10" />
                    <SPLIT distance="75" swimtime="00:00:59.33" />
                    <SPLIT distance="100" swimtime="00:01:21.48" />
                    <SPLIT distance="125" swimtime="00:01:43.98" />
                    <SPLIT distance="150" swimtime="00:02:07.23" />
                    <SPLIT distance="175" swimtime="00:02:30.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="415" reactiontime="+79" swimtime="00:01:18.92" resultid="4500" lane="1" heatid="7310" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.49" />
                    <SPLIT distance="50" swimtime="00:00:36.17" />
                    <SPLIT distance="75" swimtime="00:00:57.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="494" reactiontime="+87" swimtime="00:00:34.37" resultid="4496" lane="7" heatid="6865" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="424" reactiontime="+85" swimtime="00:00:28.32" resultid="4501" lane="1" heatid="7347" entrytime="00:00:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="4499" lane="8" heatid="7064" entrytime="00:02:18.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PREGE" name="Pregel Kaliningrad" nation="RUS">
          <CONTACT name="Terwinski" />
          <ATHLETES>
            <ATHLETE birthdate="1957-01-01" firstname="Natalia" gender="F" lastname="Aleshchenko" nation="RUS" athleteid="4513">
              <RESULTS>
                <RESULT eventid="1058" points="323" swimtime="00:12:00.03" resultid="4514" lane="8" heatid="6715" entrytime="00:12:15.00" />
                <RESULT eventid="1445" points="277" reactiontime="+86" swimtime="00:01:26.81" resultid="4517" lane="8" heatid="7014" entrytime="00:01:26.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.40" />
                    <SPLIT distance="50" swimtime="00:00:39.91" />
                    <SPLIT distance="75" swimtime="00:01:02.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="346" reactiontime="+93" swimtime="00:05:44.03" resultid="4516" lane="8" heatid="6897" entrytime="00:05:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.42" />
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                    <SPLIT distance="75" swimtime="00:00:58.73" />
                    <SPLIT distance="100" swimtime="00:01:20.13" />
                    <SPLIT distance="125" swimtime="00:01:42.20" />
                    <SPLIT distance="150" swimtime="00:02:03.78" />
                    <SPLIT distance="175" swimtime="00:02:25.70" />
                    <SPLIT distance="200" swimtime="00:02:47.65" />
                    <SPLIT distance="225" swimtime="00:03:09.82" />
                    <SPLIT distance="250" swimtime="00:03:31.96" />
                    <SPLIT distance="275" swimtime="00:03:54.16" />
                    <SPLIT distance="300" swimtime="00:04:16.19" />
                    <SPLIT distance="325" swimtime="00:04:37.67" />
                    <SPLIT distance="350" swimtime="00:04:57.92" />
                    <SPLIT distance="375" swimtime="00:05:23.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="242" reactiontime="+92" swimtime="00:03:19.13" resultid="4515" lane="5" heatid="6868" entrytime="00:03:19.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.77" />
                    <SPLIT distance="50" swimtime="00:00:41.53" />
                    <SPLIT distance="75" swimtime="00:01:05.07" />
                    <SPLIT distance="100" swimtime="00:01:29.99" />
                    <SPLIT distance="125" swimtime="00:01:56.48" />
                    <SPLIT distance="150" swimtime="00:02:26.08" />
                    <SPLIT distance="175" swimtime="00:02:53.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1581" status="DNS" swimtime="00:00:00.00" resultid="4518" lane="7" heatid="7070" entrytime="00:03:12.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-01" firstname="Yuri" gender="M" lastname="Yakovenko" nation="RUS" athleteid="4519">
              <RESULTS>
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="4520" lane="2" heatid="6734" entrytime="00:01:29.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Akim" gender="M" lastname="Denisenko" nation="RUS" athleteid="4525">
              <RESULTS>
                <RESULT eventid="1239" points="207" reactiontime="+113" swimtime="00:00:45.91" resultid="4527" lane="7" heatid="6857" entrytime="00:00:43.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="142" reactiontime="+100" swimtime="00:01:37.95" resultid="4526" lane="6" heatid="6734" entrytime="00:01:29.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.62" />
                    <SPLIT distance="50" swimtime="00:00:45.05" />
                    <SPLIT distance="75" swimtime="00:01:15.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-01-01" firstname="Alexander" gender="M" lastname="Tervinskiy" nation="RUS" athleteid="4528">
              <RESULTS>
                <RESULT eventid="1239" points="348" reactiontime="+87" swimtime="00:00:38.61" resultid="4530" lane="1" heatid="6858" entrytime="00:00:41.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="233" reactiontime="+89" swimtime="00:01:23.10" resultid="4529" heatid="6735" entrytime="00:01:26.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.37" />
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                    <SPLIT distance="75" swimtime="00:01:02.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-01-01" firstname="Vadim" gender="M" lastname="Ezkov" nation="RUS" athleteid="4535">
              <RESULTS>
                <RESULT eventid="1696" points="360" reactiontime="+79" swimtime="00:01:22.76" resultid="4539" lane="4" heatid="7307" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.77" />
                    <SPLIT distance="50" swimtime="00:00:38.55" />
                    <SPLIT distance="75" swimtime="00:01:00.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="285" reactiontime="+78" swimtime="00:00:34.87" resultid="4538" lane="2" heatid="7286" entrytime="00:00:34.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="316" reactiontime="+75" swimtime="00:03:07.09" resultid="4537" lane="7" heatid="7009" entrytime="00:03:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.87" />
                    <SPLIT distance="50" swimtime="00:00:41.71" />
                    <SPLIT distance="75" swimtime="00:01:04.76" />
                    <SPLIT distance="100" swimtime="00:01:28.53" />
                    <SPLIT distance="125" swimtime="00:01:52.91" />
                    <SPLIT distance="150" swimtime="00:02:17.79" />
                    <SPLIT distance="175" swimtime="00:02:42.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="398" reactiontime="+77" swimtime="00:00:36.92" resultid="4536" lane="1" heatid="6860" entrytime="00:00:38.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Viktor" gender="M" lastname="Lyubavin" nation="RUS" athleteid="4540">
              <RESULTS>
                <RESULT eventid="1205" points="483" reactiontime="+76" swimtime="00:00:59.95" resultid="4542" lane="5" heatid="6842" entrytime="00:01:01.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.82" />
                    <SPLIT distance="50" swimtime="00:00:29.36" />
                    <SPLIT distance="75" swimtime="00:00:44.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="349" swimtime="00:20:41.87" resultid="4541" lane="6" heatid="6752" entrytime="00:20:59.00" />
                <RESULT eventid="1696" points="404" reactiontime="+79" swimtime="00:01:19.67" resultid="4544" lane="3" heatid="7309" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.17" />
                    <SPLIT distance="50" swimtime="00:00:37.75" />
                    <SPLIT distance="75" swimtime="00:00:58.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="477" reactiontime="+79" swimtime="00:00:27.23" resultid="4545" lane="6" heatid="7350" entrytime="00:00:27.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="398" reactiontime="+82" swimtime="00:02:19.90" resultid="4543" heatid="7064" entrytime="00:02:17.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.26" />
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                    <SPLIT distance="75" swimtime="00:00:50.32" />
                    <SPLIT distance="100" swimtime="00:01:08.44" />
                    <SPLIT distance="125" swimtime="00:01:26.69" />
                    <SPLIT distance="150" swimtime="00:01:45.11" />
                    <SPLIT distance="175" swimtime="00:02:03.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-01" firstname="Vladimir" gender="M" lastname="Chekutov" nation="RUS" athleteid="4546">
              <RESULTS>
                <RESULT eventid="1307" points="366" reactiontime="+84" swimtime="00:02:39.23" resultid="4549" lane="5" heatid="6886" entrytime="00:02:38.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.94" />
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                    <SPLIT distance="75" swimtime="00:00:56.08" />
                    <SPLIT distance="100" swimtime="00:01:16.27" />
                    <SPLIT distance="125" swimtime="00:01:36.43" />
                    <SPLIT distance="150" swimtime="00:01:57.29" />
                    <SPLIT distance="175" swimtime="00:02:18.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="347" reactiontime="+91" swimtime="00:01:12.76" resultid="4547" lane="3" heatid="6740" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.58" />
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                    <SPLIT distance="75" swimtime="00:00:55.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="447" reactiontime="+76" swimtime="00:01:01.51" resultid="4548" lane="6" heatid="6842" entrytime="00:01:01.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.71" />
                    <SPLIT distance="50" swimtime="00:00:29.11" />
                    <SPLIT distance="75" swimtime="00:00:45.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" status="DNS" swimtime="00:00:00.00" resultid="4550" lane="8" heatid="7041" entrytime="00:00:32.80" />
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="4552" lane="1" heatid="7349" entrytime="00:00:27.70" />
                <RESULT eventid="1730" status="DNS" swimtime="00:00:00.00" resultid="4551" lane="4" heatid="7324" entrytime="00:01:11.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-01" firstname="Yuri" gender="M" lastname="Ushakov" nation="RUS" athleteid="4553">
              <RESULTS>
                <RESULT eventid="1075" points="347" swimtime="00:10:52.12" resultid="4554" lane="6" heatid="6721" entrytime="00:11:05.00" />
                <RESULT eventid="1375" points="356" reactiontime="+95" swimtime="00:05:10.51" resultid="4556" lane="5" heatid="6907" entrytime="00:05:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.70" />
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                    <SPLIT distance="75" swimtime="00:00:51.28" />
                    <SPLIT distance="100" swimtime="00:01:10.01" />
                    <SPLIT distance="125" swimtime="00:01:29.43" />
                    <SPLIT distance="150" swimtime="00:01:48.75" />
                    <SPLIT distance="175" swimtime="00:02:08.68" />
                    <SPLIT distance="200" swimtime="00:02:28.85" />
                    <SPLIT distance="225" swimtime="00:02:49.08" />
                    <SPLIT distance="250" swimtime="00:03:09.63" />
                    <SPLIT distance="275" swimtime="00:03:29.73" />
                    <SPLIT distance="300" swimtime="00:03:50.40" />
                    <SPLIT distance="325" swimtime="00:04:11.07" />
                    <SPLIT distance="350" swimtime="00:04:31.52" />
                    <SPLIT distance="375" swimtime="00:04:51.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="363" reactiontime="+90" swimtime="00:02:24.24" resultid="4558" heatid="7063" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.33" />
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                    <SPLIT distance="75" swimtime="00:00:49.36" />
                    <SPLIT distance="100" swimtime="00:01:07.67" />
                    <SPLIT distance="125" swimtime="00:01:25.78" />
                    <SPLIT distance="150" swimtime="00:01:45.33" />
                    <SPLIT distance="175" swimtime="00:02:05.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="378" reactiontime="+89" swimtime="00:00:29.41" resultid="4560" lane="3" heatid="7346" entrytime="00:00:28.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="406" reactiontime="+103" swimtime="00:01:03.49" resultid="4555" lane="1" heatid="6841" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.94" />
                    <SPLIT distance="50" swimtime="00:00:31.03" />
                    <SPLIT distance="75" swimtime="00:00:47.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="314" reactiontime="+96" swimtime="00:00:33.76" resultid="4559" lane="1" heatid="7287" entrytime="00:00:33.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" status="DNS" swimtime="00:00:00.00" resultid="4557" lane="4" heatid="7020" entrytime="00:01:13.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-01" firstname="Sergey" gender="M" lastname="Bolgov" nation="RUS" athleteid="4561">
              <RESULTS>
                <RESULT eventid="1496" points="379" reactiontime="+72" swimtime="00:00:33.80" resultid="4564" lane="5" heatid="7038" entrytime="00:00:35.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="385" reactiontime="+93" swimtime="00:01:10.31" resultid="4562" lane="4" heatid="6742" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.48" />
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                    <SPLIT distance="75" swimtime="00:00:54.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="531" reactiontime="+76" swimtime="00:00:26.27" resultid="4566" lane="4" heatid="7351" entrytime="00:00:26.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="492" reactiontime="+96" swimtime="00:00:59.57" resultid="4563" lane="3" heatid="6843" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.68" />
                    <SPLIT distance="50" swimtime="00:00:28.83" />
                    <SPLIT distance="75" swimtime="00:00:44.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="401" reactiontime="+80" swimtime="00:00:31.13" resultid="4565" lane="8" heatid="7288" entrytime="00:00:32.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1177" status="DNS" swimtime="00:00:00.00" resultid="4567" lane="7" heatid="6809" entrytime="00:01:59.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4553" number="1" />
                    <RELAYPOSITION athleteid="4561" number="2" />
                    <RELAYPOSITION number="3" />
                    <RELAYPOSITION athleteid="4519" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1341" points="428" reactiontime="+77" swimtime="00:02:06.68" resultid="4568" lane="6" heatid="6987" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.39" />
                    <SPLIT distance="50" swimtime="00:00:32.88" />
                    <SPLIT distance="75" swimtime="00:00:49.05" />
                    <SPLIT distance="100" swimtime="00:01:08.24" />
                    <SPLIT distance="125" swimtime="00:01:23.40" />
                    <SPLIT distance="150" swimtime="00:01:40.93" />
                    <SPLIT distance="175" swimtime="00:01:53.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4546" number="1" reactiontime="+77" />
                    <RELAYPOSITION number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="4540" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="4561" number="4" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1177" points="373" reactiontime="+76" swimtime="00:02:00.45" resultid="4569" lane="4" heatid="6808" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.62" />
                    <SPLIT distance="50" swimtime="00:00:27.82" />
                    <SPLIT distance="75" swimtime="00:00:41.04" />
                    <SPLIT distance="100" swimtime="00:00:55.35" />
                    <SPLIT distance="125" swimtime="00:01:09.97" />
                    <SPLIT distance="150" swimtime="00:01:26.56" />
                    <SPLIT distance="175" swimtime="00:01:42.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4546" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="4540" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="4528" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="4525" number="4" reactiontime="+20" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1341" status="DNS" swimtime="00:00:00.00" resultid="4570" lane="1" heatid="6986" entrytime="00:02:29.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4553" number="1" />
                    <RELAYPOSITION athleteid="4528" number="2" />
                    <RELAYPOSITION athleteid="4525" number="3" />
                    <RELAYPOSITION athleteid="4519" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SKSLU" name="Skalar Słupsk" nation="POL">
          <CONTACT name="z" />
          <ATHLETES>
            <ATHLETE birthdate="1968-01-01" firstname="Beata" gender="F" lastname="Zubel" nation="POL" athleteid="4587">
              <RESULTS>
                <RESULT eventid="1713" points="414" reactiontime="+72" swimtime="00:01:18.81" resultid="4594" lane="7" heatid="7317" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.92" />
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                    <SPLIT distance="75" swimtime="00:00:59.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="462" reactiontime="+72" swimtime="00:00:35.77" resultid="4592" lane="8" heatid="7031" entrytime="00:00:36.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="419" reactiontime="+81" swimtime="00:00:40.50" resultid="4590" lane="8" heatid="6853" entrytime="00:00:40.29">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="451" reactiontime="+78" swimtime="00:01:08.93" resultid="4589" heatid="6828" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.49" />
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                    <SPLIT distance="75" swimtime="00:00:50.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="440" swimtime="00:01:17.26" resultid="4588" lane="2" heatid="6729" entrytime="00:01:16.75">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.95" />
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                    <SPLIT distance="75" swimtime="00:00:59.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" status="DNS" swimtime="00:00:00.00" resultid="4593" lane="1" heatid="7300" entrytime="00:01:29.80" />
                <RESULT eventid="1445" status="DNS" swimtime="00:00:00.00" resultid="4591" lane="5" heatid="7014" entrytime="00:01:15.60" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SPCZL" name="Starostwo Powiatowe Człuchów" nation="POL">
          <CONTACT name="t" />
          <ATHLETES>
            <ATHLETE birthdate="1986-01-01" firstname="Paweł" gender="M" lastname="Troka" nation="POL" athleteid="4596">
              <RESULTS>
                <RESULT eventid="1075" points="478" swimtime="00:09:46.53" resultid="4597" lane="1" heatid="6722" entrytime="00:10:00.41" />
                <RESULT eventid="1273" points="412" reactiontime="+84" swimtime="00:02:30.51" resultid="4599" lane="6" heatid="6874" entrytime="00:02:30.02">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.95" />
                    <SPLIT distance="50" swimtime="00:00:30.83" />
                    <SPLIT distance="75" swimtime="00:00:48.80" />
                    <SPLIT distance="100" swimtime="00:01:07.80" />
                    <SPLIT distance="125" swimtime="00:01:27.75" />
                    <SPLIT distance="150" swimtime="00:01:48.19" />
                    <SPLIT distance="175" swimtime="00:02:09.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="553" reactiontime="+82" swimtime="00:00:57.32" resultid="4598" lane="6" heatid="6844" entrytime="00:00:59.43">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.82" />
                    <SPLIT distance="50" swimtime="00:00:27.06" />
                    <SPLIT distance="75" swimtime="00:00:42.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="UMLOD" name="UM Łódź" nation="POL">
          <CONTACT name="b" />
        </CLUB>
        <CLUB type="CLUB" code="WIKRA" name="Wisła Kraków" nation="POL">
          <CONTACT name="Krokoszyński" />
          <ATHLETES>
            <ATHLETE birthdate="1930-01-01" firstname="Stanisław" gender="M" lastname="Krokoszyński" nation="POL" athleteid="4608">
              <RESULTS>
                <RESULT eventid="1109" points="118" reactiontime="+113" swimtime="00:01:44.11" resultid="4609" lane="1" heatid="6731" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.22" />
                    <SPLIT distance="50" swimtime="00:00:49.15" />
                    <SPLIT distance="75" swimtime="00:01:21.16" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1764" points="184" reactiontime="+115" swimtime="00:00:37.38" resultid="4613" lane="4" heatid="7337" entrytime="00:00:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="113" reactiontime="+121" swimtime="00:03:55.96" resultid="4612" lane="8" heatid="7073" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.69" />
                    <SPLIT distance="50" swimtime="00:00:54.54" />
                    <SPLIT distance="75" swimtime="00:01:23.71" />
                    <SPLIT distance="100" swimtime="00:01:53.45" />
                    <SPLIT distance="125" swimtime="00:02:28.36" />
                    <SPLIT distance="150" swimtime="00:03:03.20" />
                    <SPLIT distance="175" swimtime="00:03:29.73" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1375" points="133" swimtime="00:07:10.86" resultid="4611" heatid="6900" entrytime="00:07:30.00" />
                <RESULT comment="Rekord Polski " eventid="1205" points="155" reactiontime="+110" swimtime="00:01:27.46" resultid="4610" lane="8" heatid="6832" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.25" />
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                    <SPLIT distance="75" swimtime="00:01:03.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Janusz" gender="M" lastname="Konstanty" nation="POL" athleteid="4615">
              <RESULTS>
                <RESULT eventid="1598" points="264" reactiontime="+86" swimtime="00:02:58.06" resultid="4619" lane="1" heatid="7076" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.27" />
                    <SPLIT distance="50" swimtime="00:00:36.88" />
                    <SPLIT distance="75" swimtime="00:00:59.86" />
                    <SPLIT distance="100" swimtime="00:01:22.25" />
                    <SPLIT distance="125" swimtime="00:01:48.65" />
                    <SPLIT distance="150" swimtime="00:02:16.87" />
                    <SPLIT distance="175" swimtime="00:02:38.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="260" reactiontime="+92" swimtime="00:01:20.12" resultid="4616" lane="8" heatid="6737" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.14" />
                    <SPLIT distance="50" swimtime="00:00:37.20" />
                    <SPLIT distance="75" swimtime="00:01:00.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="302" reactiontime="+74" swimtime="00:01:18.27" resultid="4620" lane="4" heatid="7322" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.53" />
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                    <SPLIT distance="75" swimtime="00:00:57.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="315" reactiontime="+78" swimtime="00:00:35.94" resultid="4618" lane="2" heatid="7037" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="289" reactiontime="+80" swimtime="00:02:52.31" resultid="4617" lane="5" heatid="6884" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.13" />
                    <SPLIT distance="50" swimtime="00:00:38.42" />
                    <SPLIT distance="75" swimtime="00:00:59.05" />
                    <SPLIT distance="100" swimtime="00:01:21.14" />
                    <SPLIT distance="150" swimtime="00:02:07.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WKPOZ" name="WKB Poznań" nation="POL">
          <CONTACT name="z" />
          <ATHLETES>
            <ATHLETE birthdate="1946-01-01" firstname="Teresa" gender="F" lastname="Zarzeczańska-Różańska" nation="POL" athleteid="4622">
              <RESULTS>
                <RESULT eventid="1126" status="DNS" swimtime="00:00:00.00" resultid="4623" lane="2" heatid="6746" entrytime="00:37:00.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WOPAB" name="WOPR Pabianice" nation="POL">
          <CONTACT name="w" />
          <ATHLETES>
            <ATHLETE birthdate="1967-01-01" firstname="Jarosław" gender="M" lastname="Wyrwa" nation="POL" athleteid="4625">
              <RESULTS>
                <RESULT eventid="1239" points="372" reactiontime="+80" swimtime="00:00:37.79" resultid="4626" heatid="6860" entrytime="00:00:39.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="274" reactiontime="+79" swimtime="00:03:16.28" resultid="4627" lane="7" heatid="7007" entrytime="00:03:25.02">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.41" />
                    <SPLIT distance="50" swimtime="00:00:43.59" />
                    <SPLIT distance="75" swimtime="00:01:07.42" />
                    <SPLIT distance="100" swimtime="00:01:31.94" />
                    <SPLIT distance="125" swimtime="00:01:58.40" />
                    <SPLIT distance="150" swimtime="00:02:24.16" />
                    <SPLIT distance="175" swimtime="00:02:50.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ALMOS" name="All Stars Moscow" nation="RUS">
          <CONTACT name="l" />
          <ATHLETES>
            <ATHLETE birthdate="1955-01-01" firstname="Ludmila" gender="F" lastname="Lukashova" nation="RUS" athleteid="4635">
              <RESULTS>
                <RESULT eventid="1713" points="126" reactiontime="+86" swimtime="00:01:57.07" resultid="4639" lane="7" heatid="7314" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.76" />
                    <SPLIT distance="50" swimtime="00:00:56.19" />
                    <SPLIT distance="75" swimtime="00:01:27.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="114" reactiontime="+80" swimtime="00:04:18.15" resultid="4637" lane="3" heatid="6876" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.00" />
                    <SPLIT distance="50" swimtime="00:00:58.47" />
                    <SPLIT distance="75" swimtime="00:01:30.10" />
                    <SPLIT distance="100" swimtime="00:02:03.41" />
                    <SPLIT distance="125" swimtime="00:02:37.49" />
                    <SPLIT distance="150" swimtime="00:03:12.83" />
                    <SPLIT distance="175" swimtime="00:03:46.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="150" reactiontime="+86" swimtime="00:00:52.02" resultid="4638" lane="6" heatid="7026" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="124" reactiontime="+113" swimtime="00:01:57.89" resultid="4636" lane="6" heatid="6724" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.70" />
                    <SPLIT distance="50" swimtime="00:00:56.40" />
                    <SPLIT distance="75" swimtime="00:01:30.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="GDANS" name="Gdańsk" nation="POL">
          <CONTACT name="n" />
          <ATHLETES>
            <ATHLETE birthdate="1977-01-01" firstname="Adam" gender="M" lastname="Nadolski" nation="POL" athleteid="4641">
              <RESULTS>
                <RESULT eventid="1411" points="410" reactiontime="+87" swimtime="00:02:51.57" resultid="4644" lane="1" heatid="7010" entrytime="00:02:57.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.70" />
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                    <SPLIT distance="75" swimtime="00:00:58.34" />
                    <SPLIT distance="100" swimtime="00:01:20.63" />
                    <SPLIT distance="125" swimtime="00:01:42.96" />
                    <SPLIT distance="150" swimtime="00:02:05.87" />
                    <SPLIT distance="175" swimtime="00:02:29.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="530" reactiontime="+85" swimtime="00:00:33.57" resultid="4642" lane="1" heatid="6865" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="422" reactiontime="+88" swimtime="00:01:18.53" resultid="4646" lane="2" heatid="7310" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.37" />
                    <SPLIT distance="50" swimtime="00:00:35.83" />
                    <SPLIT distance="75" swimtime="00:00:56.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="327" reactiontime="+90" swimtime="00:05:19.33" resultid="4643" lane="4" heatid="6906" entrytime="00:05:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.26" />
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="75" swimtime="00:00:54.17" />
                    <SPLIT distance="100" swimtime="00:01:13.91" />
                    <SPLIT distance="125" swimtime="00:01:33.62" />
                    <SPLIT distance="150" swimtime="00:01:54.11" />
                    <SPLIT distance="175" swimtime="00:02:14.25" />
                    <SPLIT distance="200" swimtime="00:02:34.66" />
                    <SPLIT distance="225" swimtime="00:02:54.70" />
                    <SPLIT distance="250" swimtime="00:03:15.43" />
                    <SPLIT distance="275" swimtime="00:03:36.13" />
                    <SPLIT distance="300" swimtime="00:03:56.92" />
                    <SPLIT distance="325" swimtime="00:04:17.41" />
                    <SPLIT distance="350" swimtime="00:04:38.47" />
                    <SPLIT distance="375" swimtime="00:04:58.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="434" reactiontime="+85" swimtime="00:00:28.09" resultid="4647" lane="4" heatid="7350" entrytime="00:00:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.57" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Z 2" eventid="1598" reactiontime="+82" status="DSQ" swimtime="00:00:00.00" resultid="4645" lane="6" heatid="7078" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.40" />
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                    <SPLIT distance="75" swimtime="00:00:53.77" />
                    <SPLIT distance="100" swimtime="00:01:15.73" />
                    <SPLIT distance="125" swimtime="00:01:38.05" />
                    <SPLIT distance="150" swimtime="00:02:00.99" />
                    <SPLIT distance="175" swimtime="00:02:22.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="GDYNI" name="Gdynia" nation="POL">
          <CONTACT name="g" />
          <ATHLETES>
            <ATHLETE birthdate="1948-01-02" firstname="Janusz" gender="M" lastname="Płonka" nation="POL" athleteid="3375">
              <RESULTS>
                <RESULT eventid="1462" points="67" reactiontime="+87" swimtime="00:02:03.68" resultid="3379" lane="3" heatid="7015" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.90" />
                    <SPLIT distance="50" swimtime="00:00:58.62" />
                    <SPLIT distance="75" swimtime="00:01:31.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="66" reactiontime="+89" swimtime="00:04:36.22" resultid="3377" lane="2" heatid="6869" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.06" />
                    <SPLIT distance="50" swimtime="00:01:01.50" />
                    <SPLIT distance="75" swimtime="00:01:38.82" />
                    <SPLIT distance="100" swimtime="00:02:16.26" />
                    <SPLIT distance="125" swimtime="00:02:53.10" />
                    <SPLIT distance="150" swimtime="00:03:31.33" />
                    <SPLIT distance="175" swimtime="00:04:04.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="58" reactiontime="+85" swimtime="00:04:54.22" resultid="3378" heatid="6881" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.63" />
                    <SPLIT distance="50" swimtime="00:01:12.74" />
                    <SPLIT distance="75" swimtime="00:03:11.60" />
                    <SPLIT distance="100" swimtime="00:02:31.58" />
                    <SPLIT distance="125" swimtime="00:04:23.27" />
                    <SPLIT distance="150" swimtime="00:03:48.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="69" reactiontime="+85" swimtime="00:04:37.86" resultid="3380" lane="8" heatid="7072" entrytime="00:04:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.49" />
                    <SPLIT distance="50" swimtime="00:01:01.68" />
                    <SPLIT distance="75" swimtime="00:01:43.04" />
                    <SPLIT distance="100" swimtime="00:02:23.94" />
                    <SPLIT distance="125" swimtime="00:02:59.30" />
                    <SPLIT distance="150" swimtime="00:03:35.26" />
                    <SPLIT distance="175" swimtime="00:04:09.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="87" reactiontime="+83" swimtime="00:00:51.74" resultid="3381" lane="6" heatid="7281" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="70" reactiontime="+94" swimtime="00:02:03.97" resultid="3376" lane="4" heatid="6730" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.67" />
                    <SPLIT distance="50" swimtime="00:01:03.57" />
                    <SPLIT distance="75" swimtime="00:01:36.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="64" reactiontime="+91" swimtime="00:10:07.57" resultid="3382" lane="1" heatid="7358" entrytime="00:10:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.10" />
                    <SPLIT distance="50" swimtime="00:01:06.16" />
                    <SPLIT distance="75" swimtime="00:01:44.12" />
                    <SPLIT distance="100" swimtime="00:02:22.70" />
                    <SPLIT distance="125" swimtime="00:03:08.98" />
                    <SPLIT distance="150" swimtime="00:03:52.31" />
                    <SPLIT distance="175" swimtime="00:04:35.32" />
                    <SPLIT distance="200" swimtime="00:05:19.21" />
                    <SPLIT distance="225" swimtime="00:05:57.55" />
                    <SPLIT distance="250" swimtime="00:06:36.82" />
                    <SPLIT distance="275" swimtime="00:07:13.12" />
                    <SPLIT distance="300" swimtime="00:07:49.62" />
                    <SPLIT distance="325" swimtime="00:08:27.74" />
                    <SPLIT distance="350" swimtime="00:09:04.20" />
                    <SPLIT distance="375" swimtime="00:09:38.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-01-01" firstname="Beata" gender="F" lastname="Galska" nation="POL" athleteid="4649">
              <RESULTS>
                <RESULT eventid="1679" status="DNS" swimtime="00:00:00.00" resultid="4654" lane="6" heatid="7298" entrytime="00:01:45.43" />
                <RESULT eventid="1222" status="DNS" swimtime="00:00:00.00" resultid="4651" lane="1" heatid="6851" entrytime="00:00:45.43" />
                <RESULT eventid="1409" status="DNS" swimtime="00:00:00.00" resultid="4652" lane="8" heatid="7000" entrytime="00:03:34.01" />
                <RESULT eventid="1547" status="DNS" swimtime="00:00:00.00" resultid="4653" lane="6" heatid="7051" entrytime="00:02:59.07" />
                <RESULT eventid="1747" status="DNS" swimtime="00:00:00.00" resultid="4655" lane="5" heatid="7331" entrytime="00:00:36.41" />
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="4650" lane="3" heatid="6825" entrytime="00:01:20.06" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KORCZ" name="Korczyna" nation="POL">
          <CONTACT name="Ż" />
          <ATHLETES>
            <ATHLETE birthdate="1966-01-01" firstname="Bogdan" gender="M" lastname="Żebracki" nation="POL" athleteid="4657">
              <RESULTS>
                <RESULT eventid="1730" points="269" reactiontime="+97" swimtime="00:01:21.36" resultid="4664" lane="5" heatid="7323" entrytime="00:01:18.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.48" />
                    <SPLIT distance="50" swimtime="00:00:39.02" />
                    <SPLIT distance="75" swimtime="00:01:00.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="317" reactiontime="+98" swimtime="00:03:06.88" resultid="4661" lane="1" heatid="7009" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.15" />
                    <SPLIT distance="50" swimtime="00:00:40.75" />
                    <SPLIT distance="75" swimtime="00:01:04.42" />
                    <SPLIT distance="100" swimtime="00:01:28.51" />
                    <SPLIT distance="125" swimtime="00:01:53.07" />
                    <SPLIT distance="150" swimtime="00:02:18.36" />
                    <SPLIT distance="175" swimtime="00:02:43.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="349" reactiontime="+84" swimtime="00:01:23.63" resultid="4663" lane="8" heatid="7309" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.81" />
                    <SPLIT distance="50" swimtime="00:00:38.65" />
                    <SPLIT distance="75" swimtime="00:01:00.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="275" reactiontime="+102" swimtime="00:02:55.11" resultid="4660" heatid="6885" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.07" />
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                    <SPLIT distance="75" swimtime="00:01:01.56" />
                    <SPLIT distance="100" swimtime="00:01:24.34" />
                    <SPLIT distance="125" swimtime="00:01:47.53" />
                    <SPLIT distance="150" swimtime="00:02:11.19" />
                    <SPLIT distance="175" swimtime="00:02:34.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="323" reactiontime="+97" swimtime="00:00:35.65" resultid="4662" lane="2" heatid="7038" entrytime="00:00:35.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="301" reactiontime="+93" swimtime="00:01:16.32" resultid="4658" lane="5" heatid="6738" entrytime="00:01:15.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.87" />
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                    <SPLIT distance="75" swimtime="00:00:58.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="394" reactiontime="+88" swimtime="00:00:37.06" resultid="4659" lane="7" heatid="6862" entrytime="00:00:37.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KORNI" name="Kórnik" nation="POL">
          <CONTACT name="t" />
          <ATHLETES>
            <ATHLETE birthdate="1972-01-01" firstname="Dominik" gender="M" lastname="Tomaszewski" nation="POL" athleteid="4666">
              <RESULTS>
                <RESULT eventid="1798" points="204" reactiontime="+107" swimtime="00:06:53.84" resultid="4673" lane="2" heatid="7360" entrytime="00:07:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.46" />
                    <SPLIT distance="50" swimtime="00:00:45.34" />
                    <SPLIT distance="75" swimtime="00:01:11.04" />
                    <SPLIT distance="100" swimtime="00:01:39.10" />
                    <SPLIT distance="125" swimtime="00:02:08.88" />
                    <SPLIT distance="150" swimtime="00:02:36.71" />
                    <SPLIT distance="175" swimtime="00:03:07.25" />
                    <SPLIT distance="200" swimtime="00:03:36.73" />
                    <SPLIT distance="225" swimtime="00:04:03.56" />
                    <SPLIT distance="250" swimtime="00:04:30.25" />
                    <SPLIT distance="275" swimtime="00:04:57.61" />
                    <SPLIT distance="300" swimtime="00:05:24.50" />
                    <SPLIT distance="325" swimtime="00:05:47.30" />
                    <SPLIT distance="350" swimtime="00:06:10.06" />
                    <SPLIT distance="375" swimtime="00:06:33.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="221" swimtime="00:12:38.22" resultid="4667" lane="3" heatid="6718" entrytime="00:12:45.00" />
                <RESULT eventid="1375" points="216" reactiontime="+109" swimtime="00:06:06.69" resultid="4669" lane="5" heatid="6902" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.79" />
                    <SPLIT distance="50" swimtime="00:00:40.28" />
                    <SPLIT distance="75" swimtime="00:01:01.29" />
                    <SPLIT distance="100" swimtime="00:01:24.01" />
                    <SPLIT distance="125" swimtime="00:01:46.88" />
                    <SPLIT distance="150" swimtime="00:02:10.70" />
                    <SPLIT distance="175" swimtime="00:02:34.34" />
                    <SPLIT distance="200" swimtime="00:02:58.32" />
                    <SPLIT distance="225" swimtime="00:03:22.16" />
                    <SPLIT distance="250" swimtime="00:03:46.46" />
                    <SPLIT distance="275" swimtime="00:04:10.48" />
                    <SPLIT distance="300" swimtime="00:04:35.22" />
                    <SPLIT distance="325" swimtime="00:04:58.96" />
                    <SPLIT distance="350" swimtime="00:05:23.11" />
                    <SPLIT distance="375" swimtime="00:05:45.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="152" reactiontime="+111" swimtime="00:01:34.35" resultid="4670" lane="5" heatid="7017" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.14" />
                    <SPLIT distance="50" swimtime="00:00:40.90" />
                    <SPLIT distance="75" swimtime="00:01:06.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="195" reactiontime="+108" swimtime="00:00:39.53" resultid="4672" lane="4" heatid="7283" entrytime="00:00:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="4668" lane="2" heatid="6833" entrytime="00:01:20.00" />
                <RESULT eventid="1598" status="DNS" swimtime="00:00:00.00" resultid="4671" lane="6" heatid="7074" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.55" />
                    <SPLIT distance="50" swimtime="00:00:42.20" />
                    <SPLIT distance="75" swimtime="00:01:10.06" />
                    <SPLIT distance="100" swimtime="00:01:39.71" />
                    <SPLIT distance="125" swimtime="00:02:09.89" />
                    <SPLIT distance="150" swimtime="00:02:40.21" />
                    <SPLIT distance="175" swimtime="00:03:03.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-01-01" firstname="Krzysztof" gender="M" lastname="Buszkiewicz" nation="POL" athleteid="6666">
              <RESULTS>
                <RESULT eventid="1764" points="430" reactiontime="+91" swimtime="00:00:28.18" resultid="7495" lane="2" heatid="7347">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="KRAKO" name="Kraków" nation="POL">
          <CONTACT name="g" />
          <ATHLETES>
            <ATHLETE birthdate="1958-01-01" firstname="Jadwiga" gender="F" lastname="Górecka-Burkot" nation="POL" athleteid="4675">
              <RESULTS>
                <RESULT eventid="1747" points="333" reactiontime="+75" swimtime="00:00:34.58" resultid="4681" heatid="7333" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="259" reactiontime="+74" swimtime="00:01:22.92" resultid="4677" lane="4" heatid="6825" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.20" />
                    <SPLIT distance="50" swimtime="00:00:39.53" />
                    <SPLIT distance="75" swimtime="00:01:02.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="245" reactiontime="+76" swimtime="00:00:40.66" resultid="4680" lane="2" heatid="7277" entrytime="00:00:44.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.80" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Z 1" eventid="1092" status="DSQ" swimtime="00:00:00.00" resultid="4676" lane="2" heatid="6725" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.33" />
                    <SPLIT distance="50" swimtime="00:00:49.80" />
                    <SPLIT distance="75" swimtime="00:01:18.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="4678" lane="6" heatid="7028" entrytime="00:00:43.00" />
                <RESULT eventid="1547" status="DNS" swimtime="00:00:00.00" resultid="4679" heatid="7051" entrytime="00:03:08.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MAGRY" name="Marlin Gryfino" nation="POL">
          <CONTACT name="g" />
          <ATHLETES>
            <ATHLETE birthdate="1953-01-01" firstname="Sławomir" gender="M" lastname="Grzeszewski" nation="POL" athleteid="4683">
              <RESULTS>
                <RESULT eventid="1411" points="279" reactiontime="+90" swimtime="00:03:15.12" resultid="4686" lane="1" heatid="7007" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.80" />
                    <SPLIT distance="50" swimtime="00:00:43.11" />
                    <SPLIT distance="75" swimtime="00:01:07.67" />
                    <SPLIT distance="100" swimtime="00:01:32.54" />
                    <SPLIT distance="125" swimtime="00:01:58.33" />
                    <SPLIT distance="150" swimtime="00:02:23.82" />
                    <SPLIT distance="175" swimtime="00:02:50.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="304" reactiontime="+83" swimtime="00:01:27.60" resultid="4687" lane="2" heatid="7307" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.43" />
                    <SPLIT distance="50" swimtime="00:00:39.69" />
                    <SPLIT distance="75" swimtime="00:01:02.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="328" reactiontime="+82" swimtime="00:00:39.38" resultid="4685" lane="6" heatid="6859" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="231" reactiontime="+81" swimtime="00:01:23.28" resultid="4684" lane="4" heatid="6735" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.61" />
                    <SPLIT distance="50" swimtime="00:00:39.86" />
                    <SPLIT distance="75" swimtime="00:01:03.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ORRAD" name="Orka Radlin" nation="POL">
          <CONTACT name="b" />
          <ATHLETES>
            <ATHLETE birthdate="1940-01-01" firstname="Rudolf" gender="M" lastname="Bugla" nation="POL" athleteid="4689">
              <RESULTS>
                <RESULT eventid="1798" points="96" reactiontime="+99" swimtime="00:08:51.98" resultid="4696" lane="7" heatid="7358" entrytime="00:08:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.11" />
                    <SPLIT distance="50" swimtime="00:00:56.78" />
                    <SPLIT distance="75" swimtime="00:01:29.02" />
                    <SPLIT distance="100" swimtime="00:02:02.69" />
                    <SPLIT distance="125" swimtime="00:02:36.22" />
                    <SPLIT distance="150" swimtime="00:03:10.65" />
                    <SPLIT distance="175" swimtime="00:03:46.44" />
                    <SPLIT distance="200" swimtime="00:04:22.58" />
                    <SPLIT distance="225" swimtime="00:04:57.96" />
                    <SPLIT distance="250" swimtime="00:05:31.74" />
                    <SPLIT distance="275" swimtime="00:06:06.89" />
                    <SPLIT distance="300" swimtime="00:06:42.85" />
                    <SPLIT distance="325" swimtime="00:07:14.58" />
                    <SPLIT distance="350" swimtime="00:07:46.87" />
                    <SPLIT distance="375" swimtime="00:08:20.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="88" reactiontime="+95" swimtime="00:04:11.86" resultid="4691" lane="7" heatid="6870" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.12" />
                    <SPLIT distance="50" swimtime="00:00:55.89" />
                    <SPLIT distance="75" swimtime="00:01:26.97" />
                    <SPLIT distance="100" swimtime="00:01:58.51" />
                    <SPLIT distance="125" swimtime="00:02:31.33" />
                    <SPLIT distance="150" swimtime="00:03:03.80" />
                    <SPLIT distance="175" swimtime="00:03:38.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="77" reactiontime="+93" swimtime="00:01:57.96" resultid="4693" lane="6" heatid="7016" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.80" />
                    <SPLIT distance="50" swimtime="00:00:52.69" />
                    <SPLIT distance="75" swimtime="00:01:24.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="96" reactiontime="+99" swimtime="00:04:09.40" resultid="4694" lane="6" heatid="7072" entrytime="00:04:04.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.81" />
                    <SPLIT distance="50" swimtime="00:00:55.13" />
                    <SPLIT distance="75" swimtime="00:01:26.47" />
                    <SPLIT distance="100" swimtime="00:01:58.87" />
                    <SPLIT distance="125" swimtime="00:02:33.03" />
                    <SPLIT distance="150" swimtime="00:03:06.69" />
                    <SPLIT distance="175" swimtime="00:03:36.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="83" reactiontime="+81" swimtime="00:02:00.33" resultid="4695" lane="5" heatid="7319" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.67" />
                    <SPLIT distance="50" swimtime="00:00:57.33" />
                    <SPLIT distance="75" swimtime="00:01:28.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="109" reactiontime="+101" swimtime="00:01:46.89" resultid="4690" lane="3" heatid="6731" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.40" />
                    <SPLIT distance="50" swimtime="00:00:52.23" />
                    <SPLIT distance="75" swimtime="00:01:21.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="74" reactiontime="+84" swimtime="00:04:30.54" resultid="4692" lane="3" heatid="6881" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.72" />
                    <SPLIT distance="50" swimtime="00:01:02.16" />
                    <SPLIT distance="75" swimtime="00:01:37.79" />
                    <SPLIT distance="100" swimtime="00:02:12.20" />
                    <SPLIT distance="125" swimtime="00:02:46.42" />
                    <SPLIT distance="150" swimtime="00:03:21.23" />
                    <SPLIT distance="175" swimtime="00:03:56.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Leon" gender="M" lastname="Irczyk" nation="POL" athleteid="4697">
              <RESULTS>
                <RESULT eventid="1564" points="114" reactiontime="+107" swimtime="00:03:31.74" resultid="4702" lane="1" heatid="7055" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.81" />
                    <SPLIT distance="50" swimtime="00:00:46.31" />
                    <SPLIT distance="75" swimtime="00:01:12.54" />
                    <SPLIT distance="100" swimtime="00:01:40.56" />
                    <SPLIT distance="125" swimtime="00:02:08.88" />
                    <SPLIT distance="150" swimtime="00:02:36.77" />
                    <SPLIT distance="175" swimtime="00:03:04.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="115" reactiontime="+138" swimtime="00:08:21.21" resultid="4704" lane="6" heatid="7358" entrytime="00:09:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.37" />
                    <SPLIT distance="50" swimtime="00:00:58.38" />
                    <SPLIT distance="75" swimtime="00:01:32.06" />
                    <SPLIT distance="100" swimtime="00:02:04.52" />
                    <SPLIT distance="125" swimtime="00:02:42.56" />
                    <SPLIT distance="150" swimtime="00:03:20.06" />
                    <SPLIT distance="175" swimtime="00:03:57.18" />
                    <SPLIT distance="200" swimtime="00:04:33.75" />
                    <SPLIT distance="225" swimtime="00:05:04.42" />
                    <SPLIT distance="250" swimtime="00:05:33.06" />
                    <SPLIT distance="275" swimtime="00:06:02.42" />
                    <SPLIT distance="300" swimtime="00:06:31.84" />
                    <SPLIT distance="325" swimtime="00:06:59.51" />
                    <SPLIT distance="350" swimtime="00:07:26.81" />
                    <SPLIT distance="375" swimtime="00:07:54.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="174" reactiontime="+108" swimtime="00:01:45.41" resultid="4703" lane="2" heatid="7304" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.85" />
                    <SPLIT distance="50" swimtime="00:00:51.59" />
                    <SPLIT distance="75" swimtime="00:01:18.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="130" swimtime="00:15:04.53" resultid="4698" lane="2" heatid="6717" entrytime="00:15:00.00" />
                <RESULT eventid="1411" points="189" reactiontime="+112" swimtime="00:03:42.08" resultid="4701" lane="2" heatid="7004" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.93" />
                    <SPLIT distance="50" swimtime="00:00:51.21" />
                    <SPLIT distance="75" swimtime="00:01:18.62" />
                    <SPLIT distance="100" swimtime="00:01:46.93" />
                    <SPLIT distance="125" swimtime="00:02:15.94" />
                    <SPLIT distance="150" swimtime="00:02:44.75" />
                    <SPLIT distance="175" swimtime="00:03:13.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="126" reactiontime="+107" swimtime="00:07:18.18" resultid="4700" lane="3" heatid="6900" entrytime="00:07:19.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.91" />
                    <SPLIT distance="50" swimtime="00:00:47.57" />
                    <SPLIT distance="75" swimtime="00:01:15.27" />
                    <SPLIT distance="100" swimtime="00:01:42.99" />
                    <SPLIT distance="125" swimtime="00:02:11.26" />
                    <SPLIT distance="150" swimtime="00:02:38.83" />
                    <SPLIT distance="175" swimtime="00:03:07.49" />
                    <SPLIT distance="200" swimtime="00:03:35.53" />
                    <SPLIT distance="225" swimtime="00:04:04.17" />
                    <SPLIT distance="250" swimtime="00:04:32.50" />
                    <SPLIT distance="275" swimtime="00:05:00.57" />
                    <SPLIT distance="300" swimtime="00:05:28.83" />
                    <SPLIT distance="325" swimtime="00:05:56.79" />
                    <SPLIT distance="350" swimtime="00:06:24.55" />
                    <SPLIT distance="375" swimtime="00:06:52.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="140" reactiontime="+113" swimtime="00:01:30.46" resultid="4699" lane="1" heatid="6831" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.14" />
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                    <SPLIT distance="75" swimtime="00:01:04.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-01-01" firstname="Jan" gender="M" lastname="Klapsia" nation="POL" athleteid="4705">
              <RESULTS>
                <RESULT eventid="1764" points="32" reactiontime="+133" swimtime="00:01:06.77" resultid="4710" lane="7" heatid="7336" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="30" reactiontime="+69" swimtime="00:02:48.30" resultid="4709" lane="3" heatid="7318" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:36.76" />
                    <SPLIT distance="50" swimtime="00:01:17.86" />
                    <SPLIT distance="75" swimtime="00:02:03.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="37" swimtime="00:01:12.91" resultid="4708" lane="4" heatid="7032" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:36.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="4706" lane="1" heatid="6830" entrytime="00:02:15.00" />
                <RESULT comment="K 8" eventid="1239" reactiontime="+140" status="DSQ" swimtime="00:01:13.88" resultid="4707" lane="7" heatid="6854" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:35.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Marian" gender="M" lastname="Otlik" nation="POL" athleteid="4711">
              <RESULTS>
                <RESULT eventid="1598" points="224" reactiontime="+68" swimtime="00:03:07.82" resultid="4716" lane="3" heatid="7076" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.46" />
                    <SPLIT distance="50" swimtime="00:00:37.37" />
                    <SPLIT distance="75" swimtime="00:01:02.34" />
                    <SPLIT distance="100" swimtime="00:01:29.26" />
                    <SPLIT distance="125" swimtime="00:01:56.73" />
                    <SPLIT distance="150" swimtime="00:02:24.34" />
                    <SPLIT distance="175" swimtime="00:02:47.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="158" reactiontime="+82" swimtime="00:01:33.11" resultid="4715" lane="1" heatid="7017" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.40" />
                    <SPLIT distance="50" swimtime="00:00:40.95" />
                    <SPLIT distance="75" swimtime="00:01:05.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="281" reactiontime="+73" swimtime="00:00:35.02" resultid="4717" lane="3" heatid="7285" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="329" reactiontime="+73" swimtime="00:01:08.15" resultid="4713" lane="5" heatid="6840" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.39" />
                    <SPLIT distance="50" swimtime="00:00:30.88" />
                    <SPLIT distance="75" swimtime="00:00:48.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="385" reactiontime="+63" swimtime="00:00:29.24" resultid="4718" lane="4" heatid="7345" entrytime="00:00:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="269" reactiontime="+80" swimtime="00:01:19.23" resultid="4712" lane="6" heatid="6739" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.61" />
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                    <SPLIT distance="75" swimtime="00:01:00.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" reactiontime="+75" status="DNF" swimtime="00:00:00.00" resultid="4714" heatid="6903" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.65" />
                    <SPLIT distance="50" swimtime="00:00:35.84" />
                    <SPLIT distance="75" swimtime="00:00:55.75" />
                    <SPLIT distance="100" swimtime="00:01:17.27" />
                    <SPLIT distance="125" swimtime="00:01:39.93" />
                    <SPLIT distance="150" swimtime="00:02:03.58" />
                    <SPLIT distance="175" swimtime="00:02:26.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1971-01-01" firstname="Sławomir" gender="M" lastname="Szurek" nation="POL" athleteid="4719">
              <RESULTS>
                <RESULT eventid="1598" points="229" reactiontime="+88" swimtime="00:03:06.54" resultid="4724" lane="1" heatid="7075" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.60" />
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                    <SPLIT distance="75" swimtime="00:01:05.71" />
                    <SPLIT distance="100" swimtime="00:01:30.45" />
                    <SPLIT distance="125" swimtime="00:01:56.83" />
                    <SPLIT distance="150" swimtime="00:02:24.55" />
                    <SPLIT distance="175" swimtime="00:02:46.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="153" reactiontime="+100" swimtime="00:03:29.24" resultid="4721" lane="8" heatid="6871" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.04" />
                    <SPLIT distance="50" swimtime="00:00:47.15" />
                    <SPLIT distance="75" swimtime="00:01:13.86" />
                    <SPLIT distance="100" swimtime="00:01:41.14" />
                    <SPLIT distance="125" swimtime="00:02:09.50" />
                    <SPLIT distance="150" swimtime="00:02:37.67" />
                    <SPLIT distance="175" swimtime="00:03:03.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="200" reactiontime="+97" swimtime="00:06:56.82" resultid="4726" lane="7" heatid="7361" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.59" />
                    <SPLIT distance="50" swimtime="00:00:45.17" />
                    <SPLIT distance="75" swimtime="00:01:11.74" />
                    <SPLIT distance="100" swimtime="00:01:39.53" />
                    <SPLIT distance="125" swimtime="00:02:07.35" />
                    <SPLIT distance="150" swimtime="00:02:34.72" />
                    <SPLIT distance="175" swimtime="00:03:03.34" />
                    <SPLIT distance="200" swimtime="00:03:30.99" />
                    <SPLIT distance="225" swimtime="00:04:00.17" />
                    <SPLIT distance="250" swimtime="00:04:28.37" />
                    <SPLIT distance="275" swimtime="00:04:57.45" />
                    <SPLIT distance="300" swimtime="00:05:26.87" />
                    <SPLIT distance="325" swimtime="00:05:49.95" />
                    <SPLIT distance="350" swimtime="00:06:12.26" />
                    <SPLIT distance="375" swimtime="00:06:35.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="258" reactiontime="+88" swimtime="00:05:45.62" resultid="4722" lane="3" heatid="6903" entrytime="00:05:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.30" />
                    <SPLIT distance="50" swimtime="00:00:37.38" />
                    <SPLIT distance="75" swimtime="00:00:57.97" />
                    <SPLIT distance="100" swimtime="00:01:19.14" />
                    <SPLIT distance="125" swimtime="00:01:40.75" />
                    <SPLIT distance="150" swimtime="00:02:02.91" />
                    <SPLIT distance="175" swimtime="00:02:25.18" />
                    <SPLIT distance="200" swimtime="00:02:47.71" />
                    <SPLIT distance="225" swimtime="00:03:10.24" />
                    <SPLIT distance="250" swimtime="00:03:32.70" />
                    <SPLIT distance="275" swimtime="00:03:54.88" />
                    <SPLIT distance="300" swimtime="00:04:17.82" />
                    <SPLIT distance="325" swimtime="00:04:40.52" />
                    <SPLIT distance="350" swimtime="00:05:03.14" />
                    <SPLIT distance="375" swimtime="00:05:26.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="235" swimtime="00:12:22.50" resultid="4720" lane="8" heatid="6719" entrytime="00:12:30.00" />
                <RESULT eventid="1564" points="258" reactiontime="+88" swimtime="00:02:41.63" resultid="4723" heatid="7058" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.99" />
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                    <SPLIT distance="75" swimtime="00:00:56.76" />
                    <SPLIT distance="100" swimtime="00:01:17.50" />
                    <SPLIT distance="125" swimtime="00:01:38.28" />
                    <SPLIT distance="150" swimtime="00:01:59.31" />
                    <SPLIT distance="175" swimtime="00:02:20.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="300" reactiontime="+86" swimtime="00:00:31.76" resultid="4725" lane="5" heatid="7342" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-01-01" firstname="Ewa" gender="F" lastname="Adamczyk" nation="POL" athleteid="4727">
              <RESULTS>
                <RESULT eventid="1747" points="197" reactiontime="+114" swimtime="00:00:41.16" resultid="4733" lane="3" heatid="7329" entrytime="00:00:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1409" points="225" reactiontime="+118" swimtime="00:03:50.49" resultid="4730" lane="7" heatid="6999" entrytime="00:04:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.12" />
                    <SPLIT distance="50" swimtime="00:00:51.98" />
                    <SPLIT distance="75" swimtime="00:01:20.86" />
                    <SPLIT distance="100" swimtime="00:01:50.41" />
                    <SPLIT distance="125" swimtime="00:02:20.25" />
                    <SPLIT distance="150" swimtime="00:02:50.59" />
                    <SPLIT distance="175" swimtime="00:03:21.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="131" reactiontime="+114" swimtime="00:03:45.72" resultid="4731" lane="6" heatid="7049" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.79" />
                    <SPLIT distance="50" swimtime="00:00:50.47" />
                    <SPLIT distance="75" swimtime="00:01:19.30" />
                    <SPLIT distance="100" swimtime="00:01:48.33" />
                    <SPLIT distance="125" swimtime="00:02:18.45" />
                    <SPLIT distance="150" swimtime="00:02:47.91" />
                    <SPLIT distance="175" swimtime="00:03:17.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="240" reactiontime="+90" swimtime="00:01:44.64" resultid="4732" lane="6" heatid="7297" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.16" />
                    <SPLIT distance="50" swimtime="00:00:49.50" />
                    <SPLIT distance="75" swimtime="00:01:16.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="267" reactiontime="+110" swimtime="00:00:47.04" resultid="4729" lane="4" heatid="6850" entrytime="00:00:49.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.92" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="04" eventid="1187" reactiontime="+73" status="DSQ" swimtime="00:01:35.07" resultid="4728" lane="2" heatid="6823" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.23" />
                    <SPLIT distance="50" swimtime="00:00:44.06" />
                    <SPLIT distance="75" swimtime="00:01:09.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1341" points="101" reactiontime="+141" swimtime="00:03:24.91" resultid="4742" lane="5" heatid="6985">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.28" />
                    <SPLIT distance="50" swimtime="00:01:11.73" />
                    <SPLIT distance="75" swimtime="00:01:38.96" />
                    <SPLIT distance="100" swimtime="00:02:08.47" />
                    <SPLIT distance="125" swimtime="00:02:25.45" />
                    <SPLIT distance="150" swimtime="00:02:46.69" />
                    <SPLIT distance="175" swimtime="00:03:03.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4705" number="1" reactiontime="+141" />
                    <RELAYPOSITION athleteid="4689" number="2" reactiontime="+70" />
                    <RELAYPOSITION athleteid="4711" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="4697" number="4" reactiontime="+69" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1177" status="DNS" swimtime="00:00:00.00" resultid="4743" lane="3" heatid="6807">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4697" number="1" />
                    <RELAYPOSITION athleteid="4705" number="2" />
                    <RELAYPOSITION athleteid="4689" number="3" />
                    <RELAYPOSITION athleteid="4711" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1615" status="DNS" swimtime="00:00:00.00" resultid="4744" heatid="7442" entrytime="00:02:18.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" />
                    <RELAYPOSITION athleteid="4719" number="2" />
                    <RELAYPOSITION athleteid="4727" number="3" />
                    <RELAYPOSITION athleteid="4711" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1815" status="DNS" swimtime="00:00:00.00" resultid="4745" lane="1" heatid="7503" entrytime="00:02:38.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" />
                    <RELAYPOSITION athleteid="4727" number="2" />
                    <RELAYPOSITION athleteid="4719" number="3" />
                    <RELAYPOSITION athleteid="4711" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="TROST" name="OTR Interkol Ostrów Wlkp" nation="POL">
          <CONTACT name="w" />
          <ATHLETES>
            <ATHLETE birthdate="1948-01-01" firstname="Henryk" gender="M" lastname="Wołowicz" nation="POL" athleteid="4752">
              <RESULTS>
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="4754" lane="1" heatid="7339" entrytime="00:00:35.00" />
                <RESULT eventid="1375" status="DNS" swimtime="00:00:00.00" resultid="4753" lane="8" heatid="6900" entrytime="00:08:00.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="BASTA" name="SKSP Barakuda Stargard Szczeciński" nation="POL">
          <CONTACT name="Ch" />
          <ATHLETES>
            <ATHLETE birthdate="1955-01-01" firstname="Jerzy" gender="M" lastname="Grzesiak" nation="POL" athleteid="4768">
              <RESULTS>
                <RESULT eventid="1143" points="122" swimtime="00:29:20.06" resultid="4769" lane="1" heatid="6749" entrytime="00:28:58.00" />
                <RESULT eventid="1496" points="91" reactiontime="+154" swimtime="00:00:54.23" resultid="4772" lane="4" heatid="7033" entrytime="00:00:54.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="143" reactiontime="+153" swimtime="00:03:16.55" resultid="4773" lane="1" heatid="7056" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.54" />
                    <SPLIT distance="50" swimtime="00:00:41.09" />
                    <SPLIT distance="75" swimtime="00:01:04.36" />
                    <SPLIT distance="100" swimtime="00:01:29.94" />
                    <SPLIT distance="125" swimtime="00:01:56.04" />
                    <SPLIT distance="150" swimtime="00:02:22.92" />
                    <SPLIT distance="175" swimtime="00:02:50.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="195" reactiontime="+110" swimtime="00:00:36.69" resultid="4775" lane="3" heatid="7339" entrytime="00:00:34.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="121" reactiontime="+109" swimtime="00:07:24.54" resultid="4771" lane="1" heatid="6901" entrytime="00:06:59.40">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.15" />
                    <SPLIT distance="50" swimtime="00:00:46.12" />
                    <SPLIT distance="75" swimtime="00:01:12.54" />
                    <SPLIT distance="100" swimtime="00:01:40.53" />
                    <SPLIT distance="125" swimtime="00:02:08.68" />
                    <SPLIT distance="150" swimtime="00:02:37.41" />
                    <SPLIT distance="175" swimtime="00:03:05.56" />
                    <SPLIT distance="200" swimtime="00:03:34.20" />
                    <SPLIT distance="225" swimtime="00:04:03.14" />
                    <SPLIT distance="250" swimtime="00:04:31.94" />
                    <SPLIT distance="275" swimtime="00:05:01.05" />
                    <SPLIT distance="300" swimtime="00:05:30.31" />
                    <SPLIT distance="325" swimtime="00:05:59.33" />
                    <SPLIT distance="350" swimtime="00:06:28.91" />
                    <SPLIT distance="375" swimtime="00:06:57.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="89" reactiontime="+137" swimtime="00:02:11.66" resultid="4774" lane="2" heatid="7303" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.24" />
                    <SPLIT distance="50" swimtime="00:01:02.12" />
                    <SPLIT distance="75" swimtime="00:01:37.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="185" reactiontime="+108" swimtime="00:01:22.47" resultid="4770" lane="4" heatid="6833" entrytime="00:01:19.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.60" />
                    <SPLIT distance="50" swimtime="00:00:38.98" />
                    <SPLIT distance="75" swimtime="00:01:00.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1956-01-01" firstname="Jerzy" gender="M" lastname="Chełstowski" nation="POL" athleteid="4776">
              <RESULTS>
                <RESULT eventid="1730" points="128" reactiontime="+156" swimtime="00:01:44.22" resultid="4782" lane="2" heatid="7320" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.82" />
                    <SPLIT distance="50" swimtime="00:00:52.18" />
                    <SPLIT distance="75" swimtime="00:01:19.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="181" swimtime="00:25:43.61" resultid="4777" lane="5" heatid="6749" entrytime="00:26:25.00" />
                <RESULT eventid="1798" points="150" reactiontime="+81" swimtime="00:07:38.46" resultid="4783" lane="3" heatid="7359" entrytime="00:07:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.16" />
                    <SPLIT distance="50" swimtime="00:00:46.80" />
                    <SPLIT distance="75" swimtime="00:01:14.25" />
                    <SPLIT distance="100" swimtime="00:01:42.99" />
                    <SPLIT distance="125" swimtime="00:02:15.25" />
                    <SPLIT distance="150" swimtime="00:02:46.32" />
                    <SPLIT distance="175" swimtime="00:03:17.95" />
                    <SPLIT distance="200" swimtime="00:03:49.67" />
                    <SPLIT distance="225" swimtime="00:04:20.81" />
                    <SPLIT distance="250" swimtime="00:04:52.11" />
                    <SPLIT distance="275" swimtime="00:05:24.01" />
                    <SPLIT distance="300" swimtime="00:05:55.21" />
                    <SPLIT distance="325" swimtime="00:06:22.09" />
                    <SPLIT distance="350" swimtime="00:06:50.10" />
                    <SPLIT distance="375" swimtime="00:07:15.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="166" reactiontime="+79" swimtime="00:03:27.63" resultid="4781" lane="3" heatid="7074" entrytime="00:03:19.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.04" />
                    <SPLIT distance="50" swimtime="00:00:42.61" />
                    <SPLIT distance="75" swimtime="00:01:11.41" />
                    <SPLIT distance="100" swimtime="00:01:39.92" />
                    <SPLIT distance="125" swimtime="00:02:10.24" />
                    <SPLIT distance="150" swimtime="00:02:41.09" />
                    <SPLIT distance="175" swimtime="00:03:06.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="180" reactiontime="+77" swimtime="00:06:29.18" resultid="4779" lane="6" heatid="6902" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.72" />
                    <SPLIT distance="50" swimtime="00:00:41.52" />
                    <SPLIT distance="75" swimtime="00:01:03.83" />
                    <SPLIT distance="100" swimtime="00:01:28.74" />
                    <SPLIT distance="125" swimtime="00:01:52.79" />
                    <SPLIT distance="150" swimtime="00:02:18.39" />
                    <SPLIT distance="175" swimtime="00:02:44.59" />
                    <SPLIT distance="200" swimtime="00:03:10.41" />
                    <SPLIT distance="225" swimtime="00:03:35.97" />
                    <SPLIT distance="250" swimtime="00:04:00.62" />
                    <SPLIT distance="275" swimtime="00:04:27.46" />
                    <SPLIT distance="300" swimtime="00:04:52.68" />
                    <SPLIT distance="325" swimtime="00:05:18.55" />
                    <SPLIT distance="350" swimtime="00:05:44.84" />
                    <SPLIT distance="375" swimtime="00:06:08.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="248" reactiontime="+79" swimtime="00:01:14.87" resultid="4778" lane="3" heatid="6833" entrytime="00:01:19.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.89" />
                    <SPLIT distance="50" swimtime="00:00:35.52" />
                    <SPLIT distance="75" swimtime="00:00:55.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" status="DNS" swimtime="00:00:00.00" resultid="4780" heatid="7017" entrytime="00:01:34.30" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TOTOR" name="Toruńczyk Toruń" nation="POL">
          <CONTACT name="d" />
          <ATHLETES>
            <ATHLETE birthdate="1980-01-01" firstname="Bartosz" gender="M" lastname="Dybowski" nation="POL" athleteid="4793">
              <RESULTS>
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="4794" lane="6" heatid="6735" entrytime="00:01:25.60" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="4795" lane="7" heatid="6863" entrytime="00:00:36.70" />
                <RESULT eventid="1496" status="DNS" swimtime="00:00:00.00" resultid="4796" lane="4" heatid="7038" entrytime="00:00:35.20" />
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="4797" lane="5" heatid="7344" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TSRUM" name="Tri-Saucony Rumia" nation="POL">
          <CONTACT name="g" />
        </CLUB>
        <CLUB type="CLUB" code="WOKAT" name="UKS Wodnik 29 Katowice" nation="POL">
          <CONTACT name="mr" />
          <ATHLETES>
            <ATHLETE birthdate="1981-01-01" firstname="Anna" gender="F" lastname="Duda" nation="POL" athleteid="4807">
              <RESULTS>
                <RESULT eventid="1747" points="517" reactiontime="+71" swimtime="00:00:29.85" resultid="4811" heatid="7335" entrytime="00:00:30.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="487" reactiontime="+83" swimtime="00:00:32.36" resultid="4810" lane="3" heatid="7280" entrytime="00:00:31.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1445" points="366" reactiontime="+91" swimtime="00:01:19.13" resultid="4809" lane="1" heatid="7014" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.87" />
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                    <SPLIT distance="75" swimtime="00:00:57.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="466" reactiontime="+95" swimtime="00:01:08.19" resultid="4808" lane="8" heatid="6828" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.76" />
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                    <SPLIT distance="75" swimtime="00:00:49.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1952-01-01" firstname="Krzysztof" gender="M" lastname="Kulczyk" nation="POL" athleteid="4817">
              <RESULTS>
                <RESULT eventid="1645" points="334" reactiontime="+86" swimtime="00:00:33.09" resultid="4820" lane="4" heatid="7288" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="221" reactiontime="+89" swimtime="00:01:23.33" resultid="4819" lane="4" heatid="7018" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.49" />
                    <SPLIT distance="50" swimtime="00:00:37.08" />
                    <SPLIT distance="75" swimtime="00:00:59.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="312" reactiontime="+88" swimtime="00:00:31.37" resultid="4821" lane="2" heatid="7343" entrytime="00:00:30.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="298" reactiontime="+103" swimtime="00:01:10.42" resultid="4818" lane="4" heatid="6835" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.43" />
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                    <SPLIT distance="75" swimtime="00:00:51.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Jerzy" gender="M" lastname="Mroziński" nation="POL" athleteid="4822">
              <RESULTS>
                <RESULT eventid="1411" points="326" reactiontime="+93" swimtime="00:03:05.26" resultid="4825" lane="3" heatid="7008" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.63" />
                    <SPLIT distance="50" swimtime="00:00:41.42" />
                    <SPLIT distance="75" swimtime="00:01:04.42" />
                    <SPLIT distance="100" swimtime="00:01:28.54" />
                    <SPLIT distance="125" swimtime="00:01:52.77" />
                    <SPLIT distance="150" swimtime="00:02:17.40" />
                    <SPLIT distance="175" swimtime="00:02:41.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="391" reactiontime="+85" swimtime="00:01:20.50" resultid="4827" lane="1" heatid="7309" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.91" />
                    <SPLIT distance="50" swimtime="00:00:37.31" />
                    <SPLIT distance="75" swimtime="00:00:58.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="415" reactiontime="+86" swimtime="00:00:36.43" resultid="4824" lane="3" heatid="6862" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="294" reactiontime="+93" swimtime="00:01:16.87" resultid="4823" heatid="6737" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.37" />
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                    <SPLIT distance="75" swimtime="00:00:57.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" status="DNS" swimtime="00:00:00.00" resultid="4826" lane="1" heatid="7077" entrytime="00:02:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1979-01-01" firstname="Edyta" gender="F" lastname="Mróz" nation="POL" athleteid="4828">
              <RESULTS>
                <RESULT eventid="1058" points="366" swimtime="00:11:30.33" resultid="4829" lane="7" heatid="6715" entrytime="00:12:00.00" />
                <RESULT eventid="1290" points="362" reactiontime="+82" swimtime="00:02:55.65" resultid="4831" lane="7" heatid="6879" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.31" />
                    <SPLIT distance="50" swimtime="00:00:39.91" />
                    <SPLIT distance="75" swimtime="00:01:01.91" />
                    <SPLIT distance="100" swimtime="00:01:24.46" />
                    <SPLIT distance="125" swimtime="00:01:47.37" />
                    <SPLIT distance="150" swimtime="00:02:10.67" />
                    <SPLIT distance="175" swimtime="00:02:33.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="336" reactiontime="+87" swimtime="00:02:45.06" resultid="4833" lane="3" heatid="7052" entrytime="00:02:38.13">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.80" />
                    <SPLIT distance="50" swimtime="00:00:36.34" />
                    <SPLIT distance="75" swimtime="00:00:55.88" />
                    <SPLIT distance="100" swimtime="00:01:18.34" />
                    <SPLIT distance="125" swimtime="00:01:42.48" />
                    <SPLIT distance="150" swimtime="00:02:03.69" />
                    <SPLIT distance="175" swimtime="00:02:24.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="348" reactiontime="+88" swimtime="00:00:36.19" resultid="4834" lane="4" heatid="7278" entrytime="00:00:37.49">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="382" reactiontime="+77" swimtime="00:01:20.93" resultid="4835" lane="4" heatid="7316" entrytime="00:01:22.72">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.74" />
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                    <SPLIT distance="75" swimtime="00:01:00.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="412" reactiontime="+75" swimtime="00:00:37.17" resultid="4832" lane="2" heatid="7030" entrytime="00:00:38.43">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="379" reactiontime="+87" swimtime="00:01:13.06" resultid="4830" lane="1" heatid="6827" entrytime="00:01:12.47">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.15" />
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                    <SPLIT distance="75" swimtime="00:00:53.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1940-01-01" firstname="Krystyna" gender="F" lastname="Nicpoń" nation="POL" athleteid="4840">
              <RESULTS>
                <RESULT comment="Rekord Polski " eventid="1713" points="138" reactiontime="+112" swimtime="00:01:53.66" resultid="4845" heatid="7314" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.75" />
                    <SPLIT distance="50" swimtime="00:00:54.08" />
                    <SPLIT distance="75" swimtime="00:01:23.17" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1479" points="142" reactiontime="+77" swimtime="00:00:52.97" resultid="4844" lane="4" heatid="7026" entrytime="00:00:54.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.95" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1358" points="104" reactiontime="+94" swimtime="00:08:32.59" resultid="4843" lane="1" heatid="6894" entrytime="00:09:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.92" />
                    <SPLIT distance="50" swimtime="00:00:55.35" />
                    <SPLIT distance="75" swimtime="00:01:27.57" />
                    <SPLIT distance="100" swimtime="00:02:02.19" />
                    <SPLIT distance="125" swimtime="00:02:35.60" />
                    <SPLIT distance="150" swimtime="00:03:08.60" />
                    <SPLIT distance="175" swimtime="00:03:41.00" />
                    <SPLIT distance="200" swimtime="00:04:14.23" />
                    <SPLIT distance="225" swimtime="00:04:47.47" />
                    <SPLIT distance="250" swimtime="00:05:20.50" />
                    <SPLIT distance="275" swimtime="00:05:53.35" />
                    <SPLIT distance="300" swimtime="00:06:26.10" />
                    <SPLIT distance="325" swimtime="00:06:58.78" />
                    <SPLIT distance="350" swimtime="00:07:31.56" />
                    <SPLIT distance="375" swimtime="00:08:02.31" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1058" points="86" swimtime="00:18:38.78" resultid="4841" lane="4" heatid="6713" entrytime="00:19:00.00" />
                <RESULT comment="Rekord Polski " eventid="1290" points="135" reactiontime="+80" swimtime="00:04:03.80" resultid="4842" lane="4" heatid="6876" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.01" />
                    <SPLIT distance="50" swimtime="00:00:55.73" />
                    <SPLIT distance="75" swimtime="00:01:25.58" />
                    <SPLIT distance="100" swimtime="00:01:56.81" />
                    <SPLIT distance="125" swimtime="00:02:29.25" />
                    <SPLIT distance="150" swimtime="00:03:01.68" />
                    <SPLIT distance="175" swimtime="00:03:33.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Tomasz" gender="M" lastname="Skoczylas" nation="POL" athleteid="4846">
              <RESULTS>
                <RESULT eventid="1143" points="373" swimtime="00:20:14.77" resultid="4847" lane="7" heatid="6752" entrytime="00:21:10.00" />
                <RESULT eventid="1496" points="398" reactiontime="+81" swimtime="00:00:33.25" resultid="4850" lane="6" heatid="7040" entrytime="00:00:33.05">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="329" reactiontime="+83" swimtime="00:02:44.90" resultid="4849" lane="3" heatid="6884" entrytime="00:02:57.75">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.04" />
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                    <SPLIT distance="75" swimtime="00:00:56.84" />
                    <SPLIT distance="100" swimtime="00:01:18.13" />
                    <SPLIT distance="125" swimtime="00:01:39.68" />
                    <SPLIT distance="150" swimtime="00:02:01.66" />
                    <SPLIT distance="175" swimtime="00:02:23.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="361" reactiontime="+85" swimtime="00:01:13.75" resultid="4852" lane="7" heatid="7324" entrytime="00:01:16.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.59" />
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                    <SPLIT distance="75" swimtime="00:00:54.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="411" reactiontime="+90" swimtime="00:02:18.44" resultid="4851" lane="2" heatid="7062" entrytime="00:02:26.32">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.97" />
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                    <SPLIT distance="75" swimtime="00:00:49.21" />
                    <SPLIT distance="100" swimtime="00:01:07.28" />
                    <SPLIT distance="125" swimtime="00:01:25.59" />
                    <SPLIT distance="150" swimtime="00:01:44.19" />
                    <SPLIT distance="175" swimtime="00:02:01.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="460" reactiontime="+86" swimtime="00:01:00.91" resultid="4848" lane="7" heatid="6843" entrytime="00:01:00.77">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.90" />
                    <SPLIT distance="50" swimtime="00:00:29.09" />
                    <SPLIT distance="75" swimtime="00:00:44.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="451" reactiontime="+85" swimtime="00:00:27.73" resultid="4853" lane="2" heatid="7348" entrytime="00:00:27.92">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Marcin" gender="M" lastname="Szczypiński" nation="POL" athleteid="4854">
              <RESULTS>
                <RESULT eventid="1375" points="589" reactiontime="+86" swimtime="00:04:22.47" resultid="4857" lane="3" heatid="6909" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.82" />
                    <SPLIT distance="50" swimtime="00:00:29.56" />
                    <SPLIT distance="75" swimtime="00:00:45.36" />
                    <SPLIT distance="100" swimtime="00:01:01.90" />
                    <SPLIT distance="125" swimtime="00:01:18.42" />
                    <SPLIT distance="150" swimtime="00:01:35.44" />
                    <SPLIT distance="175" swimtime="00:01:52.09" />
                    <SPLIT distance="200" swimtime="00:02:09.06" />
                    <SPLIT distance="225" swimtime="00:02:25.50" />
                    <SPLIT distance="250" swimtime="00:02:42.50" />
                    <SPLIT distance="275" swimtime="00:02:59.04" />
                    <SPLIT distance="300" swimtime="00:03:15.95" />
                    <SPLIT distance="325" swimtime="00:03:32.47" />
                    <SPLIT distance="350" swimtime="00:03:49.51" />
                    <SPLIT distance="375" swimtime="00:04:06.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="558" swimtime="00:09:17.09" resultid="4855" lane="4" heatid="6722" entrytime="00:09:00.00" />
                <RESULT eventid="1205" points="649" reactiontime="+80" swimtime="00:00:54.34" resultid="4856" lane="5" heatid="6846" entrytime="00:00:54.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.60" />
                    <SPLIT distance="50" swimtime="00:00:26.61" />
                    <SPLIT distance="75" swimtime="00:00:40.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="583" reactiontime="+80" swimtime="00:02:03.22" resultid="4858" lane="6" heatid="7066" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.18" />
                    <SPLIT distance="50" swimtime="00:00:28.11" />
                    <SPLIT distance="75" swimtime="00:00:43.56" />
                    <SPLIT distance="100" swimtime="00:00:59.63" />
                    <SPLIT distance="125" swimtime="00:01:15.46" />
                    <SPLIT distance="150" swimtime="00:01:31.80" />
                    <SPLIT distance="175" swimtime="00:01:47.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="628" reactiontime="+78" swimtime="00:00:26.81" resultid="4859" heatid="7294" entrytime="00:00:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1934-01-01" firstname="Maria" gender="F" lastname="Śmiglewska" nation="POL" athleteid="4860">
              <RESULTS>
                <RESULT eventid="1222" points="36" swimtime="00:01:31.63" resultid="4861" lane="1" heatid="6848" entrytime="00:01:28.06">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:45.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1409" points="39" swimtime="00:06:51.19" resultid="4862" lane="8" heatid="6998" entrytime="00:07:11.73">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:49.85" />
                    <SPLIT distance="50" swimtime="00:01:40.59" />
                    <SPLIT distance="75" swimtime="00:02:33.24" />
                    <SPLIT distance="100" swimtime="00:03:25.46" />
                    <SPLIT distance="125" swimtime="00:04:17.69" />
                    <SPLIT distance="150" swimtime="00:05:08.82" />
                    <SPLIT distance="175" swimtime="00:06:00.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="34" swimtime="00:03:19.56" resultid="4863" lane="8" heatid="7296" entrytime="00:03:15.85">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:48.14" />
                    <SPLIT distance="50" swimtime="00:01:38.19" />
                    <SPLIT distance="75" swimtime="00:02:29.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1932-01-01" firstname="Urszula" gender="F" lastname="Walkowicz" nation="POL" athleteid="4864">
              <RESULTS>
                <RESULT eventid="1747" points="61" reactiontime="+129" swimtime="00:01:00.67" resultid="4870" lane="6" heatid="7328" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="65" reactiontime="+90" swimtime="00:02:25.45" resultid="4869" lane="1" heatid="7313" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:31.86" />
                    <SPLIT distance="50" swimtime="00:01:10.09" />
                    <SPLIT distance="75" swimtime="00:01:50.00" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rekord Polski " eventid="1479" points="82" reactiontime="+92" swimtime="00:01:03.49" resultid="4868" lane="5" heatid="7025" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="55" reactiontime="+132" swimtime="00:10:33.12" resultid="4867" lane="8" heatid="6894" entrytime="00:13:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:31.14" />
                    <SPLIT distance="50" swimtime="00:01:07.38" />
                    <SPLIT distance="75" swimtime="00:01:47.87" />
                    <SPLIT distance="100" swimtime="00:02:28.40" />
                    <SPLIT distance="125" swimtime="00:03:09.14" />
                    <SPLIT distance="150" swimtime="00:03:50.35" />
                    <SPLIT distance="175" swimtime="00:04:31.19" />
                    <SPLIT distance="200" swimtime="00:05:11.67" />
                    <SPLIT distance="225" swimtime="00:05:53.72" />
                    <SPLIT distance="250" swimtime="00:06:34.21" />
                    <SPLIT distance="275" swimtime="00:07:15.43" />
                    <SPLIT distance="300" swimtime="00:07:56.15" />
                    <SPLIT distance="325" swimtime="00:08:37.75" />
                    <SPLIT distance="350" swimtime="00:09:18.25" />
                    <SPLIT distance="375" swimtime="00:09:57.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1058" points="52" swimtime="00:22:02.77" resultid="4865" lane="3" heatid="6713" entrytime="00:24:30.00" />
                <RESULT eventid="1290" points="58" reactiontime="+90" swimtime="00:05:23.29" resultid="4866" lane="4" heatid="6875" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:33.81" />
                    <SPLIT distance="50" swimtime="00:01:14.85" />
                    <SPLIT distance="75" swimtime="00:01:56.69" />
                    <SPLIT distance="100" swimtime="00:02:39.61" />
                    <SPLIT distance="125" swimtime="00:03:22.55" />
                    <SPLIT distance="150" swimtime="00:04:04.43" />
                    <SPLIT distance="175" swimtime="00:04:45.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Olga" gender="F" lastname="Załuska" nation="POL" athleteid="4871">
              <RESULTS>
                <RESULT eventid="1641" points="437" reactiontime="+71" swimtime="00:00:33.55" resultid="4873" lane="5" heatid="7280" entrytime="00:00:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1445" points="396" reactiontime="+78" swimtime="00:01:17.07" resultid="4872" lane="3" heatid="7014" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.18" />
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                    <SPLIT distance="75" swimtime="00:00:55.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" status="DNS" swimtime="00:00:00.00" resultid="4874" lane="5" heatid="7334" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1341" points="404" reactiontime="+79" swimtime="00:02:09.18" resultid="4875" lane="2" heatid="6987" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.07" />
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                    <SPLIT distance="75" swimtime="00:00:51.67" />
                    <SPLIT distance="100" swimtime="00:01:11.55" />
                    <SPLIT distance="125" swimtime="00:01:23.72" />
                    <SPLIT distance="150" swimtime="00:01:38.39" />
                    <SPLIT distance="175" swimtime="00:01:52.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4846" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="4822" number="2" reactiontime="+53" />
                    <RELAYPOSITION athleteid="4854" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="4817" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1615" reactiontime="+79" swimtime="00:01:55.78" resultid="4876" heatid="7443" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.07" />
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                    <SPLIT distance="75" swimtime="00:00:47.91" />
                    <SPLIT distance="100" swimtime="00:01:03.71" />
                    <SPLIT distance="125" swimtime="00:01:16.93" />
                    <SPLIT distance="150" swimtime="00:01:31.19" />
                    <SPLIT distance="175" swimtime="00:01:42.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4828" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="4807" number="2" reactiontime="+32" />
                    <RELAYPOSITION athleteid="4846" number="3" reactiontime="+30" />
                    <RELAYPOSITION athleteid="4854" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WARSZ" name="Warszawa" nation="POL">
          <CONTACT name="d" />
          <ATHLETES>
            <ATHLETE birthdate="1953-01-01" firstname="Bogdan" gender="M" lastname="Dubiński" nation="POL" athleteid="4880">
              <RESULTS>
                <RESULT eventid="1496" points="289" reactiontime="+74" swimtime="00:00:36.98" resultid="4884" lane="7" heatid="7037" entrytime="00:00:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="187" reactiontime="+90" swimtime="00:03:19.09" resultid="4883" lane="3" heatid="6883" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:01:11.34" />
                    <SPLIT distance="50" swimtime="00:00:46.71" />
                    <SPLIT distance="75" swimtime="00:02:03.00" />
                    <SPLIT distance="100" swimtime="00:01:37.12" />
                    <SPLIT distance="125" swimtime="00:02:54.70" />
                    <SPLIT distance="150" swimtime="00:02:28.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="227" reactiontime="+80" swimtime="00:01:26.12" resultid="4886" lane="7" heatid="7322" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.52" />
                    <SPLIT distance="50" swimtime="00:00:42.62" />
                    <SPLIT distance="75" swimtime="00:01:04.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="176" reactiontime="+99" swimtime="00:07:14.89" resultid="4887" lane="1" heatid="7359" entrytime="00:07:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.54" />
                    <SPLIT distance="50" swimtime="00:00:54.64" />
                    <SPLIT distance="75" swimtime="00:01:25.87" />
                    <SPLIT distance="100" swimtime="00:01:57.94" />
                    <SPLIT distance="125" swimtime="00:02:26.13" />
                    <SPLIT distance="150" swimtime="00:02:52.95" />
                    <SPLIT distance="175" swimtime="00:03:19.82" />
                    <SPLIT distance="200" swimtime="00:03:45.95" />
                    <SPLIT distance="225" swimtime="00:04:17.28" />
                    <SPLIT distance="250" swimtime="00:04:48.48" />
                    <SPLIT distance="275" swimtime="00:05:18.83" />
                    <SPLIT distance="300" swimtime="00:05:48.44" />
                    <SPLIT distance="325" swimtime="00:06:12.05" />
                    <SPLIT distance="350" swimtime="00:06:33.89" />
                    <SPLIT distance="375" swimtime="00:06:55.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="187" reactiontime="+97" swimtime="00:03:19.68" resultid="4885" lane="6" heatid="7075" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.32" />
                    <SPLIT distance="50" swimtime="00:00:44.15" />
                    <SPLIT distance="75" swimtime="00:01:10.20" />
                    <SPLIT distance="100" swimtime="00:01:34.97" />
                    <SPLIT distance="125" swimtime="00:02:05.77" />
                    <SPLIT distance="150" swimtime="00:02:35.56" />
                    <SPLIT distance="175" swimtime="00:02:59.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="202" reactiontime="+103" swimtime="00:01:27.07" resultid="4881" lane="7" heatid="6735" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.30" />
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                    <SPLIT distance="75" swimtime="00:01:05.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="273" reactiontime="+95" swimtime="00:01:12.47" resultid="4882" lane="5" heatid="6835" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.08" />
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                    <SPLIT distance="75" swimtime="00:00:52.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1928-01-01" firstname="Wiesław" gender="M" lastname="Osiński" nation="POL" athleteid="4909">
              <RESULTS>
                <RESULT eventid="1730" points="7" reactiontime="+103" swimtime="00:04:24.56" resultid="4911" lane="2" heatid="7318" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:55.89" />
                    <SPLIT distance="50" swimtime="00:02:04.10" />
                    <SPLIT distance="75" swimtime="00:03:13.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="6" reactiontime="+152" swimtime="00:02:13.01" resultid="4910" lane="5" heatid="7032" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:59.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WMWAR" name="WMT Warszawa" nation="POL">
          <CONTACT name="w" />
          <ATHLETES>
            <ATHLETE birthdate="1980-01-01" firstname="Maciej" gender="M" lastname="Szymański" nation="POL" athleteid="4763">
              <RESULTS>
                <RESULT eventid="1764" points="597" reactiontime="+71" swimtime="00:00:25.27" resultid="4766" heatid="7354" entrytime="00:00:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="528" reactiontime="+80" swimtime="00:00:30.27" resultid="4765" heatid="7043" entrytime="00:00:29.99">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="485" reactiontime="+77" swimtime="00:00:34.58" resultid="4764" lane="8" heatid="6866" entrytime="00:00:32.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-01-01" firstname="Mirosław" gender="M" lastname="Warchoł" nation="POL" athleteid="4896">
              <RESULTS>
                <RESULT eventid="1496" points="342" reactiontime="+70" swimtime="00:00:34.99" resultid="4900" lane="3" heatid="7038" entrytime="00:00:35.33">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="437" reactiontime="+80" swimtime="00:00:28.03" resultid="4903" lane="6" heatid="7346" entrytime="00:00:28.55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="372" reactiontime="+69" swimtime="00:01:13.02" resultid="4902" lane="1" heatid="7323" entrytime="00:01:19.88">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.24" />
                    <SPLIT distance="50" swimtime="00:00:35.40" />
                    <SPLIT distance="75" swimtime="00:00:54.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="361" reactiontime="+73" swimtime="00:02:39.90" resultid="4899" lane="8" heatid="6886" entrytime="00:02:44.15">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.32" />
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                    <SPLIT distance="75" swimtime="00:00:57.36" />
                    <SPLIT distance="100" swimtime="00:01:17.49" />
                    <SPLIT distance="125" swimtime="00:01:37.90" />
                    <SPLIT distance="150" swimtime="00:01:58.53" />
                    <SPLIT distance="175" swimtime="00:02:19.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="402" reactiontime="+83" swimtime="00:02:19.44" resultid="4901" lane="6" heatid="7063" entrytime="00:02:19.55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.35" />
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                    <SPLIT distance="75" swimtime="00:00:49.55" />
                    <SPLIT distance="100" swimtime="00:01:07.54" />
                    <SPLIT distance="125" swimtime="00:01:25.43" />
                    <SPLIT distance="150" swimtime="00:01:43.70" />
                    <SPLIT distance="175" swimtime="00:02:02.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="419" reactiontime="+84" swimtime="00:01:02.83" resultid="4898" lane="6" heatid="6840" entrytime="00:01:05.88">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.24" />
                    <SPLIT distance="50" swimtime="00:00:30.13" />
                    <SPLIT distance="75" swimtime="00:00:46.42" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Z 2" eventid="1109" reactiontime="+84" status="DSQ" swimtime="00:01:12.57" resultid="4897" heatid="6740" entrytime="00:01:13.55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.81" />
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                    <SPLIT distance="75" swimtime="00:00:56.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1341" points="467" reactiontime="+69" swimtime="00:02:03.02" resultid="6981" lane="5" heatid="6988" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.21" />
                    <SPLIT distance="50" swimtime="00:00:32.38" />
                    <SPLIT distance="75" swimtime="00:00:46.77" />
                    <SPLIT distance="100" swimtime="00:01:04.28" />
                    <SPLIT distance="125" swimtime="00:01:17.68" />
                    <SPLIT distance="150" swimtime="00:01:33.18" />
                    <SPLIT distance="175" swimtime="00:01:47.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2678" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="2666" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="2588" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="2536" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1341" points="547" reactiontime="+69" swimtime="00:01:56.73" resultid="6982" lane="2" heatid="6988" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.32" />
                    <SPLIT distance="50" swimtime="00:00:31.20" />
                    <SPLIT distance="75" swimtime="00:00:45.80" />
                    <SPLIT distance="100" swimtime="00:01:03.63" />
                    <SPLIT distance="125" swimtime="00:01:16.26" />
                    <SPLIT distance="150" swimtime="00:01:31.46" />
                    <SPLIT distance="175" swimtime="00:01:39.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2560" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="2651" number="2" reactiontime="+73" />
                    <RELAYPOSITION athleteid="2615" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="4763" number="4" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1341" points="203" reactiontime="+80" swimtime="00:02:42.39" resultid="6983" lane="5" heatid="6987" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:01:06.59" />
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                    <SPLIT distance="75" swimtime="00:01:50.45" />
                    <SPLIT distance="100" swimtime="00:01:33.41" />
                    <SPLIT distance="125" swimtime="00:02:26.28" />
                    <SPLIT distance="150" swimtime="00:02:11.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2598" number="1" reactiontime="+80" />
                    <RELAYPOSITION athleteid="2633" number="2" reactiontime="+95" />
                    <RELAYPOSITION athleteid="2581" number="3" reactiontime="-1" />
                    <RELAYPOSITION athleteid="2576" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1177" points="426" reactiontime="+90" swimtime="00:01:55.26" resultid="6659" lane="7" heatid="6808" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.32" />
                    <SPLIT distance="50" swimtime="00:00:27.41" />
                    <SPLIT distance="75" swimtime="00:00:42.10" />
                    <SPLIT distance="100" swimtime="00:00:58.35" />
                    <SPLIT distance="125" swimtime="00:01:12.91" />
                    <SPLIT distance="150" swimtime="00:01:29.33" />
                    <SPLIT distance="175" swimtime="00:01:41.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2666" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="2576" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="2536" number="3" reactiontime="+65" />
                    <RELAYPOSITION athleteid="2615" number="4" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1341" points="143" reactiontime="+76" swimtime="00:03:02.61" resultid="6984" lane="7" heatid="6986" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.39" />
                    <SPLIT distance="50" swimtime="00:00:58.46" />
                    <SPLIT distance="75" swimtime="00:01:21.34" />
                    <SPLIT distance="100" swimtime="00:01:46.32" />
                    <SPLIT distance="125" swimtime="00:02:01.60" />
                    <SPLIT distance="150" swimtime="00:02:21.17" />
                    <SPLIT distance="175" swimtime="00:02:40.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2528" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="2628" number="2" reactiontime="+103" />
                    <RELAYPOSITION athleteid="4896" number="3" reactiontime="+39" />
                    <RELAYPOSITION athleteid="2593" number="4" reactiontime="+91" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1324" points="347" reactiontime="+90" swimtime="00:02:34.12" resultid="6977" lane="3" heatid="6979" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.94" />
                    <SPLIT distance="50" swimtime="00:00:46.32" />
                    <SPLIT distance="75" swimtime="00:01:04.32" />
                    <SPLIT distance="100" swimtime="00:01:24.66" />
                    <SPLIT distance="125" swimtime="00:01:40.92" />
                    <SPLIT distance="150" swimtime="00:02:00.30" />
                    <SPLIT distance="175" swimtime="00:02:16.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2568" number="1" reactiontime="+90" />
                    <RELAYPOSITION athleteid="2622" number="2" reactiontime="+63" />
                    <RELAYPOSITION athleteid="2659" number="3" reactiontime="+51" />
                    <RELAYPOSITION athleteid="2685" number="4" reactiontime="+65" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1815" reactiontime="+66" swimtime="00:02:06.86" resultid="7499" lane="3" heatid="7504" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.31" />
                    <SPLIT distance="50" swimtime="00:00:29.29" />
                    <SPLIT distance="75" swimtime="00:00:43.34" />
                    <SPLIT distance="100" swimtime="00:01:00.48" />
                    <SPLIT distance="125" swimtime="00:01:16.44" />
                    <SPLIT distance="150" swimtime="00:01:35.69" />
                    <SPLIT distance="175" swimtime="00:01:50.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2615" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="2666" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="2659" number="3" reactiontime="+50" />
                    <RELAYPOSITION athleteid="2622" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1615" reactiontime="+93" swimtime="00:02:05.57" resultid="7268" lane="4" heatid="7443" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.23" />
                    <SPLIT distance="50" swimtime="00:00:31.92" />
                    <SPLIT distance="75" swimtime="00:00:46.32" />
                    <SPLIT distance="100" swimtime="00:01:02.77" />
                    <SPLIT distance="125" swimtime="00:01:19.00" />
                    <SPLIT distance="150" swimtime="00:01:37.37" />
                    <SPLIT distance="175" swimtime="00:01:51.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2638" number="1" reactiontime="+93" />
                    <RELAYPOSITION athleteid="2536" number="2" reactiontime="+63" />
                    <RELAYPOSITION athleteid="2685" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="2560" number="4" reactiontime="+72" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1815" reactiontime="+77" swimtime="00:02:24.04" resultid="7500" lane="2" heatid="7504" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.32" />
                    <SPLIT distance="50" swimtime="00:00:37.38" />
                    <SPLIT distance="75" swimtime="00:00:57.80" />
                    <SPLIT distance="100" swimtime="00:01:21.59" />
                    <SPLIT distance="125" swimtime="00:01:34.85" />
                    <SPLIT distance="150" swimtime="00:01:50.75" />
                    <SPLIT distance="175" swimtime="00:02:06.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2536" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="2568" number="2" reactiontime="+60" />
                    <RELAYPOSITION athleteid="2588" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="2685" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1615" status="DNS" swimtime="00:00:00.00" resultid="7269" lane="3" heatid="7443" entrytime="00:01:51.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2622" number="1" />
                    <RELAYPOSITION athleteid="2685" number="2" />
                    <RELAYPOSITION athleteid="2588" number="3" />
                    <RELAYPOSITION athleteid="4896" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1615" status="DNS" swimtime="00:00:00.00" resultid="7270" lane="8" heatid="7443" entrytime="00:02:07.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2610" number="1" />
                    <RELAYPOSITION athleteid="2568" number="2" />
                    <RELAYPOSITION athleteid="2555" number="3" />
                    <RELAYPOSITION athleteid="2560" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="1615" status="DNS" swimtime="00:00:00.00" resultid="7271" lane="1" heatid="7442" entrytime="00:02:15.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2672" number="1" />
                    <RELAYPOSITION athleteid="2654" number="2" />
                    <RELAYPOSITION athleteid="2643" number="3" />
                    <RELAYPOSITION athleteid="2598" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="WROCL" name="Wrocław" nation="POL">
          <CONTACT name="f" />
          <ATHLETES>
            <ATHLETE birthdate="1989-01-01" firstname="Bartłomiej" gender="M" lastname="Jankowski" nation="POL" athleteid="4905">
              <RESULTS>
                <RESULT eventid="1696" points="382" reactiontime="+95" swimtime="00:01:21.14" resultid="4906" lane="5" heatid="7308" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.08" />
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                    <SPLIT distance="75" swimtime="00:00:58.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="384" reactiontime="+95" swimtime="00:01:10.34" resultid="4908" lane="1" heatid="6737" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.60" />
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                    <SPLIT distance="75" swimtime="00:00:53.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="MIELE" name="Mielec" shortname="Miele">
          <ATHLETES>
            <ATHLETE birthdate="1988-01-01" firstname="Daniel" gender="M" lastname="Paduch" nation="POL" athleteid="4912">
              <RESULTS>
                <RESULT eventid="1273" points="556" reactiontime="+76" swimtime="00:02:16.23" resultid="4915" lane="3" heatid="6874" entrytime="00:02:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.68" />
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                    <SPLIT distance="75" swimtime="00:00:47.00" />
                    <SPLIT distance="100" swimtime="00:01:04.75" />
                    <SPLIT distance="125" swimtime="00:01:22.35" />
                    <SPLIT distance="150" swimtime="00:01:40.29" />
                    <SPLIT distance="175" swimtime="00:01:58.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="534" swimtime="00:09:25.10" resultid="4914" lane="3" heatid="6722" entrytime="00:09:16.00" />
                <RESULT eventid="1462" points="512" reactiontime="+76" swimtime="00:01:02.96" resultid="4917" heatid="7023" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.50" />
                    <SPLIT distance="50" swimtime="00:00:29.58" />
                    <SPLIT distance="75" swimtime="00:00:46.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="512" reactiontime="+74" swimtime="00:02:08.69" resultid="4918" lane="8" heatid="7066" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.62" />
                    <SPLIT distance="50" swimtime="00:00:29.18" />
                    <SPLIT distance="75" swimtime="00:00:45.47" />
                    <SPLIT distance="100" swimtime="00:01:02.20" />
                    <SPLIT distance="125" swimtime="00:01:18.58" />
                    <SPLIT distance="150" swimtime="00:01:35.70" />
                    <SPLIT distance="175" swimtime="00:01:52.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="543" reactiontime="+73" swimtime="00:04:29.72" resultid="4916" lane="2" heatid="6909" entrytime="00:04:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.93" />
                    <SPLIT distance="50" swimtime="00:00:30.15" />
                    <SPLIT distance="75" swimtime="00:00:47.06" />
                    <SPLIT distance="100" swimtime="00:01:04.08" />
                    <SPLIT distance="125" swimtime="00:01:20.91" />
                    <SPLIT distance="150" swimtime="00:01:38.20" />
                    <SPLIT distance="175" swimtime="00:01:55.27" />
                    <SPLIT distance="200" swimtime="00:02:12.82" />
                    <SPLIT distance="225" swimtime="00:02:29.70" />
                    <SPLIT distance="250" swimtime="00:02:46.85" />
                    <SPLIT distance="275" swimtime="00:03:04.01" />
                    <SPLIT distance="300" swimtime="00:03:21.75" />
                    <SPLIT distance="325" swimtime="00:03:39.03" />
                    <SPLIT distance="350" swimtime="00:03:56.41" />
                    <SPLIT distance="375" swimtime="00:04:13.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="4919" lane="3" heatid="7292" entrytime="00:00:28.40" />
                <RESULT eventid="1798" status="DNS" swimtime="00:00:00.00" resultid="4920" lane="4" heatid="7364" entrytime="00:04:58.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WOWASF" name="WOPR Warszawa SPORT-Figielski" nation="POL" region="MAZ">
          <CONTACT city="Warszawa" email="sport-figielski@o2.pl" fax="22-403-2788" internet="www.sport-figielski.pl" name="Grzegorz Figielski" phone="501-29-44-77" state="MAZ" street="Sarmacka 21 m. 41" zip="02-972" />
          <ATHLETES>
            <ATHLETE birthdate="1953-12-27" firstname="Grzegorz" gender="M" lastname="Figielski" nation="POL" athleteid="4923">
              <RESULTS>
                <RESULT eventid="1798" points="150" reactiontime="+105" swimtime="00:07:38.04" resultid="4929" heatid="7359" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.26" />
                    <SPLIT distance="50" swimtime="00:00:53.02" />
                    <SPLIT distance="75" swimtime="00:01:21.59" />
                    <SPLIT distance="100" swimtime="00:01:52.87" />
                    <SPLIT distance="125" swimtime="00:02:25.36" />
                    <SPLIT distance="150" swimtime="00:02:55.23" />
                    <SPLIT distance="175" swimtime="00:03:25.05" />
                    <SPLIT distance="200" swimtime="00:03:57.43" />
                    <SPLIT distance="225" swimtime="00:04:27.36" />
                    <SPLIT distance="250" swimtime="00:04:59.42" />
                    <SPLIT distance="275" swimtime="00:05:30.36" />
                    <SPLIT distance="300" swimtime="00:06:01.50" />
                    <SPLIT distance="325" swimtime="00:06:26.10" />
                    <SPLIT distance="350" swimtime="00:06:50.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="212" reactiontime="+94" swimtime="00:02:52.50" resultid="4927" lane="4" heatid="7055" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.31" />
                    <SPLIT distance="50" swimtime="00:00:38.68" />
                    <SPLIT distance="75" swimtime="00:00:59.50" />
                    <SPLIT distance="100" swimtime="00:01:21.56" />
                    <SPLIT distance="125" swimtime="00:01:43.64" />
                    <SPLIT distance="150" swimtime="00:02:06.86" />
                    <SPLIT distance="175" swimtime="00:02:30.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="203" reactiontime="+108" swimtime="00:06:14.12" resultid="4926" lane="4" heatid="6901" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.77" />
                    <SPLIT distance="50" swimtime="00:00:41.59" />
                    <SPLIT distance="75" swimtime="00:01:03.66" />
                    <SPLIT distance="100" swimtime="00:01:26.18" />
                    <SPLIT distance="125" swimtime="00:01:49.21" />
                    <SPLIT distance="150" swimtime="00:02:12.09" />
                    <SPLIT distance="175" swimtime="00:02:35.70" />
                    <SPLIT distance="200" swimtime="00:02:59.05" />
                    <SPLIT distance="225" swimtime="00:03:23.18" />
                    <SPLIT distance="250" swimtime="00:03:48.01" />
                    <SPLIT distance="275" swimtime="00:04:11.96" />
                    <SPLIT distance="300" swimtime="00:04:35.90" />
                    <SPLIT distance="325" swimtime="00:05:00.76" />
                    <SPLIT distance="350" swimtime="00:05:25.67" />
                    <SPLIT distance="375" swimtime="00:05:50.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="242" reactiontime="+97" swimtime="00:00:34.11" resultid="4928" lane="7" heatid="7340" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="4925" lane="6" heatid="6834" entrytime="00:01:15.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-02-05" firstname="Agata" gender="F" lastname="Figielska" nation="POL" athleteid="4930">
              <RESULTS>
                <RESULT eventid="1679" points="122" reactiontime="+113" swimtime="00:02:10.95" resultid="4933" lane="6" heatid="7296" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.99" />
                    <SPLIT distance="50" swimtime="00:01:02.86" />
                    <SPLIT distance="75" swimtime="00:01:38.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="137" reactiontime="+116" swimtime="00:00:58.75" resultid="4932" heatid="6849" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="70" reactiontime="+129" swimtime="00:00:58.01" resultid="4934" lane="4" heatid="7328" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="4931" lane="2" heatid="6822" entrytime="00:02:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1953-08-29" firstname="Michał" gender="M" lastname="Chojecki" nation="POL" athleteid="4935">
              <RESULTS>
                <RESULT eventid="1109" points="249" reactiontime="+98" swimtime="00:01:21.24" resultid="4936" lane="1" heatid="6736" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.30" />
                    <SPLIT distance="50" swimtime="00:00:39.42" />
                    <SPLIT distance="75" swimtime="00:01:02.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="230" reactiontime="+98" swimtime="00:03:06.28" resultid="4940" lane="4" heatid="7075" entrytime="00:03:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.50" />
                    <SPLIT distance="50" swimtime="00:00:39.40" />
                    <SPLIT distance="75" swimtime="00:01:04.31" />
                    <SPLIT distance="100" swimtime="00:01:30.01" />
                    <SPLIT distance="125" swimtime="00:01:56.87" />
                    <SPLIT distance="150" swimtime="00:02:23.70" />
                    <SPLIT distance="175" swimtime="00:02:45.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="305" reactiontime="+94" swimtime="00:01:27.48" resultid="4941" lane="1" heatid="7307" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.98" />
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                    <SPLIT distance="75" swimtime="00:01:04.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="334" reactiontime="+94" swimtime="00:00:30.67" resultid="4942" lane="5" heatid="7343" entrytime="00:00:30.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="264" reactiontime="+95" swimtime="00:03:18.55" resultid="4939" lane="4" heatid="7007" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.32" />
                    <SPLIT distance="50" swimtime="00:00:44.39" />
                    <SPLIT distance="75" swimtime="00:01:09.13" />
                    <SPLIT distance="100" swimtime="00:01:34.58" />
                    <SPLIT distance="125" swimtime="00:01:59.95" />
                    <SPLIT distance="150" swimtime="00:02:25.82" />
                    <SPLIT distance="175" swimtime="00:02:51.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="316" reactiontime="+100" swimtime="00:01:09.04" resultid="4937" lane="7" heatid="6836" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.21" />
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                    <SPLIT distance="75" swimtime="00:00:50.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="316" reactiontime="+94" swimtime="00:00:39.87" resultid="4938" lane="4" heatid="6858" entrytime="00:00:40.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1958-03-19" firstname="Andrzej" gender="M" lastname="Gryboś" nation="POL" athleteid="4943">
              <RESULTS>
                <RESULT eventid="1143" points="177" swimtime="00:25:57.44" resultid="4944" lane="8" heatid="6750" entrytime="00:24:30.00" />
                <RESULT eventid="1375" points="203" reactiontime="+99" swimtime="00:06:14.18" resultid="4945" lane="3" heatid="6902" entrytime="00:06:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.18" />
                    <SPLIT distance="50" swimtime="00:00:38.87" />
                    <SPLIT distance="75" swimtime="00:01:00.85" />
                    <SPLIT distance="100" swimtime="00:01:23.50" />
                    <SPLIT distance="125" swimtime="00:01:47.41" />
                    <SPLIT distance="150" swimtime="00:02:12.20" />
                    <SPLIT distance="175" swimtime="00:02:37.21" />
                    <SPLIT distance="200" swimtime="00:03:02.50" />
                    <SPLIT distance="225" swimtime="00:03:27.44" />
                    <SPLIT distance="250" swimtime="00:03:52.37" />
                    <SPLIT distance="275" swimtime="00:04:16.86" />
                    <SPLIT distance="300" swimtime="00:04:40.86" />
                    <SPLIT distance="325" swimtime="00:05:05.10" />
                    <SPLIT distance="350" swimtime="00:05:29.01" />
                    <SPLIT distance="375" swimtime="00:05:52.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="4946" lane="7" heatid="7058" entrytime="00:02:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-03-13" firstname="Alina" gender="F" lastname="Kraśniewska" nation="POL" athleteid="4947">
              <RESULTS>
                <RESULT eventid="1641" status="DNS" swimtime="00:00:00.00" resultid="4953" lane="6" heatid="7275" entrytime="00:01:22.00" />
                <RESULT eventid="1126" status="DNS" swimtime="00:00:00.00" resultid="4948" lane="1" heatid="6746" entrytime="00:40:00.00" />
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="4949" lane="4" heatid="6822" entrytime="00:02:00.00" />
                <RESULT eventid="1358" status="DNS" swimtime="00:00:00.00" resultid="4950" lane="6" heatid="6894" entrytime="00:08:56.00" />
                <RESULT eventid="1445" status="DNS" swimtime="00:00:00.00" resultid="4951" lane="6" heatid="7012" entrytime="00:03:30.00" />
                <RESULT eventid="1581" status="DNS" swimtime="00:00:00.00" resultid="4952" lane="5" heatid="7067" entrytime="00:05:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1945-03-07" firstname="Barbara" gender="F" lastname="Czabańska" nation="POL" athleteid="4954">
              <RESULTS>
                <RESULT eventid="1358" points="49" reactiontime="+112" swimtime="00:10:57.11" resultid="4957" heatid="6894" entrytime="00:10:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.88" />
                    <SPLIT distance="50" swimtime="00:02:41.31" />
                    <SPLIT distance="75" swimtime="00:01:57.69" />
                    <SPLIT distance="100" swimtime="00:04:06.33" />
                    <SPLIT distance="125" swimtime="00:03:23.37" />
                    <SPLIT distance="150" swimtime="00:05:29.95" />
                    <SPLIT distance="175" swimtime="00:04:47.90" />
                    <SPLIT distance="200" swimtime="00:06:52.99" />
                    <SPLIT distance="225" swimtime="00:06:11.42" />
                    <SPLIT distance="250" swimtime="00:08:18.02" />
                    <SPLIT distance="275" swimtime="00:07:33.95" />
                    <SPLIT distance="325" swimtime="00:08:58.87" />
                    <SPLIT distance="350" swimtime="00:09:41.43" />
                    <SPLIT distance="375" swimtime="00:10:20.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1445" points="12" reactiontime="+122" swimtime="00:04:06.47" resultid="4958" lane="2" heatid="7012" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:59.59" />
                    <SPLIT distance="50" swimtime="00:02:03.83" />
                    <SPLIT distance="75" swimtime="00:03:05.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="39" reactiontime="+136" swimtime="00:02:52.28" resultid="4955" lane="3" heatid="6723" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:41.97" />
                    <SPLIT distance="50" swimtime="00:01:34.32" />
                    <SPLIT distance="75" swimtime="00:02:16.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="52" reactiontime="+112" swimtime="00:02:21.64" resultid="4956" lane="6" heatid="6822" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.45" />
                    <SPLIT distance="50" swimtime="00:01:08.49" />
                    <SPLIT distance="75" swimtime="00:01:46.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1581" status="DNS" swimtime="00:00:00.00" resultid="4959" lane="2" heatid="7067" entrytime="00:06:00.00" />
                <RESULT eventid="1713" status="DNS" swimtime="00:00:00.00" resultid="4960" lane="6" heatid="7313" entrytime="00:02:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1942-01-05" firstname="Anna" gender="F" lastname="Zielińska" nation="POL" athleteid="4961">
              <RESULTS>
                <RESULT eventid="1290" points="48" reactiontime="+89" swimtime="00:05:42.63" resultid="4962" lane="7" heatid="6876" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:41.83" />
                    <SPLIT distance="50" swimtime="00:01:25.49" />
                    <SPLIT distance="75" swimtime="00:02:09.43" />
                    <SPLIT distance="100" swimtime="00:02:53.78" />
                    <SPLIT distance="125" swimtime="00:03:36.45" />
                    <SPLIT distance="150" swimtime="00:04:18.24" />
                    <SPLIT distance="175" swimtime="00:05:00.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="43" swimtime="00:05:26.67" resultid="4964" lane="3" heatid="7048" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.81" />
                    <SPLIT distance="50" swimtime="00:01:13.74" />
                    <SPLIT distance="75" swimtime="00:01:53.41" />
                    <SPLIT distance="100" swimtime="00:02:36.23" />
                    <SPLIT distance="125" swimtime="00:03:19.78" />
                    <SPLIT distance="150" swimtime="00:04:02.05" />
                    <SPLIT distance="175" swimtime="00:04:46.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="49" reactiontime="+88" swimtime="00:02:40.55" resultid="4965" lane="7" heatid="7313" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:37.65" />
                    <SPLIT distance="50" swimtime="00:01:17.34" />
                    <SPLIT distance="75" swimtime="00:01:58.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1409" points="63" swimtime="00:05:51.44" resultid="4963" heatid="6998" entrytime="00:06:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:41.29" />
                    <SPLIT distance="50" swimtime="00:01:23.76" />
                    <SPLIT distance="75" swimtime="00:02:07.71" />
                    <SPLIT distance="100" swimtime="00:02:52.11" />
                    <SPLIT distance="125" swimtime="00:03:38.02" />
                    <SPLIT distance="150" swimtime="00:04:22.39" />
                    <SPLIT distance="175" swimtime="00:05:07.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="51" swimtime="00:01:04.56" resultid="4966" lane="2" heatid="7328" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-02-25" firstname="Fabian" gender="M" lastname="Filipiak" nation="POL" athleteid="4967">
              <RESULTS>
                <RESULT eventid="1462" points="70" reactiontime="+90" swimtime="00:02:02.23" resultid="4970" lane="4" heatid="7015" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.50" />
                    <SPLIT distance="50" swimtime="00:00:55.71" />
                    <SPLIT distance="75" swimtime="00:01:28.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="93" swimtime="00:04:11.93" resultid="4971" lane="1" heatid="7072" entrytime="00:04:04.00" />
                <RESULT eventid="1307" points="84" reactiontime="+110" swimtime="00:04:19.29" resultid="4969" lane="8" heatid="6882" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.15" />
                    <SPLIT distance="50" swimtime="00:01:00.00" />
                    <SPLIT distance="75" swimtime="00:01:32.46" />
                    <SPLIT distance="100" swimtime="00:02:04.29" />
                    <SPLIT distance="125" swimtime="00:02:39.76" />
                    <SPLIT distance="150" swimtime="00:03:12.13" />
                    <SPLIT distance="175" swimtime="00:03:45.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="70" reactiontime="+95" swimtime="00:04:31.14" resultid="4968" lane="4" heatid="6869" entrytime="00:04:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.70" />
                    <SPLIT distance="50" swimtime="00:00:59.31" />
                    <SPLIT distance="75" swimtime="00:01:32.88" />
                    <SPLIT distance="100" swimtime="00:02:07.80" />
                    <SPLIT distance="125" swimtime="00:02:44.31" />
                    <SPLIT distance="150" swimtime="00:03:20.61" />
                    <SPLIT distance="175" swimtime="00:03:57.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="108" swimtime="00:16:01.43" resultid="6712" heatid="6718" entrytime="00:14:00.00" />
                <RESULT eventid="1798" points="92" reactiontime="+101" swimtime="00:08:59.23" resultid="4973" lane="2" heatid="7358" entrytime="00:08:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.83" />
                    <SPLIT distance="50" swimtime="00:01:03.64" />
                    <SPLIT distance="75" swimtime="00:01:38.83" />
                    <SPLIT distance="100" swimtime="00:02:14.05" />
                    <SPLIT distance="125" swimtime="00:02:48.05" />
                    <SPLIT distance="150" swimtime="00:03:24.15" />
                    <SPLIT distance="175" swimtime="00:03:59.12" />
                    <SPLIT distance="200" swimtime="00:04:32.07" />
                    <SPLIT distance="225" swimtime="00:05:09.89" />
                    <SPLIT distance="250" swimtime="00:05:46.01" />
                    <SPLIT distance="275" swimtime="00:06:23.63" />
                    <SPLIT distance="300" swimtime="00:07:00.62" />
                    <SPLIT distance="325" swimtime="00:07:29.84" />
                    <SPLIT distance="350" swimtime="00:08:00.16" />
                    <SPLIT distance="375" swimtime="00:08:30.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="74" reactiontime="+111" swimtime="00:02:05.13" resultid="4972" lane="2" heatid="7319" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.91" />
                    <SPLIT distance="50" swimtime="00:01:00.03" />
                    <SPLIT distance="75" swimtime="00:01:32.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-04-21" firstname="Damian" gender="M" lastname="Kądzielewski" nation="POL" athleteid="4974">
              <RESULTS>
                <RESULT eventid="1530" points="198" reactiontime="+97" swimtime="00:00:36.49" resultid="4975" lane="6" heatid="7047" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-10-01" firstname="Beata" gender="F" lastname="Kądzielewska" nation="POL" athleteid="4976">
              <RESULTS>
                <RESULT eventid="1581" points="249" reactiontime="+96" swimtime="00:03:24.17" resultid="4979" lane="7" heatid="7068" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.40" />
                    <SPLIT distance="50" swimtime="00:00:44.42" />
                    <SPLIT distance="75" swimtime="00:01:10.06" />
                    <SPLIT distance="100" swimtime="00:01:35.41" />
                    <SPLIT distance="125" swimtime="00:02:05.03" />
                    <SPLIT distance="150" swimtime="00:02:34.00" />
                    <SPLIT distance="175" swimtime="00:02:59.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="281" reactiontime="+76" swimtime="00:00:42.24" resultid="4978" lane="3" heatid="7028" entrytime="00:00:42.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="264" reactiontime="+72" swimtime="00:01:31.56" resultid="4980" lane="4" heatid="7315" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.40" />
                    <SPLIT distance="50" swimtime="00:00:44.62" />
                    <SPLIT distance="75" swimtime="00:01:08.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="263" reactiontime="+76" swimtime="00:03:15.36" resultid="4977" lane="1" heatid="6878" entrytime="00:03:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.73" />
                    <SPLIT distance="50" swimtime="00:00:44.40" />
                    <SPLIT distance="75" swimtime="00:01:08.54" />
                    <SPLIT distance="100" swimtime="00:01:33.69" />
                    <SPLIT distance="125" swimtime="00:01:59.13" />
                    <SPLIT distance="150" swimtime="00:02:25.20" />
                    <SPLIT distance="175" swimtime="00:02:50.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1177" points="198" reactiontime="+105" swimtime="00:02:28.86" resultid="4982" lane="8" heatid="6808" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.91" />
                    <SPLIT distance="50" swimtime="00:00:36.54" />
                    <SPLIT distance="75" swimtime="00:00:57.94" />
                    <SPLIT distance="100" swimtime="00:01:22.92" />
                    <SPLIT distance="125" swimtime="00:01:39.20" />
                    <SPLIT distance="150" swimtime="00:01:56.97" />
                    <SPLIT distance="175" swimtime="00:02:12.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4943" number="1" reactiontime="+105" />
                    <RELAYPOSITION athleteid="4967" number="2" reactiontime="+51" />
                    <RELAYPOSITION athleteid="4923" number="3" reactiontime="+57" />
                    <RELAYPOSITION athleteid="4935" number="4" reactiontime="+66" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1341" points="150" reactiontime="+104" swimtime="00:02:59.56" resultid="4984" lane="4" heatid="6985" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.83" />
                    <SPLIT distance="50" swimtime="00:00:58.62" />
                    <SPLIT distance="75" swimtime="00:01:18.72" />
                    <SPLIT distance="100" swimtime="00:01:41.31" />
                    <SPLIT distance="125" swimtime="00:01:59.44" />
                    <SPLIT distance="150" swimtime="00:02:20.06" />
                    <SPLIT distance="175" swimtime="00:02:38.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4967" number="1" reactiontime="+104" />
                    <RELAYPOSITION athleteid="4935" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="4923" number="3" reactiontime="+93" />
                    <RELAYPOSITION athleteid="4943" number="4" reactiontime="+90" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1160" points="76" swimtime="00:03:51.28" resultid="4981" lane="7" heatid="6813" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.21" />
                    <SPLIT distance="50" swimtime="00:01:07.09" />
                    <SPLIT distance="75" swimtime="00:01:38.87" />
                    <SPLIT distance="100" swimtime="00:02:12.80" />
                    <SPLIT distance="125" swimtime="00:02:40.20" />
                    <SPLIT distance="150" swimtime="00:03:11.63" />
                    <SPLIT distance="175" swimtime="00:03:30.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4961" number="1" />
                    <RELAYPOSITION athleteid="4954" number="2" reactiontime="+43" />
                    <RELAYPOSITION athleteid="4930" number="3" reactiontime="+106" />
                    <RELAYPOSITION athleteid="4976" number="4" reactiontime="+67" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="F" number="3">
              <RESULTS>
                <RESULT eventid="1324" points="66" reactiontime="+73" swimtime="00:04:27.80" resultid="4983" heatid="6979" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:33.20" />
                    <SPLIT distance="50" swimtime="00:01:11.61" />
                    <SPLIT distance="75" swimtime="00:01:37.65" />
                    <SPLIT distance="100" swimtime="00:02:08.69" />
                    <SPLIT distance="125" swimtime="00:02:54.96" />
                    <SPLIT distance="150" swimtime="00:03:47.66" />
                    <SPLIT distance="175" swimtime="00:04:07.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4961" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="4930" number="2" reactiontime="+36" />
                    <RELAYPOSITION athleteid="4954" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="4976" number="4" reactiontime="+78" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="X" number="5">
              <RESULTS>
                <RESULT eventid="1615" status="DNS" swimtime="00:00:00.00" resultid="4985" lane="2" heatid="7441" entrytime="00:03:00.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4947" number="1" />
                    <RELAYPOSITION athleteid="4954" number="2" />
                    <RELAYPOSITION athleteid="4923" number="3" />
                    <RELAYPOSITION athleteid="4935" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="X" number="6">
              <RESULTS>
                <RESULT eventid="1615" status="DNS" swimtime="00:00:00.00" resultid="4986" lane="5" heatid="7441" entrytime="00:03:00.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4961" number="1" />
                    <RELAYPOSITION athleteid="4967" number="2" />
                    <RELAYPOSITION athleteid="4976" number="3" />
                    <RELAYPOSITION athleteid="4943" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="X" number="7">
              <RESULTS>
                <RESULT eventid="1815" status="DNS" swimtime="00:00:00.00" resultid="4987" lane="7" heatid="7503" entrytime="00:03:30.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4954" number="1" />
                    <RELAYPOSITION athleteid="4935" number="2" />
                    <RELAYPOSITION athleteid="4923" number="3" />
                    <RELAYPOSITION athleteid="4947" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="X" number="8">
              <RESULTS>
                <RESULT eventid="1815" status="DNS" swimtime="00:00:00.00" resultid="4988" heatid="7503" entrytime="00:04:00.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4976" number="1" />
                    <RELAYPOSITION athleteid="4961" number="2" />
                    <RELAYPOSITION athleteid="4967" number="3" />
                    <RELAYPOSITION athleteid="4943" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="TRKOL" name="MLUKS Triathlon Koło">
          <ATHLETES>
            <ATHLETE birthdate="1962-01-01" firstname="Tomasz" gender="M" lastname="Brett" nation="POL" athleteid="5024">
              <RESULTS>
                <RESULT eventid="1143" points="312" swimtime="00:21:28.64" resultid="5026" lane="2" heatid="6752" entrytime="00:20:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WAPOZ" name="KS Warta Poznań" nation="POL" region="WIE">
          <CONTACT name="Jacek Thiem" />
          <ATHLETES>
            <ATHLETE birthdate="1963-02-17" firstname="Jacek" gender="M" lastname="Thiem" nation="POL" athleteid="5028">
              <RESULTS>
                <RESULT eventid="1075" points="232" swimtime="00:12:25.55" resultid="5029" heatid="6719" entrytime="00:12:30.00" />
                <RESULT eventid="1273" points="217" reactiontime="+106" swimtime="00:03:06.19" resultid="5031" lane="2" heatid="6872" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.34" />
                    <SPLIT distance="50" swimtime="00:00:42.19" />
                    <SPLIT distance="75" swimtime="00:01:05.51" />
                    <SPLIT distance="100" swimtime="00:01:29.15" />
                    <SPLIT distance="125" swimtime="00:01:52.92" />
                    <SPLIT distance="150" swimtime="00:02:17.29" />
                    <SPLIT distance="175" swimtime="00:02:41.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="185" reactiontime="+80" swimtime="00:01:32.07" resultid="5035" heatid="7322" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.15" />
                    <SPLIT distance="50" swimtime="00:00:45.97" />
                    <SPLIT distance="75" swimtime="00:01:09.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="210" reactiontime="+105" swimtime="00:01:24.77" resultid="5032" lane="2" heatid="7018" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.22" />
                    <SPLIT distance="50" swimtime="00:00:40.06" />
                    <SPLIT distance="75" swimtime="00:01:02.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="244" reactiontime="+90" swimtime="00:00:36.74" resultid="5034" lane="6" heatid="7285" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="240" reactiontime="+104" swimtime="00:02:45.61" resultid="5033" lane="3" heatid="7059" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.58" />
                    <SPLIT distance="50" swimtime="00:00:38.44" />
                    <SPLIT distance="75" swimtime="00:00:59.47" />
                    <SPLIT distance="100" swimtime="00:01:20.87" />
                    <SPLIT distance="125" swimtime="00:01:42.23" />
                    <SPLIT distance="150" swimtime="00:02:03.61" />
                    <SPLIT distance="175" swimtime="00:02:24.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="285" reactiontime="+93" swimtime="00:01:11.46" resultid="5030" heatid="6835" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.08" />
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                    <SPLIT distance="75" swimtime="00:00:52.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-01-01" firstname="Anna" gender="F" lastname="Kotecka" nation="POL" athleteid="5036">
              <RESULTS>
                <RESULT eventid="1058" points="268" swimtime="00:12:45.68" resultid="5037" lane="3" heatid="6714" entrytime="00:13:10.00" />
                <RESULT eventid="1358" points="288" swimtime="00:06:05.36" resultid="5039" lane="6" heatid="6896" entrytime="00:06:15.01">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.83" />
                    <SPLIT distance="50" swimtime="00:00:40.36" />
                    <SPLIT distance="75" swimtime="00:01:01.42" />
                    <SPLIT distance="100" swimtime="00:01:23.71" />
                    <SPLIT distance="125" swimtime="00:01:46.23" />
                    <SPLIT distance="150" swimtime="00:02:09.35" />
                    <SPLIT distance="175" swimtime="00:02:32.46" />
                    <SPLIT distance="200" swimtime="00:02:55.72" />
                    <SPLIT distance="225" swimtime="00:03:19.04" />
                    <SPLIT distance="250" swimtime="00:03:42.62" />
                    <SPLIT distance="275" swimtime="00:04:06.03" />
                    <SPLIT distance="300" swimtime="00:04:30.65" />
                    <SPLIT distance="325" swimtime="00:04:54.20" />
                    <SPLIT distance="350" swimtime="00:05:18.33" />
                    <SPLIT distance="375" swimtime="00:05:42.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="262" swimtime="00:00:37.44" resultid="5043" lane="1" heatid="7331" entrytime="00:00:37.46">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" points="297" swimtime="00:02:52.02" resultid="5041" lane="7" heatid="7051" entrytime="00:03:01.53">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.50" />
                    <SPLIT distance="50" swimtime="00:00:39.79" />
                    <SPLIT distance="75" swimtime="00:01:01.08" />
                    <SPLIT distance="100" swimtime="00:01:23.05" />
                    <SPLIT distance="125" swimtime="00:01:45.00" />
                    <SPLIT distance="150" swimtime="00:02:07.55" />
                    <SPLIT distance="175" swimtime="00:02:30.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="245" reactiontime="+98" swimtime="00:03:19.92" resultid="5038" heatid="6878" entrytime="00:03:20.82">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.51" />
                    <SPLIT distance="50" swimtime="00:00:46.74" />
                    <SPLIT distance="75" swimtime="00:01:11.44" />
                    <SPLIT distance="100" swimtime="00:01:37.34" />
                    <SPLIT distance="125" swimtime="00:02:04.04" />
                    <SPLIT distance="150" swimtime="00:02:29.76" />
                    <SPLIT distance="175" swimtime="00:02:56.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="242" reactiontime="+81" swimtime="00:01:34.18" resultid="5042" lane="5" heatid="7315" entrytime="00:01:33.79">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.50" />
                    <SPLIT distance="50" swimtime="00:00:45.93" />
                    <SPLIT distance="75" swimtime="00:01:10.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" status="DNS" swimtime="00:00:00.00" resultid="5040" lane="3" heatid="7027" entrytime="00:00:46.11" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-01" firstname="Paweł" gender="M" lastname="Olszewski" nation="POL" athleteid="5044">
              <RESULTS>
                <RESULT eventid="1764" points="488" reactiontime="+69" swimtime="00:00:27.02" resultid="5048" lane="5" heatid="7350" entrytime="00:00:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="424" reactiontime="+80" swimtime="00:02:16.99" resultid="5047" lane="5" heatid="7064" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.81" />
                    <SPLIT distance="50" swimtime="00:00:30.97" />
                    <SPLIT distance="75" swimtime="00:00:48.00" />
                    <SPLIT distance="100" swimtime="00:01:05.73" />
                    <SPLIT distance="125" swimtime="00:01:23.65" />
                    <SPLIT distance="150" swimtime="00:01:42.13" />
                    <SPLIT distance="175" swimtime="00:02:00.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="479" reactiontime="+79" swimtime="00:01:00.10" resultid="5046" lane="4" heatid="6843" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.63" />
                    <SPLIT distance="50" swimtime="00:00:28.35" />
                    <SPLIT distance="75" swimtime="00:00:43.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="344" reactiontime="+80" swimtime="00:01:12.95" resultid="5045" lane="8" heatid="6739" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.57" />
                    <SPLIT distance="50" swimtime="00:00:33.35" />
                    <SPLIT distance="75" swimtime="00:00:56.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-01-01" firstname="Piotr" gender="M" lastname="Kodur" nation="POL" athleteid="5049">
              <RESULTS>
                <RESULT eventid="1730" points="529" reactiontime="+65" swimtime="00:01:04.93" resultid="5056" lane="7" heatid="7325" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.32" />
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                    <SPLIT distance="75" swimtime="00:00:48.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="507" reactiontime="+70" swimtime="00:02:22.89" resultid="5052" lane="4" heatid="6885" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.92" />
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                    <SPLIT distance="75" swimtime="00:00:51.13" />
                    <SPLIT distance="100" swimtime="00:01:09.31" />
                    <SPLIT distance="125" swimtime="00:01:27.46" />
                    <SPLIT distance="150" swimtime="00:01:45.97" />
                    <SPLIT distance="175" swimtime="00:02:04.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="523" reactiontime="+77" swimtime="00:01:02.55" resultid="5053" lane="4" heatid="7022" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.02" />
                    <SPLIT distance="50" swimtime="00:00:28.71" />
                    <SPLIT distance="75" swimtime="00:00:45.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="566" reactiontime="+77" swimtime="00:00:32.85" resultid="5051" lane="5" heatid="6865" entrytime="00:00:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="501" reactiontime="+77" swimtime="00:01:04.39" resultid="5050" lane="2" heatid="6741" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.72" />
                    <SPLIT distance="50" swimtime="00:00:28.60" />
                    <SPLIT distance="75" swimtime="00:00:48.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="460" reactiontime="+81" swimtime="00:00:29.74" resultid="5055" lane="2" heatid="7289" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" status="DNS" swimtime="00:00:00.00" resultid="5054" lane="6" heatid="7080" entrytime="00:02:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1981-01-01" firstname="Piotr" gender="M" lastname="Kurek" nation="POL" athleteid="5057">
              <RESULTS>
                <RESULT eventid="1375" points="381" reactiontime="+69" swimtime="00:05:03.50" resultid="5059" lane="7" heatid="6907" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.76" />
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                    <SPLIT distance="75" swimtime="00:00:50.14" />
                    <SPLIT distance="100" swimtime="00:01:08.57" />
                    <SPLIT distance="125" swimtime="00:01:27.36" />
                    <SPLIT distance="150" swimtime="00:01:46.71" />
                    <SPLIT distance="175" swimtime="00:02:06.00" />
                    <SPLIT distance="200" swimtime="00:02:25.82" />
                    <SPLIT distance="225" swimtime="00:02:45.83" />
                    <SPLIT distance="250" swimtime="00:03:05.68" />
                    <SPLIT distance="275" swimtime="00:03:25.71" />
                    <SPLIT distance="300" swimtime="00:03:45.91" />
                    <SPLIT distance="325" swimtime="00:04:05.89" />
                    <SPLIT distance="350" swimtime="00:04:25.51" />
                    <SPLIT distance="375" swimtime="00:04:45.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="407" reactiontime="+65" swimtime="00:01:07.97" resultid="5060" lane="8" heatid="7021" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.21" />
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                    <SPLIT distance="75" swimtime="00:00:49.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="336" swimtime="00:10:59.25" resultid="5058" lane="2" heatid="6721" entrytime="00:11:00.00" />
                <RESULT eventid="1564" points="400" reactiontime="+67" swimtime="00:02:19.67" resultid="5061" lane="5" heatid="7061" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.92" />
                    <SPLIT distance="50" swimtime="00:00:29.92" />
                    <SPLIT distance="75" swimtime="00:00:47.11" />
                    <SPLIT distance="100" swimtime="00:01:05.00" />
                    <SPLIT distance="125" swimtime="00:01:23.39" />
                    <SPLIT distance="150" swimtime="00:01:42.70" />
                    <SPLIT distance="175" swimtime="00:02:01.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="456" reactiontime="+66" swimtime="00:00:29.81" resultid="5062" lane="4" heatid="7291" entrytime="00:00:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="463" reactiontime="+68" swimtime="00:00:27.49" resultid="5063" lane="4" heatid="7347" entrytime="00:00:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-01" firstname="Tomasz" gender="M" lastname="Rybak" nation="POL" athleteid="5064">
              <RESULTS>
                <RESULT eventid="1730" points="343" reactiontime="+71" swimtime="00:01:15.04" resultid="5070" lane="8" heatid="7323" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.58" />
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                    <SPLIT distance="75" swimtime="00:00:55.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="334" reactiontime="+69" swimtime="00:02:44.13" resultid="5066" lane="7" heatid="6884" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.76" />
                    <SPLIT distance="50" swimtime="00:00:36.62" />
                    <SPLIT distance="75" swimtime="00:00:56.42" />
                    <SPLIT distance="100" swimtime="00:01:16.86" />
                    <SPLIT distance="125" swimtime="00:01:38.62" />
                    <SPLIT distance="150" swimtime="00:02:00.44" />
                    <SPLIT distance="175" swimtime="00:02:22.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="332" reactiontime="+82" swimtime="00:02:44.86" resultid="5069" lane="2" heatid="7076" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.27" />
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                    <SPLIT distance="75" swimtime="00:00:52.96" />
                    <SPLIT distance="100" swimtime="00:01:14.19" />
                    <SPLIT distance="125" swimtime="00:01:39.93" />
                    <SPLIT distance="150" swimtime="00:02:05.51" />
                    <SPLIT distance="175" swimtime="00:02:25.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="345" reactiontime="+81" swimtime="00:01:11.80" resultid="5068" lane="7" heatid="7020" entrytime="00:01:16.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.15" />
                    <SPLIT distance="50" swimtime="00:00:33.16" />
                    <SPLIT distance="75" swimtime="00:00:52.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="326" reactiontime="+80" swimtime="00:01:14.26" resultid="5065" lane="3" heatid="6737" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.65" />
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                    <SPLIT distance="75" swimtime="00:00:57.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" status="DNS" swimtime="00:00:00.00" resultid="5071" lane="7" heatid="7362" entrytime="00:06:30.00" />
                <RESULT eventid="1375" status="DNS" swimtime="00:00:00.00" resultid="5067" lane="7" heatid="6906" entrytime="00:05:34.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1980-01-01" firstname="Błażej" gender="M" lastname="Wachowski" nation="POL" athleteid="5072">
              <RESULTS>
                <RESULT eventid="1798" points="177" swimtime="00:07:14.26" resultid="5079" lane="1" heatid="7360" entrytime="00:07:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.78" />
                    <SPLIT distance="50" swimtime="00:00:46.83" />
                    <SPLIT distance="75" swimtime="00:01:11.78" />
                    <SPLIT distance="100" swimtime="00:01:38.01" />
                    <SPLIT distance="125" swimtime="00:02:08.05" />
                    <SPLIT distance="150" swimtime="00:02:34.75" />
                    <SPLIT distance="175" swimtime="00:03:01.68" />
                    <SPLIT distance="200" swimtime="00:03:28.61" />
                    <SPLIT distance="225" swimtime="00:04:03.25" />
                    <SPLIT distance="250" swimtime="00:04:37.01" />
                    <SPLIT distance="275" swimtime="00:05:11.71" />
                    <SPLIT distance="300" swimtime="00:05:45.93" />
                    <SPLIT distance="325" swimtime="00:06:08.39" />
                    <SPLIT distance="350" swimtime="00:06:30.91" />
                    <SPLIT distance="375" swimtime="00:06:52.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="165" swimtime="00:03:23.86" resultid="5074" lane="1" heatid="6871" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.45" />
                    <SPLIT distance="50" swimtime="00:00:46.13" />
                    <SPLIT distance="75" swimtime="00:01:10.47" />
                    <SPLIT distance="100" swimtime="00:01:36.07" />
                    <SPLIT distance="125" swimtime="00:02:01.69" />
                    <SPLIT distance="150" swimtime="00:02:28.70" />
                    <SPLIT distance="175" swimtime="00:02:56.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="188" reactiontime="+111" swimtime="00:01:31.65" resultid="5078" lane="8" heatid="7321" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.53" />
                    <SPLIT distance="50" swimtime="00:00:45.43" />
                    <SPLIT distance="75" swimtime="00:01:09.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="172" swimtime="00:01:30.57" resultid="5076" lane="2" heatid="7017" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.66" />
                    <SPLIT distance="50" swimtime="00:00:42.31" />
                    <SPLIT distance="75" swimtime="00:01:05.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="238" swimtime="00:02:46.06" resultid="5077" lane="3" heatid="7056" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.26" />
                    <SPLIT distance="50" swimtime="00:00:39.29" />
                    <SPLIT distance="75" swimtime="00:01:00.30" />
                    <SPLIT distance="100" swimtime="00:01:21.69" />
                    <SPLIT distance="125" swimtime="00:01:42.99" />
                    <SPLIT distance="150" swimtime="00:02:04.20" />
                    <SPLIT distance="175" swimtime="00:02:25.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="237" swimtime="00:05:55.16" resultid="5075" lane="6" heatid="6903" entrytime="00:05:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.23" />
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                    <SPLIT distance="75" swimtime="00:01:01.19" />
                    <SPLIT distance="100" swimtime="00:01:23.18" />
                    <SPLIT distance="125" swimtime="00:01:45.63" />
                    <SPLIT distance="150" swimtime="00:02:07.60" />
                    <SPLIT distance="175" swimtime="00:02:30.13" />
                    <SPLIT distance="200" swimtime="00:02:52.92" />
                    <SPLIT distance="225" swimtime="00:03:15.57" />
                    <SPLIT distance="250" swimtime="00:03:38.60" />
                    <SPLIT distance="275" swimtime="00:04:01.87" />
                    <SPLIT distance="300" swimtime="00:04:25.30" />
                    <SPLIT distance="325" swimtime="00:04:48.17" />
                    <SPLIT distance="350" swimtime="00:05:11.29" />
                    <SPLIT distance="375" swimtime="00:05:33.41" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="przekroczony limit 12:15:00" eventid="1075" status="DSQ" swimtime="00:12:15.50" resultid="5073" lane="2" heatid="6720" entrytime="00:12:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="ADRIAN" gender="M" lastname="SOBKOWIAK" nation="POL" athleteid="5080">
              <RESULTS>
                <RESULT eventid="1696" points="229" reactiontime="+94" swimtime="00:01:36.17" resultid="5083" lane="7" heatid="7302" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.99" />
                    <SPLIT distance="50" swimtime="00:00:45.26" />
                    <SPLIT distance="75" swimtime="00:01:10.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="254" reactiontime="+85" swimtime="00:00:42.91" resultid="5081" lane="2" heatid="6857" entrytime="00:00:42.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" status="DNS" swimtime="00:00:00.00" resultid="5082" lane="2" heatid="7002" entrytime="00:05:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-01" firstname="RADOSŁAW" gender="M" lastname="SOBKOWIAK" nation="POL" athleteid="5084">
              <RESULTS>
                <RESULT eventid="1764" points="325" swimtime="00:00:30.93" resultid="5086" lane="2" heatid="7342" entrytime="00:00:31.00" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="5085" lane="5" heatid="6833" entrytime="00:01:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Grzegorz" gender="M" lastname="Witt" nation="POL" athleteid="5087">
              <RESULTS>
                <RESULT eventid="1375" points="184" reactiontime="+125" swimtime="00:06:26.86" resultid="5089" lane="8" heatid="6903" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.97" />
                    <SPLIT distance="50" swimtime="00:00:40.23" />
                    <SPLIT distance="75" swimtime="00:01:02.36" />
                    <SPLIT distance="100" swimtime="00:01:25.28" />
                    <SPLIT distance="125" swimtime="00:01:49.41" />
                    <SPLIT distance="150" swimtime="00:02:14.19" />
                    <SPLIT distance="175" swimtime="00:02:38.57" />
                    <SPLIT distance="200" swimtime="00:03:03.99" />
                    <SPLIT distance="225" swimtime="00:03:29.00" />
                    <SPLIT distance="250" swimtime="00:03:54.57" />
                    <SPLIT distance="275" swimtime="00:04:19.90" />
                    <SPLIT distance="300" swimtime="00:04:45.56" />
                    <SPLIT distance="325" swimtime="00:05:11.03" />
                    <SPLIT distance="350" swimtime="00:05:36.81" />
                    <SPLIT distance="375" swimtime="00:06:02.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="127" reactiontime="+82" swimtime="00:01:44.45" resultid="5092" lane="3" heatid="7320" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.38" />
                    <SPLIT distance="50" swimtime="00:00:51.58" />
                    <SPLIT distance="75" swimtime="00:01:18.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="103" reactiontime="+102" swimtime="00:04:02.58" resultid="5088" lane="1" heatid="6883" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.99" />
                    <SPLIT distance="50" swimtime="00:00:58.36" />
                    <SPLIT distance="75" swimtime="00:01:29.71" />
                    <SPLIT distance="100" swimtime="00:02:00.58" />
                    <SPLIT distance="125" swimtime="00:02:31.84" />
                    <SPLIT distance="150" swimtime="00:03:02.77" />
                    <SPLIT distance="175" swimtime="00:03:33.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="197" reactiontime="+123" swimtime="00:02:56.75" resultid="5090" lane="8" heatid="7057" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.27" />
                    <SPLIT distance="50" swimtime="00:00:38.89" />
                    <SPLIT distance="75" swimtime="00:01:00.76" />
                    <SPLIT distance="100" swimtime="00:01:23.44" />
                    <SPLIT distance="125" swimtime="00:01:47.42" />
                    <SPLIT distance="150" swimtime="00:02:10.70" />
                    <SPLIT distance="175" swimtime="00:02:34.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" status="DNS" swimtime="00:00:00.00" resultid="5093" lane="6" heatid="7360" entrytime="00:07:15.00" />
                <RESULT eventid="1598" status="DNS" swimtime="00:00:00.00" resultid="5091" lane="2" heatid="7072" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.67" />
                    <SPLIT distance="50" swimtime="00:00:59.68" />
                    <SPLIT distance="75" swimtime="00:01:30.19" />
                    <SPLIT distance="100" swimtime="00:02:03.21" />
                    <SPLIT distance="125" swimtime="00:02:40.19" />
                    <SPLIT distance="150" swimtime="00:03:16.48" />
                    <SPLIT distance="175" swimtime="00:03:43.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-01" firstname="Piotr" gender="M" lastname="Witt" nation="POL" athleteid="5094">
              <RESULTS>
                <RESULT eventid="1307" points="346" reactiontime="+71" swimtime="00:02:42.22" resultid="5097" lane="4" heatid="6886" entrytime="00:02:34.54">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.94" />
                    <SPLIT distance="50" swimtime="00:00:36.00" />
                    <SPLIT distance="75" swimtime="00:00:56.17" />
                    <SPLIT distance="100" swimtime="00:01:17.29" />
                    <SPLIT distance="125" swimtime="00:01:38.47" />
                    <SPLIT distance="150" swimtime="00:02:00.38" />
                    <SPLIT distance="175" swimtime="00:02:22.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="387" reactiontime="+70" swimtime="00:01:12.06" resultid="5100" lane="3" heatid="7324" entrytime="00:01:13.32">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.97" />
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                    <SPLIT distance="75" swimtime="00:00:53.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="417" reactiontime="+63" swimtime="00:00:32.73" resultid="5098" heatid="7041" entrytime="00:00:32.12">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="525" reactiontime="+81" swimtime="00:00:58.31" resultid="5096" lane="1" heatid="6844" entrytime="00:00:59.66">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.94" />
                    <SPLIT distance="50" swimtime="00:00:27.65" />
                    <SPLIT distance="75" swimtime="00:00:42.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="390" reactiontime="+86" swimtime="00:01:09.98" resultid="5095" lane="6" heatid="6737" entrytime="00:01:19.88">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.74" />
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                    <SPLIT distance="75" swimtime="00:00:53.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="518" reactiontime="+80" swimtime="00:00:26.48" resultid="5101" heatid="7350" entrytime="00:00:27.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" status="DNS" swimtime="00:00:00.00" resultid="5099" lane="7" heatid="7078" entrytime="00:02:45.91" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-01" firstname="Maciej" gender="M" lastname="Kopka" nation="POL" license="MOO11520002" athleteid="5102">
              <RESULTS>
                <RESULT eventid="1496" points="397" reactiontime="+73" swimtime="00:00:33.27" resultid="5107" lane="3" heatid="7035" entrytime="00:00:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="325" reactiontime="+70" swimtime="00:02:45.62" resultid="5105" lane="4" heatid="6883" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.44" />
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                    <SPLIT distance="75" swimtime="00:00:58.99" />
                    <SPLIT distance="100" swimtime="00:01:19.84" />
                    <SPLIT distance="125" swimtime="00:01:40.93" />
                    <SPLIT distance="150" swimtime="00:02:02.61" />
                    <SPLIT distance="175" swimtime="00:02:24.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="526" reactiontime="+76" swimtime="00:00:33.66" resultid="5104" lane="5" heatid="6859" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="323" reactiontime="+79" swimtime="00:03:05.82" resultid="5106" lane="2" heatid="7007" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.87" />
                    <SPLIT distance="50" swimtime="00:00:41.65" />
                    <SPLIT distance="75" swimtime="00:01:04.80" />
                    <SPLIT distance="100" swimtime="00:01:28.30" />
                    <SPLIT distance="125" swimtime="00:01:52.42" />
                    <SPLIT distance="150" swimtime="00:02:16.71" />
                    <SPLIT distance="175" swimtime="00:02:41.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="381" reactiontime="+79" swimtime="00:01:10.51" resultid="5103" lane="4" heatid="6733" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.43" />
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                    <SPLIT distance="75" swimtime="00:00:52.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="5109" lane="7" heatid="7339" entrytime="00:00:35.00" />
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="5108" lane="6" heatid="7283" entrytime="00:00:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1983-01-01" firstname="JAKUB" gender="M" lastname="STANOCH" nation="POL" athleteid="5110">
              <RESULTS>
                <RESULT eventid="1645" points="509" reactiontime="+61" swimtime="00:00:28.75" resultid="5112" lane="8" heatid="7293" entrytime="00:00:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="518" reactiontime="+62" swimtime="00:00:26.48" resultid="5113" heatid="7348" entrytime="00:00:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="5111" lane="5" heatid="6844" entrytime="00:00:59.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-01-01" firstname="Przemysław" gender="M" lastname="Isalski" nation="POL" athleteid="5114">
              <RESULTS>
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="5115" lane="7" heatid="7350" entrytime="00:00:27.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1947-01-01" firstname="Karol" gender="M" lastname="Ziółkowski" nation="POL" athleteid="5116">
              <RESULTS>
                <RESULT eventid="1764" points="96" reactiontime="+105" swimtime="00:00:46.40" resultid="5122" lane="8" heatid="7337" entrytime="00:00:46.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="5120" lane="8" heatid="7055" entrytime="00:03:50.00" />
                <RESULT comment="K 12" eventid="1696" reactiontime="+95" status="DSQ" swimtime="00:00:00.00" resultid="5121" lane="3" heatid="7302" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.30" />
                    <SPLIT distance="50" swimtime="00:00:56.63" />
                    <SPLIT distance="75" swimtime="00:01:30.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" status="DNS" swimtime="00:00:00.00" resultid="5119" lane="4" heatid="7002" entrytime="00:04:30.00" />
                <RESULT eventid="1375" status="DNS" swimtime="00:00:00.00" resultid="5118" lane="1" heatid="6900" entrytime="00:07:30.00" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="5117" heatid="6855" entrytime="00:00:52.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1984-01-01" firstname="Rafał" gender="M" lastname="Liszewski" nation="POL" athleteid="5123">
              <RESULTS>
                <RESULT eventid="1496" points="511" reactiontime="+76" swimtime="00:00:30.60" resultid="5126" lane="8" heatid="7040" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="574" reactiontime="+75" swimtime="00:00:25.60" resultid="5128" heatid="7351" entrytime="00:00:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="466" reactiontime="+77" swimtime="00:00:29.60" resultid="5127" heatid="7292" entrytime="00:00:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="5124" lane="4" heatid="6743" entrytime="00:01:07.00" />
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="5125" lane="4" heatid="6864" entrytime="00:00:34.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Jakub" gender="M" lastname="Romel" nation="POL" athleteid="5129">
              <RESULTS>
                <RESULT eventid="1798" points="461" reactiontime="+69" swimtime="00:05:15.43" resultid="5133" lane="6" heatid="7364" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.78" />
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="75" swimtime="00:00:50.73" />
                    <SPLIT distance="100" swimtime="00:01:09.98" />
                    <SPLIT distance="125" swimtime="00:01:30.97" />
                    <SPLIT distance="150" swimtime="00:01:51.15" />
                    <SPLIT distance="175" swimtime="00:02:11.23" />
                    <SPLIT distance="200" swimtime="00:02:31.35" />
                    <SPLIT distance="225" swimtime="00:02:54.13" />
                    <SPLIT distance="250" swimtime="00:03:17.17" />
                    <SPLIT distance="275" swimtime="00:03:39.92" />
                    <SPLIT distance="300" swimtime="00:04:03.36" />
                    <SPLIT distance="325" swimtime="00:04:22.41" />
                    <SPLIT distance="350" swimtime="00:04:40.84" />
                    <SPLIT distance="375" swimtime="00:04:58.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="415" reactiontime="+68" swimtime="00:02:30.15" resultid="5130" lane="2" heatid="6874" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.54" />
                    <SPLIT distance="50" swimtime="00:00:31.73" />
                    <SPLIT distance="75" swimtime="00:00:49.88" />
                    <SPLIT distance="100" swimtime="00:01:08.64" />
                    <SPLIT distance="125" swimtime="00:01:28.03" />
                    <SPLIT distance="150" swimtime="00:01:48.08" />
                    <SPLIT distance="175" swimtime="00:02:08.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="447" reactiontime="+69" swimtime="00:04:47.74" resultid="5131" lane="7" heatid="6908" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.12" />
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                    <SPLIT distance="75" swimtime="00:00:50.50" />
                    <SPLIT distance="100" swimtime="00:01:08.41" />
                    <SPLIT distance="125" swimtime="00:01:26.55" />
                    <SPLIT distance="150" swimtime="00:01:44.75" />
                    <SPLIT distance="175" swimtime="00:02:03.10" />
                    <SPLIT distance="200" swimtime="00:02:21.32" />
                    <SPLIT distance="225" swimtime="00:02:39.65" />
                    <SPLIT distance="250" swimtime="00:02:58.02" />
                    <SPLIT distance="275" swimtime="00:03:16.50" />
                    <SPLIT distance="300" swimtime="00:03:35.04" />
                    <SPLIT distance="325" swimtime="00:03:53.36" />
                    <SPLIT distance="350" swimtime="00:04:11.82" />
                    <SPLIT distance="375" swimtime="00:04:30.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="450" reactiontime="+68" swimtime="00:01:05.76" resultid="5132" lane="3" heatid="7022" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.13" />
                    <SPLIT distance="50" swimtime="00:00:30.59" />
                    <SPLIT distance="75" swimtime="00:00:48.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1982-01-01" firstname="MICHAŁ" gender="M" lastname="STOLARSKI" nation="POL" athleteid="5134">
              <RESULTS>
                <RESULT eventid="1205" points="500" reactiontime="+78" swimtime="00:00:59.27" resultid="5135" heatid="6845" entrytime="00:00:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.04" />
                    <SPLIT distance="50" swimtime="00:00:27.47" />
                    <SPLIT distance="75" swimtime="00:00:43.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="5137" lane="3" heatid="7347" entrytime="00:00:28.00" />
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="5136" lane="2" heatid="7065" entrytime="00:02:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-01" firstname="MARCIN" gender="M" lastname="STACHOWIAK" nation="POL" athleteid="5138">
              <RESULTS>
                <RESULT eventid="1411" points="492" reactiontime="+72" swimtime="00:02:41.45" resultid="5139" lane="5" heatid="7011" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.61" />
                    <SPLIT distance="50" swimtime="00:00:34.89" />
                    <SPLIT distance="75" swimtime="00:00:54.74" />
                    <SPLIT distance="100" swimtime="00:01:15.34" />
                    <SPLIT distance="125" swimtime="00:01:36.43" />
                    <SPLIT distance="150" swimtime="00:01:58.16" />
                    <SPLIT distance="175" swimtime="00:02:19.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="558" reactiontime="+74" swimtime="00:01:11.53" resultid="5140" lane="7" heatid="7311" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.94" />
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                    <SPLIT distance="75" swimtime="00:00:51.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="5141" lane="6" heatid="7353" entrytime="00:00:25.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-01" firstname="Michał" gender="M" lastname="Skrzypczak" nation="POL" athleteid="5142">
              <RESULTS>
                <RESULT eventid="1109" points="435" reactiontime="+76" swimtime="00:01:07.48" resultid="5143" lane="1" heatid="6743" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.31" />
                    <SPLIT distance="50" swimtime="00:00:30.45" />
                    <SPLIT distance="75" swimtime="00:00:50.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="494" reactiontime="+77" swimtime="00:00:29.04" resultid="5145" lane="4" heatid="7292" entrytime="00:00:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="494" reactiontime="+76" swimtime="00:00:59.48" resultid="5144" lane="5" heatid="6843" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.18" />
                    <SPLIT distance="50" swimtime="00:00:27.85" />
                    <SPLIT distance="75" swimtime="00:00:43.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="528" reactiontime="+73" swimtime="00:00:26.32" resultid="5146" lane="3" heatid="7351" entrytime="00:00:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1978-01-01" firstname="Marcin" gender="M" lastname="Chałupka" nation="RUS" athleteid="6701">
              <RESULTS>
                <RESULT eventid="1496" status="DNS" swimtime="00:00:00.00" resultid="6703" lane="6" heatid="7042" entrytime="00:00:30.50" />
                <RESULT eventid="1730" status="DNS" swimtime="00:00:00.00" resultid="6704" heatid="7325" entrytime="00:01:10.00" />
                <RESULT eventid="1307" status="DNS" swimtime="00:00:00.00" resultid="6702" lane="7" heatid="6886" entrytime="00:02:40.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1177" points="541" reactiontime="+67" swimtime="00:01:46.47" resultid="6658" lane="6" heatid="6810" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.87" />
                    <SPLIT distance="50" swimtime="00:00:27.17" />
                    <SPLIT distance="75" swimtime="00:00:39.67" />
                    <SPLIT distance="100" swimtime="00:00:53.42" />
                    <SPLIT distance="125" swimtime="00:01:05.73" />
                    <SPLIT distance="150" swimtime="00:01:19.51" />
                    <SPLIT distance="175" swimtime="00:01:32.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5114" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="5110" number="2" reactiontime="+50" />
                    <RELAYPOSITION athleteid="5049" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="5044" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1341" points="514" reactiontime="+70" swimtime="00:01:59.20" resultid="6660" lane="7" heatid="6987" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.43" />
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                    <SPLIT distance="75" swimtime="00:00:46.04" />
                    <SPLIT distance="100" swimtime="00:01:05.33" />
                    <SPLIT distance="125" swimtime="00:01:18.07" />
                    <SPLIT distance="150" swimtime="00:01:33.17" />
                    <SPLIT distance="175" swimtime="00:01:45.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5049" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="5102" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="5110" number="3" reactiontime="+46" />
                    <RELAYPOSITION athleteid="5142" number="4" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="159" agemin="120" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1177" points="524" reactiontime="+74" swimtime="00:01:47.64" resultid="1906" lane="8" heatid="6809" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.77" />
                    <SPLIT distance="50" swimtime="00:00:27.10" />
                    <SPLIT distance="75" swimtime="00:00:39.84" />
                    <SPLIT distance="100" swimtime="00:00:53.42" />
                    <SPLIT distance="125" swimtime="00:01:06.50" />
                    <SPLIT distance="150" swimtime="00:01:20.99" />
                    <SPLIT distance="175" swimtime="00:01:33.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5138" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="5142" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="5057" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="5129" number="4" reactiontime="+20" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1341" points="280" reactiontime="+105" swimtime="00:02:25.84" resultid="6661" lane="3" heatid="6986" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.27" />
                    <SPLIT distance="50" swimtime="00:00:43.26" />
                    <SPLIT distance="75" swimtime="00:01:00.55" />
                    <SPLIT distance="100" swimtime="00:01:21.05" />
                    <SPLIT distance="125" swimtime="00:01:38.86" />
                    <SPLIT distance="150" swimtime="00:01:59.03" />
                    <SPLIT distance="175" swimtime="00:02:11.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5072" number="1" reactiontime="+105" />
                    <RELAYPOSITION athleteid="5129" number="2" reactiontime="+26" />
                    <RELAYPOSITION athleteid="5028" number="3" reactiontime="+80" />
                    <RELAYPOSITION athleteid="5064" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="OLPOZ" name="TS Olimpia Poznań" nation="POL">
          <CONTACT name="Pietraszewski" />
          <ATHLETES>
            <ATHLETE birthdate="1939-01-01" firstname="Barbara" gender="F" lastname="Wojtuś- Nowak" nation="POL" athleteid="5148">
              <RESULTS>
                <RESULT eventid="1747" reactiontime="+98" status="DNS" swimtime="00:00:00.00" resultid="5149" heatid="7329" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1948-01-01" firstname="Teresa" gender="F" lastname="Barełkowska" nation="POL" athleteid="5150">
              <RESULTS>
                <RESULT eventid="1479" points="101" reactiontime="+77" swimtime="00:00:59.26" resultid="5152" lane="1" heatid="7026" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="178" reactiontime="+112" swimtime="00:00:53.84" resultid="5151" lane="5" heatid="6848" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" status="DNS" swimtime="00:00:00.00" resultid="5153" lane="3" heatid="7296" entrytime="00:02:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1950-01-01" firstname="Maria" gender="F" lastname="Łutowicz" nation="POL" athleteid="5154">
              <RESULTS>
                <RESULT eventid="1547" points="210" reactiontime="+95" swimtime="00:03:13.13" resultid="5157" lane="8" heatid="7051" entrytime="00:03:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.75" />
                    <SPLIT distance="50" swimtime="00:00:45.82" />
                    <SPLIT distance="75" swimtime="00:01:11.74" />
                    <SPLIT distance="100" swimtime="00:01:37.67" />
                    <SPLIT distance="125" swimtime="00:02:02.74" />
                    <SPLIT distance="150" swimtime="00:02:26.98" />
                    <SPLIT distance="175" swimtime="00:02:51.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="248" reactiontime="+91" swimtime="00:00:38.15" resultid="5159" lane="6" heatid="7331" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="181" reactiontime="+90" swimtime="00:01:43.84" resultid="5155" lane="5" heatid="6725" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.22" />
                    <SPLIT distance="50" swimtime="00:00:48.59" />
                    <SPLIT distance="75" swimtime="00:01:19.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="222" reactiontime="+93" swimtime="00:01:27.32" resultid="5156" lane="2" heatid="6824" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.48" />
                    <SPLIT distance="50" swimtime="00:00:41.24" />
                    <SPLIT distance="75" swimtime="00:01:04.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" status="DNS" swimtime="00:00:00.00" resultid="5158" heatid="7277" entrytime="00:00:49.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1954-01-01" firstname="Małgorzata" gender="F" lastname="Łasińska" nation="POL" athleteid="5160">
              <RESULTS>
                <RESULT eventid="1445" points="97" reactiontime="+110" swimtime="00:02:03.08" resultid="5163" lane="3" heatid="7012" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.09" />
                    <SPLIT distance="50" swimtime="00:00:56.87" />
                    <SPLIT distance="75" swimtime="00:01:29.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="124" reactiontime="+74" swimtime="00:01:57.62" resultid="5166" lane="5" heatid="7314" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.27" />
                    <SPLIT distance="50" swimtime="00:00:56.88" />
                    <SPLIT distance="75" swimtime="00:01:27.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1641" points="136" reactiontime="+106" swimtime="00:00:49.44" resultid="5165" lane="3" heatid="7276" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="106" reactiontime="+90" swimtime="00:04:24.31" resultid="5162" lane="7" heatid="6877" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.84" />
                    <SPLIT distance="75" swimtime="00:01:32.50" />
                    <SPLIT distance="125" swimtime="00:02:40.99" />
                    <SPLIT distance="175" swimtime="00:03:50.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="158" swimtime="00:01:48.58" resultid="5161" lane="2" heatid="6724" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.03" />
                    <SPLIT distance="50" swimtime="00:00:51.31" />
                    <SPLIT distance="75" swimtime="00:01:23.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1581" status="DNS" swimtime="00:00:00.00" resultid="5164" heatid="7068" entrytime="00:04:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Krystyna" gender="F" lastname="Strzelecka" nation="POL" athleteid="5167">
              <RESULTS>
                <RESULT eventid="1126" points="160" swimtime="00:28:54.50" resultid="5168" lane="3" heatid="6746" entrytime="00:30:00.00" />
                <RESULT eventid="1222" points="180" reactiontime="+94" swimtime="00:00:53.59" resultid="5170" lane="8" heatid="6849" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="185" reactiontime="+97" swimtime="00:01:32.76" resultid="5169" lane="6" heatid="6824" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.19" />
                    <SPLIT distance="50" swimtime="00:00:42.88" />
                    <SPLIT distance="75" swimtime="00:01:07.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="214" reactiontime="+94" swimtime="00:00:40.05" resultid="5171" lane="3" heatid="7330" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1957-01-01" firstname="Grażyna" gender="F" lastname="Cabaj-Drela" nation="POL" athleteid="5172">
              <RESULTS>
                <RESULT eventid="1092" points="323" reactiontime="+84" swimtime="00:01:25.67" resultid="5173" heatid="6728" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.63" />
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                    <SPLIT distance="75" swimtime="00:01:03.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="288" reactiontime="+82" swimtime="00:03:09.52" resultid="5175" lane="8" heatid="6879" entrytime="00:03:06.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.59" />
                    <SPLIT distance="50" swimtime="00:00:44.22" />
                    <SPLIT distance="75" swimtime="00:01:07.83" />
                    <SPLIT distance="100" swimtime="00:01:31.59" />
                    <SPLIT distance="125" swimtime="00:01:55.88" />
                    <SPLIT distance="150" swimtime="00:02:20.78" />
                    <SPLIT distance="175" swimtime="00:02:45.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="305" reactiontime="+77" swimtime="00:01:27.27" resultid="5177" lane="8" heatid="7316" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.05" />
                    <SPLIT distance="50" swimtime="00:00:42.61" />
                    <SPLIT distance="75" swimtime="00:01:05.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="332" reactiontime="+71" swimtime="00:00:39.93" resultid="5176" lane="1" heatid="7029" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="321" reactiontime="+78" swimtime="00:00:35.00" resultid="5178" lane="1" heatid="7333" entrytime="00:00:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1222" points="366" reactiontime="+84" swimtime="00:00:42.34" resultid="5174" lane="3" heatid="6852" entrytime="00:00:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1962-01-01" firstname="Ilona" gender="F" lastname="Kamińska" nation="POL" athleteid="5179">
              <RESULTS>
                <RESULT eventid="1222" points="391" reactiontime="+87" swimtime="00:00:41.42" resultid="5181" lane="5" heatid="6852" entrytime="00:00:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="302" reactiontime="+80" swimtime="00:01:27.62" resultid="5180" lane="5" heatid="6726" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.72" />
                    <SPLIT distance="50" swimtime="00:00:42.64" />
                    <SPLIT distance="75" swimtime="00:01:06.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-01" firstname="Paulina" gender="F" lastname="Nuckowska" nation="POL" athleteid="5182">
              <RESULTS>
                <RESULT eventid="1713" points="268" swimtime="00:01:31.09" resultid="5184" lane="4" heatid="7314" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.24" />
                    <SPLIT distance="50" swimtime="00:00:44.23" />
                    <SPLIT distance="75" swimtime="00:01:07.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="268" reactiontime="+95" swimtime="00:01:21.99" resultid="5183" lane="4" heatid="6824" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.24" />
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                    <SPLIT distance="75" swimtime="00:01:00.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1747" points="304" reactiontime="+88" swimtime="00:00:35.63" resultid="5185" heatid="7331" entrytime="00:00:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-01" firstname="Agnieszka" gender="F" lastname="Rybak-Starczak" nation="POL" athleteid="5186">
              <RESULTS>
                <RESULT eventid="1679" points="363" reactiontime="+93" swimtime="00:01:31.20" resultid="5189" lane="6" heatid="7299" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.85" />
                    <SPLIT distance="50" swimtime="00:00:43.73" />
                    <SPLIT distance="75" swimtime="00:01:07.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1409" points="330" reactiontime="+104" swimtime="00:03:22.71" resultid="5188" lane="3" heatid="7000" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.15" />
                    <SPLIT distance="50" swimtime="00:00:46.18" />
                    <SPLIT distance="75" swimtime="00:01:11.93" />
                    <SPLIT distance="100" swimtime="00:01:38.37" />
                    <SPLIT distance="125" swimtime="00:02:05.12" />
                    <SPLIT distance="150" swimtime="00:02:32.01" />
                    <SPLIT distance="175" swimtime="00:02:57.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="326" reactiontime="+94" swimtime="00:01:25.40" resultid="5187" lane="4" heatid="6727" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.95" />
                    <SPLIT distance="50" swimtime="00:00:40.33" />
                    <SPLIT distance="75" swimtime="00:01:05.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1934-01-01" firstname="Jan" gender="M" lastname="Kosmowski" nation="POL" athleteid="5190">
              <RESULTS>
                <RESULT eventid="1239" points="169" reactiontime="+102" swimtime="00:00:49.16" resultid="5191" lane="3" heatid="6855" entrytime="00:00:49.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-01" firstname="Katarzyna" gender="F" lastname="Kaczmarek" nation="POL" athleteid="5192">
              <RESULTS>
                <RESULT eventid="1747" status="DNS" swimtime="00:00:00.00" resultid="5194" lane="8" heatid="7331" entrytime="00:00:38.00" />
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="5193" lane="6" heatid="6714" entrytime="00:14:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1936-01-01" firstname="Zygmunt" gender="M" lastname="Bocian" nation="POL" athleteid="5195">
              <RESULTS>
                <RESULT eventid="1764" points="86" reactiontime="+107" swimtime="00:00:48.20" resultid="5198" lane="3" heatid="7336" entrytime="00:00:48.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="61" reactiontime="+81" swimtime="00:01:01.97" resultid="5197" lane="7" heatid="7033" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.63" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="K 8" eventid="1239" reactiontime="+116" status="DSQ" swimtime="00:01:01.17" resultid="5196" lane="6" heatid="6855" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1938-01-01" firstname="Lech" gender="M" lastname="Sarnowski" nation="POL" athleteid="5199">
              <RESULTS>
                <RESULT eventid="1496" points="104" reactiontime="+67" swimtime="00:00:51.92" resultid="5201" lane="2" heatid="7034" entrytime="00:00:49.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="187" reactiontime="+98" swimtime="00:00:47.46" resultid="5200" heatid="6856" entrytime="00:00:46.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="5203" heatid="7337" entrytime="00:00:43.00" />
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="5202" lane="5" heatid="7281" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1941-01-01" firstname="Maciej" gender="M" lastname="Durka" nation="POL" athleteid="5204">
              <RESULTS>
                <RESULT eventid="1496" points="103" reactiontime="+81" swimtime="00:00:52.06" resultid="5205" lane="1" heatid="7034" entrytime="00:00:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="5206" lane="1" heatid="7281" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1942-01-01" firstname="Bogusław" gender="M" lastname="Kujawa" nation="POL" athleteid="5207">
              <RESULTS>
                <RESULT eventid="1496" points="117" reactiontime="+94" swimtime="00:00:49.97" resultid="5210" lane="3" heatid="7034" entrytime="00:00:48.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="125" reactiontime="+76" swimtime="00:01:42.20" resultid="5208" heatid="6732" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.72" />
                    <SPLIT distance="50" swimtime="00:00:54.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="163" reactiontime="+84" swimtime="00:00:38.92" resultid="5211" lane="3" heatid="7337" entrytime="00:00:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="142" reactiontime="+86" swimtime="00:01:30.06" resultid="5209" lane="4" heatid="6831" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.73" />
                    <SPLIT distance="50" swimtime="00:00:40.58" />
                    <SPLIT distance="75" swimtime="00:01:04.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1942-01-01" firstname="Janisław" gender="M" lastname="Osięgłowski" nation="POL" athleteid="5212">
              <RESULTS>
                <RESULT eventid="1496" points="164" reactiontime="+91" swimtime="00:00:44.69" resultid="5213" lane="7" heatid="7035" entrytime="00:00:47.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1942-01-01" firstname="Zdzisław" gender="M" lastname="Gacek" nation="POL" athleteid="5214">
              <RESULTS>
                <RESULT eventid="1696" points="135" reactiontime="+105" swimtime="00:01:54.80" resultid="5217" lane="7" heatid="7304" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.87" />
                    <SPLIT distance="50" swimtime="00:00:52.38" />
                    <SPLIT distance="75" swimtime="00:01:22.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="174" reactiontime="+103" swimtime="00:00:48.62" resultid="5216" lane="7" heatid="6856" entrytime="00:00:46.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="152" reactiontime="+107" swimtime="00:00:39.83" resultid="5218" lane="1" heatid="7337" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="5215" lane="6" heatid="6831" entrytime="00:01:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1944-01-01" firstname="Jacek" gender="M" lastname="Lesiński" nation="POL" athleteid="5219">
              <RESULTS>
                <RESULT eventid="1307" points="161" reactiontime="+83" swimtime="00:03:29.26" resultid="5221" lane="7" heatid="6883" entrytime="00:03:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.13" />
                    <SPLIT distance="50" swimtime="00:00:47.83" />
                    <SPLIT distance="75" swimtime="00:01:13.79" />
                    <SPLIT distance="100" swimtime="00:01:41.10" />
                    <SPLIT distance="125" swimtime="00:02:08.79" />
                    <SPLIT distance="150" swimtime="00:02:36.68" />
                    <SPLIT distance="175" swimtime="00:03:04.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="173" reactiontime="+73" swimtime="00:01:34.21" resultid="5224" lane="5" heatid="7321" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.16" />
                    <SPLIT distance="50" swimtime="00:00:44.68" />
                    <SPLIT distance="75" swimtime="00:01:09.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="189" reactiontime="+107" swimtime="00:01:29.10" resultid="5220" lane="1" heatid="6733" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.76" />
                    <SPLIT distance="50" swimtime="00:00:41.53" />
                    <SPLIT distance="75" swimtime="00:01:07.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="184" reactiontime="+85" swimtime="00:00:42.99" resultid="5222" lane="6" heatid="7036" entrytime="00:00:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" status="DNS" swimtime="00:00:00.00" resultid="5223" lane="3" heatid="7073" entrytime="00:03:33.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-01" firstname="Henryk" gender="M" lastname="Ratajczak" nation="POL" athleteid="5225">
              <RESULTS>
                <RESULT eventid="1598" points="155" reactiontime="+117" swimtime="00:03:32.34" resultid="5229" heatid="7073" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.41" />
                    <SPLIT distance="50" swimtime="00:00:49.92" />
                    <SPLIT distance="75" swimtime="00:01:20.85" />
                    <SPLIT distance="100" swimtime="00:01:50.85" />
                    <SPLIT distance="125" swimtime="00:02:18.54" />
                    <SPLIT distance="150" swimtime="00:02:46.39" />
                    <SPLIT distance="175" swimtime="00:03:11.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="123" reactiontime="+93" swimtime="00:03:44.79" resultid="5227" lane="3" heatid="6869" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.55" />
                    <SPLIT distance="50" swimtime="00:00:49.66" />
                    <SPLIT distance="75" swimtime="00:01:17.99" />
                    <SPLIT distance="100" swimtime="00:01:47.20" />
                    <SPLIT distance="125" swimtime="00:02:16.45" />
                    <SPLIT distance="150" swimtime="00:02:46.09" />
                    <SPLIT distance="175" swimtime="00:03:16.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="228" reactiontime="+103" swimtime="00:01:36.35" resultid="5230" lane="4" heatid="7304" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.93" />
                    <SPLIT distance="50" swimtime="00:00:46.77" />
                    <SPLIT distance="75" swimtime="00:01:11.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="163" reactiontime="+103" swimtime="00:07:25.75" resultid="5231" lane="8" heatid="7359" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.22" />
                    <SPLIT distance="50" swimtime="00:00:52.08" />
                    <SPLIT distance="75" swimtime="00:01:21.19" />
                    <SPLIT distance="100" swimtime="00:01:50.26" />
                    <SPLIT distance="125" swimtime="00:02:22.15" />
                    <SPLIT distance="150" swimtime="00:02:52.41" />
                    <SPLIT distance="175" swimtime="00:03:23.13" />
                    <SPLIT distance="200" swimtime="00:03:53.07" />
                    <SPLIT distance="225" swimtime="00:04:20.83" />
                    <SPLIT distance="250" swimtime="00:04:47.89" />
                    <SPLIT distance="275" swimtime="00:05:15.19" />
                    <SPLIT distance="300" swimtime="00:05:42.58" />
                    <SPLIT distance="325" swimtime="00:06:09.57" />
                    <SPLIT distance="350" swimtime="00:06:36.06" />
                    <SPLIT distance="375" swimtime="00:07:02.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="216" reactiontime="+112" swimtime="00:03:32.47" resultid="5228" lane="1" heatid="7004" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.49" />
                    <SPLIT distance="50" swimtime="00:00:49.16" />
                    <SPLIT distance="75" swimtime="00:01:16.32" />
                    <SPLIT distance="100" swimtime="00:01:44.13" />
                    <SPLIT distance="125" swimtime="00:02:11.59" />
                    <SPLIT distance="150" swimtime="00:02:39.37" />
                    <SPLIT distance="175" swimtime="00:03:05.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="175" reactiontime="+104" swimtime="00:01:31.34" resultid="5226" lane="6" heatid="6732" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.21" />
                    <SPLIT distance="50" swimtime="00:00:44.78" />
                    <SPLIT distance="75" swimtime="00:01:10.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1951-01-01" firstname="Jerzy" gender="M" lastname="Boryski" nation="POL" athleteid="5232">
              <RESULTS>
                <RESULT eventid="1730" points="201" reactiontime="+65" swimtime="00:01:29.59" resultid="5236" lane="4" heatid="7321" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.31" />
                    <SPLIT distance="50" swimtime="00:00:44.08" />
                    <SPLIT distance="75" swimtime="00:01:07.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="226" reactiontime="+70" swimtime="00:00:40.14" resultid="5235" lane="3" heatid="7036" entrytime="00:00:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" status="DNS" swimtime="00:00:00.00" resultid="5234" lane="6" heatid="6883" entrytime="00:03:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Zbigniew" gender="M" lastname="Pietraszewski" nation="POL" athleteid="5237">
              <RESULTS>
                <RESULT eventid="1798" points="246" reactiontime="+94" swimtime="00:06:28.81" resultid="5239" lane="5" heatid="7361" entrytime="00:06:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.44" />
                    <SPLIT distance="50" swimtime="00:00:45.54" />
                    <SPLIT distance="75" swimtime="00:01:11.93" />
                    <SPLIT distance="100" swimtime="00:01:38.58" />
                    <SPLIT distance="125" swimtime="00:02:03.33" />
                    <SPLIT distance="150" swimtime="00:02:26.73" />
                    <SPLIT distance="175" swimtime="00:02:50.92" />
                    <SPLIT distance="200" swimtime="00:03:14.70" />
                    <SPLIT distance="225" swimtime="00:03:41.32" />
                    <SPLIT distance="250" swimtime="00:04:08.36" />
                    <SPLIT distance="275" swimtime="00:04:35.33" />
                    <SPLIT distance="300" swimtime="00:05:01.65" />
                    <SPLIT distance="325" swimtime="00:05:24.85" />
                    <SPLIT distance="350" swimtime="00:05:46.81" />
                    <SPLIT distance="375" swimtime="00:06:09.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="242" reactiontime="+92" swimtime="00:03:03.29" resultid="5238" lane="5" heatid="7076" entrytime="00:03:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.26" />
                    <SPLIT distance="50" swimtime="00:00:42.74" />
                    <SPLIT distance="75" swimtime="00:01:06.40" />
                    <SPLIT distance="100" swimtime="00:01:29.30" />
                    <SPLIT distance="125" swimtime="00:01:54.41" />
                    <SPLIT distance="150" swimtime="00:02:19.95" />
                    <SPLIT distance="175" swimtime="00:02:42.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Wojciech" gender="M" lastname="Niewitecki" nation="POL" athleteid="5240">
              <RESULTS>
                <RESULT eventid="1307" points="246" reactiontime="+78" swimtime="00:03:01.71" resultid="5241" lane="2" heatid="6884" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.62" />
                    <SPLIT distance="50" swimtime="00:00:43.67" />
                    <SPLIT distance="75" swimtime="00:01:06.28" />
                    <SPLIT distance="100" swimtime="00:01:29.63" />
                    <SPLIT distance="125" swimtime="00:01:53.25" />
                    <SPLIT distance="150" swimtime="00:02:17.09" />
                    <SPLIT distance="175" swimtime="00:02:40.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="284" reactiontime="+79" swimtime="00:01:19.84" resultid="5243" lane="7" heatid="7323" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.63" />
                    <SPLIT distance="50" swimtime="00:00:39.93" />
                    <SPLIT distance="75" swimtime="00:01:00.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="293" reactiontime="+81" swimtime="00:00:36.84" resultid="5242" lane="6" heatid="7037" entrytime="00:00:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1959-01-01" firstname="Marek" gender="M" lastname="Piekara" nation="POL" athleteid="5244">
              <RESULTS>
                <RESULT eventid="1075" points="304" swimtime="00:11:21.56" resultid="5245" lane="1" heatid="6720" entrytime="00:12:00.00" />
                <RESULT eventid="1798" points="280" reactiontime="+93" swimtime="00:06:12.42" resultid="5247" lane="5" heatid="7362" entrytime="00:06:19.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.04" />
                    <SPLIT distance="50" swimtime="00:00:39.24" />
                    <SPLIT distance="75" swimtime="00:01:01.60" />
                    <SPLIT distance="100" swimtime="00:01:25.08" />
                    <SPLIT distance="125" swimtime="00:01:51.93" />
                    <SPLIT distance="150" swimtime="00:02:17.65" />
                    <SPLIT distance="175" swimtime="00:02:43.43" />
                    <SPLIT distance="200" swimtime="00:03:08.95" />
                    <SPLIT distance="225" swimtime="00:03:35.11" />
                    <SPLIT distance="250" swimtime="00:04:01.09" />
                    <SPLIT distance="275" swimtime="00:04:26.90" />
                    <SPLIT distance="300" swimtime="00:04:52.50" />
                    <SPLIT distance="325" swimtime="00:05:13.99" />
                    <SPLIT distance="350" swimtime="00:05:34.24" />
                    <SPLIT distance="375" swimtime="00:05:53.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="305" reactiontime="+99" swimtime="00:05:26.89" resultid="5246" lane="1" heatid="6905" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.79" />
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                    <SPLIT distance="75" swimtime="00:00:57.13" />
                    <SPLIT distance="100" swimtime="00:01:17.43" />
                    <SPLIT distance="125" swimtime="00:01:37.87" />
                    <SPLIT distance="150" swimtime="00:01:58.42" />
                    <SPLIT distance="175" swimtime="00:02:19.07" />
                    <SPLIT distance="200" swimtime="00:02:40.11" />
                    <SPLIT distance="225" swimtime="00:03:01.16" />
                    <SPLIT distance="250" swimtime="00:03:22.34" />
                    <SPLIT distance="275" swimtime="00:03:43.07" />
                    <SPLIT distance="300" swimtime="00:04:04.15" />
                    <SPLIT distance="325" swimtime="00:04:24.76" />
                    <SPLIT distance="350" swimtime="00:04:45.99" />
                    <SPLIT distance="375" swimtime="00:05:07.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1949-01-01" firstname="Ryszard" gender="M" lastname="Krzyżanowski" nation="POL" athleteid="5248">
              <RESULTS>
                <RESULT eventid="1645" points="260" reactiontime="+100" swimtime="00:00:35.95" resultid="5251" lane="8" heatid="7285" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="201" swimtime="00:13:01.75" resultid="5249" lane="7" heatid="6718" entrytime="00:14:00.00" />
                <RESULT eventid="1205" points="275" reactiontime="+107" swimtime="00:01:12.30" resultid="5250" lane="6" heatid="6839" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.42" />
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="75" swimtime="00:00:52.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="5252" lane="3" heatid="7341" entrytime="00:00:32.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1966-01-01" firstname="Sławomir" gender="M" lastname="Cybertowicz" nation="POL" athleteid="5253">
              <RESULTS>
                <RESULT eventid="1411" points="382" reactiontime="+81" swimtime="00:02:55.72" resultid="5257" lane="6" heatid="7010" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.64" />
                    <SPLIT distance="50" swimtime="00:00:39.09" />
                    <SPLIT distance="75" swimtime="00:01:01.72" />
                    <SPLIT distance="100" swimtime="00:01:24.72" />
                    <SPLIT distance="125" swimtime="00:01:48.08" />
                    <SPLIT distance="150" swimtime="00:02:11.72" />
                    <SPLIT distance="175" swimtime="00:02:34.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="427" reactiontime="+79" swimtime="00:01:18.22" resultid="5259" heatid="7310" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.87" />
                    <SPLIT distance="50" swimtime="00:00:36.97" />
                    <SPLIT distance="75" swimtime="00:00:57.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="475" reactiontime="+80" swimtime="00:00:34.83" resultid="5255" lane="2" heatid="6864" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="384" reactiontime="+83" swimtime="00:02:21.65" resultid="5258" lane="3" heatid="7062" entrytime="00:02:23.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.01" />
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                    <SPLIT distance="75" swimtime="00:00:49.40" />
                    <SPLIT distance="100" swimtime="00:01:07.45" />
                    <SPLIT distance="125" swimtime="00:01:25.70" />
                    <SPLIT distance="150" swimtime="00:01:44.99" />
                    <SPLIT distance="175" swimtime="00:02:03.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="410" reactiontime="+82" swimtime="00:01:03.29" resultid="5254" lane="3" heatid="6841" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.02" />
                    <SPLIT distance="50" swimtime="00:00:30.09" />
                    <SPLIT distance="75" swimtime="00:00:46.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" status="DNS" swimtime="00:00:00.00" resultid="5256" lane="3" heatid="6907" entrytime="00:05:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1968-01-01" firstname="Radosław" gender="M" lastname="Pierz" nation="POL" athleteid="5260">
              <RESULTS>
                <RESULT eventid="1496" points="194" reactiontime="+80" swimtime="00:00:42.23" resultid="5263" lane="5" heatid="7035" entrytime="00:00:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="203" reactiontime="+82" swimtime="00:01:27.02" resultid="5261" lane="8" heatid="6736" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.60" />
                    <SPLIT distance="50" swimtime="00:00:39.33" />
                    <SPLIT distance="75" swimtime="00:01:03.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="306" reactiontime="+87" swimtime="00:00:40.33" resultid="5262" lane="8" heatid="6857" entrytime="00:00:44.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" status="DNS" swimtime="00:00:00.00" resultid="5264" lane="5" heatid="7074" entrytime="00:03:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1963-01-01" firstname="Przemysław" gender="M" lastname="Bekas" nation="POL" athleteid="5272">
              <RESULTS>
                <RESULT eventid="1764" points="418" reactiontime="+80" swimtime="00:00:28.44" resultid="5274" lane="7" heatid="7347" entrytime="00:00:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="351" reactiontime="+80" swimtime="00:00:38.52" resultid="5273" lane="3" heatid="6863" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1976-01-01" firstname="Norbert" gender="M" lastname="Szentner" nation="POL" athleteid="5275">
              <RESULTS>
                <RESULT eventid="1645" points="500" reactiontime="+81" swimtime="00:00:28.91" resultid="5280" lane="1" heatid="7293" entrytime="00:00:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="424" reactiontime="+81" swimtime="00:00:32.56" resultid="5279" lane="8" heatid="7039" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="363" reactiontime="+83" swimtime="00:01:13.60" resultid="5281" heatid="7324" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.57" />
                    <SPLIT distance="50" swimtime="00:00:36.05" />
                    <SPLIT distance="75" swimtime="00:00:55.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="358" reactiontime="+83" swimtime="00:01:10.96" resultid="5278" lane="2" heatid="7021" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.54" />
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                    <SPLIT distance="75" swimtime="00:00:51.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1972-01-01" firstname="Sława" gender="F" lastname="Mróz" nation="POL" athleteid="5282">
              <RESULTS>
                <RESULT eventid="1641" points="39" reactiontime="+105" swimtime="00:01:15.01" resultid="5286" lane="8" heatid="7276" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:33.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1713" points="46" reactiontime="+84" swimtime="00:02:43.58" resultid="5287" lane="3" heatid="7313" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:39.24" />
                    <SPLIT distance="50" swimtime="00:01:18.35" />
                    <SPLIT distance="75" swimtime="00:02:00.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1479" points="47" reactiontime="+92" swimtime="00:01:16.26" resultid="5284" lane="7" heatid="7026" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:37.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="78" reactiontime="+96" swimtime="00:02:03.68" resultid="5283" lane="8" heatid="6823" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.80" />
                    <SPLIT distance="50" swimtime="00:00:57.26" />
                    <SPLIT distance="75" swimtime="00:01:29.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1513" points="80" swimtime="00:00:55.43" resultid="7266" heatid="7044" />
                <RESULT eventid="1547" status="DNS" swimtime="00:00:00.00" resultid="5285" lane="1" heatid="7049" entrytime="00:04:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-01-01" firstname="Jacek" gender="M" lastname="Matyszczak" nation="POL" athleteid="6568" />
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1341" points="188" reactiontime="+75" swimtime="00:02:46.67" resultid="5292" lane="3" heatid="6985" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.45" />
                    <SPLIT distance="50" swimtime="00:00:42.83" />
                    <SPLIT distance="75" swimtime="00:01:01.91" />
                    <SPLIT distance="100" swimtime="00:01:23.66" />
                    <SPLIT distance="125" swimtime="00:01:43.61" />
                    <SPLIT distance="150" swimtime="00:02:06.15" />
                    <SPLIT distance="175" swimtime="00:02:25.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5219" number="1" reactiontime="+75" />
                    <RELAYPOSITION athleteid="5244" number="2" reactiontime="+76" />
                    <RELAYPOSITION athleteid="5225" number="3" reactiontime="+81" />
                    <RELAYPOSITION athleteid="5207" number="4" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1177" status="DNS" swimtime="00:00:00.00" resultid="5293" lane="5" heatid="6808" entrytime="00:02:05.00" />
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1341" points="254" reactiontime="+74" swimtime="00:02:30.74" resultid="5290" lane="5" heatid="6986" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.33" />
                    <SPLIT distance="50" swimtime="00:00:37.13" />
                    <SPLIT distance="75" swimtime="00:01:00.68" />
                    <SPLIT distance="100" swimtime="00:01:26.98" />
                    <SPLIT distance="125" swimtime="00:01:42.03" />
                    <SPLIT distance="150" swimtime="00:01:59.87" />
                    <SPLIT distance="175" swimtime="00:02:14.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5240" number="1" reactiontime="+74" />
                    <RELAYPOSITION athleteid="5272" number="2" reactiontime="+87" />
                    <RELAYPOSITION athleteid="5253" number="3" reactiontime="+63" />
                    <RELAYPOSITION athleteid="5248" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1177" points="202" reactiontime="+89" swimtime="00:02:27.78" resultid="5291" lane="4" heatid="6807" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.02" />
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                    <SPLIT distance="75" swimtime="00:00:57.72" />
                    <SPLIT distance="100" swimtime="00:01:19.68" />
                    <SPLIT distance="125" swimtime="00:01:37.28" />
                    <SPLIT distance="150" swimtime="00:01:56.85" />
                    <SPLIT distance="175" swimtime="00:02:11.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5207" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="5214" number="2" reactiontime="+81" />
                    <RELAYPOSITION athleteid="5219" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="5248" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1160" points="280" reactiontime="+85" swimtime="00:02:30.10" resultid="5294" lane="5" heatid="6813" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.95" />
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="75" swimtime="00:00:55.57" />
                    <SPLIT distance="100" swimtime="00:00:38.20" />
                    <SPLIT distance="125" swimtime="00:01:35.93" />
                    <SPLIT distance="150" swimtime="00:01:17.21" />
                    <SPLIT distance="175" swimtime="00:02:12.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5179" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="5160" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="5154" number="3" />
                    <RELAYPOSITION athleteid="5172" number="4" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1324" points="238" reactiontime="+76" swimtime="00:02:54.65" resultid="5295" lane="6" heatid="6979" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:01:12.12" />
                    <SPLIT distance="50" swimtime="00:00:52.25" />
                    <SPLIT distance="75" swimtime="00:01:53.78" />
                    <SPLIT distance="100" swimtime="00:01:35.21" />
                    <SPLIT distance="125" swimtime="00:02:34.66" />
                    <SPLIT distance="150" swimtime="00:02:16.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5160" number="1" reactiontime="+76" />
                    <RELAYPOSITION athleteid="5172" number="2" reactiontime="+59" />
                    <RELAYPOSITION athleteid="5179" number="3" reactiontime="+45" />
                    <RELAYPOSITION athleteid="5154" number="4" reactiontime="+75" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="5289" lane="6" heatid="6813" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:30.55" />
                    <SPLIT distance="100" swimtime="00:02:17.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1815" reactiontime="+73" swimtime="00:02:31.64" resultid="5297" lane="1" heatid="7502">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.42" />
                    <SPLIT distance="50" swimtime="00:00:40.55" />
                    <SPLIT distance="75" swimtime="00:00:58.71" />
                    <SPLIT distance="100" swimtime="00:01:19.57" />
                    <SPLIT distance="125" swimtime="00:01:34.30" />
                    <SPLIT distance="150" swimtime="00:01:52.25" />
                    <SPLIT distance="175" swimtime="00:02:10.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5172" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="5272" number="2" reactiontime="+73" />
                    <RELAYPOSITION athleteid="5253" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="5154" number="4" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1815" reactiontime="+63" swimtime="00:03:19.65" resultid="5299" lane="2" heatid="7502">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.14" />
                    <SPLIT distance="50" swimtime="00:00:58.00" />
                    <SPLIT distance="75" swimtime="00:01:23.20" />
                    <SPLIT distance="100" swimtime="00:01:51.95" />
                    <SPLIT distance="125" swimtime="00:02:12.04" />
                    <SPLIT distance="150" swimtime="00:02:36.20" />
                    <SPLIT distance="175" swimtime="00:02:57.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5150" number="1" reactiontime="+63" />
                    <RELAYPOSITION athleteid="5160" number="2" reactiontime="+76" />
                    <RELAYPOSITION athleteid="5225" number="3" reactiontime="+67" />
                    <RELAYPOSITION athleteid="5207" number="4" reactiontime="+81" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1615" reactiontime="+82" swimtime="00:02:12.51" resultid="5296" lane="5" heatid="7442" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.91" />
                    <SPLIT distance="50" swimtime="00:00:28.70" />
                    <SPLIT distance="75" swimtime="00:00:45.91" />
                    <SPLIT distance="100" swimtime="00:01:05.01" />
                    <SPLIT distance="125" swimtime="00:01:23.82" />
                    <SPLIT distance="150" swimtime="00:01:44.43" />
                    <SPLIT distance="175" swimtime="00:01:57.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5253" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="5172" number="2" reactiontime="+69" />
                    <RELAYPOSITION athleteid="5154" number="3" reactiontime="+77" />
                    <RELAYPOSITION athleteid="5275" number="4" reactiontime="+63" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="239" agemin="200" agetotalmax="-1" agetotalmin="-1" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="1615" swimtime="00:02:42.89" resultid="5298" lane="3" heatid="7440">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5240" number="1" />
                    <RELAYPOSITION athleteid="5160" number="2" />
                    <RELAYPOSITION athleteid="5282" number="3" />
                    <RELAYPOSITION athleteid="5248" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="279" agemin="240" agetotalmax="-1" agetotalmin="-1" gender="X" number="5">
              <RESULTS>
                <RESULT eventid="1615" reactiontime="+102" status="DNS" swimtime="00:00:00.00" resultid="5300" lane="4" heatid="7440">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.99" />
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                    <SPLIT distance="75" swimtime="00:00:54.97" />
                    <SPLIT distance="100" swimtime="00:01:17.61" />
                    <SPLIT distance="125" swimtime="00:01:43.51" />
                    <SPLIT distance="150" swimtime="00:02:11.71" />
                    <SPLIT distance="175" swimtime="00:02:26.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" reactiontime="+102" />
                    <RELAYPOSITION number="2" reactiontime="+66" />
                    <RELAYPOSITION number="3" reactiontime="+33" />
                    <RELAYPOSITION number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SSPOZ" name="SSI Start Poznań" nation="POL">
          <CONTACT name="Łukaszewicz" />
          <ATHLETES>
            <ATHLETE birthdate="1960-01-01" firstname="Jacek" gender="M" lastname="Adamski" nation="POL" athleteid="5328">
              <RESULTS>
                <RESULT eventid="1696" points="275" reactiontime="+111" swimtime="00:01:30.57" resultid="5331" lane="7" heatid="7307" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.69" />
                    <SPLIT distance="50" swimtime="00:00:42.46" />
                    <SPLIT distance="75" swimtime="00:01:06.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="260" reactiontime="+117" swimtime="00:03:19.66" resultid="5330" lane="1" heatid="7006" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.54" />
                    <SPLIT distance="50" swimtime="00:00:44.70" />
                    <SPLIT distance="75" swimtime="00:01:09.52" />
                    <SPLIT distance="100" swimtime="00:01:35.45" />
                    <SPLIT distance="125" swimtime="00:02:02.07" />
                    <SPLIT distance="150" swimtime="00:02:29.05" />
                    <SPLIT distance="175" swimtime="00:02:54.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="300" reactiontime="+118" swimtime="00:00:40.59" resultid="5329" lane="3" heatid="6859" entrytime="00:00:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1970-01-01" firstname="Tomasz" gender="M" lastname="Tobolski" nation="POL" athleteid="5332">
              <RESULTS>
                <RESULT eventid="1273" points="225" reactiontime="+82" swimtime="00:03:03.97" resultid="5335" lane="2" heatid="6873" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.22" />
                    <SPLIT distance="50" swimtime="00:00:37.57" />
                    <SPLIT distance="75" swimtime="00:00:59.89" />
                    <SPLIT distance="100" swimtime="00:01:23.82" />
                    <SPLIT distance="125" swimtime="00:01:49.00" />
                    <SPLIT distance="150" swimtime="00:02:14.57" />
                    <SPLIT distance="175" swimtime="00:02:40.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="398" reactiontime="+81" swimtime="00:00:36.93" resultid="5334" lane="3" heatid="6856" entrytime="00:00:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="322" reactiontime="+82" swimtime="00:01:14.55" resultid="5333" lane="8" heatid="6741" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.70" />
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="75" swimtime="00:00:56.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="375" reactiontime="+79" swimtime="00:00:31.82" resultid="5338" lane="4" heatid="7289" entrytime="00:00:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" points="293" reactiontime="+78" swimtime="00:00:36.82" resultid="5337" lane="4" heatid="7037" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="329" reactiontime="+76" swimtime="00:01:12.96" resultid="5336" lane="6" heatid="7020" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.04" />
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                    <SPLIT distance="75" swimtime="00:00:52.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1798" points="264" reactiontime="+81" swimtime="00:06:20.07" resultid="5339" lane="8" heatid="7363" entrytime="00:06:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.17" />
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                    <SPLIT distance="75" swimtime="00:00:56.45" />
                    <SPLIT distance="100" swimtime="00:01:18.25" />
                    <SPLIT distance="125" swimtime="00:01:43.14" />
                    <SPLIT distance="150" swimtime="00:02:08.71" />
                    <SPLIT distance="175" swimtime="00:02:33.60" />
                    <SPLIT distance="200" swimtime="00:02:58.68" />
                    <SPLIT distance="225" swimtime="00:03:25.88" />
                    <SPLIT distance="250" swimtime="00:03:53.62" />
                    <SPLIT distance="275" swimtime="00:04:21.90" />
                    <SPLIT distance="300" swimtime="00:04:50.87" />
                    <SPLIT distance="325" swimtime="00:05:13.54" />
                    <SPLIT distance="350" swimtime="00:05:36.41" />
                    <SPLIT distance="375" swimtime="00:05:59.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1975-01-01" firstname="Tomasz" gender="M" lastname="Lutkowski" nation="POL" athleteid="5340">
              <RESULTS>
                <RESULT eventid="1273" points="186" reactiontime="+111" swimtime="00:03:16.14" resultid="5342" lane="2" heatid="6870" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.93" />
                    <SPLIT distance="50" swimtime="00:00:43.23" />
                    <SPLIT distance="75" swimtime="00:01:07.53" />
                    <SPLIT distance="100" swimtime="00:01:32.70" />
                    <SPLIT distance="125" swimtime="00:01:58.14" />
                    <SPLIT distance="150" swimtime="00:02:23.49" />
                    <SPLIT distance="175" swimtime="00:02:49.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1462" points="259" reactiontime="+101" swimtime="00:01:18.99" resultid="5343" lane="2" heatid="7019" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.42" />
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                    <SPLIT distance="75" swimtime="00:00:55.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="287" reactiontime="+93" swimtime="00:02:35.92" resultid="5344" lane="6" heatid="7060" entrytime="00:02:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.56" />
                    <SPLIT distance="50" swimtime="00:00:34.89" />
                    <SPLIT distance="75" swimtime="00:00:53.71" />
                    <SPLIT distance="100" swimtime="00:01:13.15" />
                    <SPLIT distance="125" swimtime="00:01:32.82" />
                    <SPLIT distance="150" swimtime="00:01:53.74" />
                    <SPLIT distance="175" swimtime="00:02:15.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="315" reactiontime="+89" swimtime="00:01:09.08" resultid="5341" lane="8" heatid="6838" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.75" />
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                    <SPLIT distance="75" swimtime="00:00:51.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="277" reactiontime="+93" swimtime="00:00:35.22" resultid="5345" lane="1" heatid="7285" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="307" reactiontime="+99" swimtime="00:00:31.52" resultid="5346" lane="4" heatid="7340" entrytime="00:00:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1946-01-01" firstname="Janusz" gender="M" lastname="Woch" nation="POL" athleteid="5347">
              <RESULTS>
                <RESULT eventid="1411" points="178" reactiontime="+86" swimtime="00:03:46.29" resultid="5351" lane="7" heatid="7005" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.41" />
                    <SPLIT distance="50" swimtime="00:00:49.26" />
                    <SPLIT distance="75" swimtime="00:01:17.31" />
                    <SPLIT distance="100" swimtime="00:01:47.65" />
                    <SPLIT distance="125" swimtime="00:02:17.79" />
                    <SPLIT distance="150" swimtime="00:02:47.35" />
                    <SPLIT distance="175" swimtime="00:03:17.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="223" reactiontime="+79" swimtime="00:01:37.13" resultid="5353" heatid="7305" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.10" />
                    <SPLIT distance="50" swimtime="00:00:45.58" />
                    <SPLIT distance="75" swimtime="00:01:11.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="144" reactiontime="+83" swimtime="00:03:37.44" resultid="5352" lane="1" heatid="7073" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.88" />
                    <SPLIT distance="50" swimtime="00:00:45.57" />
                    <SPLIT distance="75" swimtime="00:01:15.57" />
                    <SPLIT distance="100" swimtime="00:01:43.95" />
                    <SPLIT distance="125" swimtime="00:02:13.50" />
                    <SPLIT distance="150" swimtime="00:02:42.44" />
                    <SPLIT distance="175" swimtime="00:03:12.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="159" reactiontime="+81" swimtime="00:03:29.94" resultid="5350" lane="8" heatid="6883" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.14" />
                    <SPLIT distance="50" swimtime="00:00:47.63" />
                    <SPLIT distance="75" swimtime="00:01:13.83" />
                    <SPLIT distance="100" swimtime="00:01:41.60" />
                    <SPLIT distance="125" swimtime="00:02:09.39" />
                    <SPLIT distance="150" swimtime="00:02:36.76" />
                    <SPLIT distance="175" swimtime="00:03:04.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="281" reactiontime="+75" swimtime="00:00:41.49" resultid="5349" lane="5" heatid="6858" entrytime="00:00:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="167" reactiontime="+87" swimtime="00:01:35.32" resultid="5354" lane="6" heatid="7321" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.47" />
                    <SPLIT distance="50" swimtime="00:00:46.37" />
                    <SPLIT distance="75" swimtime="00:01:10.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="189" reactiontime="+93" swimtime="00:01:29.11" resultid="5348" heatid="6733" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.85" />
                    <SPLIT distance="50" swimtime="00:00:41.78" />
                    <SPLIT distance="75" swimtime="00:01:07.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-01" firstname="Jacek" gender="M" lastname="Beszterda" nation="POL" athleteid="5355">
              <RESULTS>
                <RESULT eventid="1075" points="242" swimtime="00:12:15.72" resultid="5356" heatid="6720" entrytime="00:12:10.00" />
                <RESULT eventid="1564" points="232" reactiontime="+88" swimtime="00:02:47.55" resultid="5359" lane="8" heatid="7059" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.18" />
                    <SPLIT distance="50" swimtime="00:00:38.26" />
                    <SPLIT distance="75" swimtime="00:00:58.95" />
                    <SPLIT distance="100" swimtime="00:01:20.28" />
                    <SPLIT distance="125" swimtime="00:01:42.05" />
                    <SPLIT distance="150" swimtime="00:02:04.47" />
                    <SPLIT distance="175" swimtime="00:02:26.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="227" reactiontime="+77" swimtime="00:01:17.07" resultid="5357" lane="8" heatid="6835" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.23" />
                    <SPLIT distance="50" swimtime="00:00:36.58" />
                    <SPLIT distance="75" swimtime="00:00:56.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="226" reactiontime="+88" swimtime="00:00:34.92" resultid="5361" lane="6" heatid="7339" entrytime="00:00:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1645" points="123" reactiontime="+88" swimtime="00:00:46.08" resultid="5360" lane="4" heatid="7282" entrytime="00:00:42.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.38" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="04" eventid="1375" reactiontime="+41" status="DSQ" swimtime="00:05:55.80" resultid="5358" lane="7" heatid="6904" entrytime="00:05:52.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.48" />
                    <SPLIT distance="50" swimtime="00:00:37.43" />
                    <SPLIT distance="75" swimtime="00:00:59.30" />
                    <SPLIT distance="100" swimtime="00:01:21.21" />
                    <SPLIT distance="125" swimtime="00:01:44.13" />
                    <SPLIT distance="150" swimtime="00:02:07.00" />
                    <SPLIT distance="175" swimtime="00:02:30.62" />
                    <SPLIT distance="200" swimtime="00:02:53.98" />
                    <SPLIT distance="225" swimtime="00:03:16.96" />
                    <SPLIT distance="250" swimtime="00:03:40.11" />
                    <SPLIT distance="275" swimtime="00:04:03.24" />
                    <SPLIT distance="300" swimtime="00:04:26.33" />
                    <SPLIT distance="325" swimtime="00:04:49.16" />
                    <SPLIT distance="350" swimtime="00:05:11.52" />
                    <SPLIT distance="375" swimtime="00:05:34.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-01" firstname="Piotr" gender="M" lastname="Monczak" nation="POL" athleteid="5362">
              <RESULTS>
                <RESULT eventid="1798" points="433" reactiontime="+70" swimtime="00:05:22.10" resultid="5369" lane="2" heatid="7364" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.80" />
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                    <SPLIT distance="75" swimtime="00:00:52.18" />
                    <SPLIT distance="100" swimtime="00:01:11.93" />
                    <SPLIT distance="125" swimtime="00:01:33.13" />
                    <SPLIT distance="150" swimtime="00:01:53.78" />
                    <SPLIT distance="175" swimtime="00:02:14.29" />
                    <SPLIT distance="200" swimtime="00:02:35.40" />
                    <SPLIT distance="225" swimtime="00:02:58.82" />
                    <SPLIT distance="250" swimtime="00:03:22.31" />
                    <SPLIT distance="275" swimtime="00:03:46.43" />
                    <SPLIT distance="300" swimtime="00:04:10.13" />
                    <SPLIT distance="325" swimtime="00:04:28.77" />
                    <SPLIT distance="350" swimtime="00:04:46.66" />
                    <SPLIT distance="375" swimtime="00:05:04.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="538" reactiontime="+70" swimtime="00:00:26.15" resultid="5368" lane="2" heatid="7352" entrytime="00:00:26.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" points="464" reactiontime="+71" swimtime="00:04:44.12" resultid="5365" lane="4" heatid="6908" entrytime="00:04:47.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.77" />
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                    <SPLIT distance="75" swimtime="00:00:49.78" />
                    <SPLIT distance="100" swimtime="00:01:07.43" />
                    <SPLIT distance="125" swimtime="00:01:25.48" />
                    <SPLIT distance="150" swimtime="00:01:43.99" />
                    <SPLIT distance="175" swimtime="00:02:02.30" />
                    <SPLIT distance="200" swimtime="00:02:20.78" />
                    <SPLIT distance="225" swimtime="00:02:38.51" />
                    <SPLIT distance="250" swimtime="00:02:56.81" />
                    <SPLIT distance="275" swimtime="00:03:15.08" />
                    <SPLIT distance="300" swimtime="00:03:33.60" />
                    <SPLIT distance="325" swimtime="00:03:51.52" />
                    <SPLIT distance="350" swimtime="00:04:09.75" />
                    <SPLIT distance="375" swimtime="00:04:26.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="411" reactiontime="+74" swimtime="00:02:33.56" resultid="5367" heatid="7080" entrytime="00:02:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.76" />
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                    <SPLIT distance="75" swimtime="00:00:52.98" />
                    <SPLIT distance="100" swimtime="00:01:12.72" />
                    <SPLIT distance="125" swimtime="00:01:35.09" />
                    <SPLIT distance="150" swimtime="00:01:58.36" />
                    <SPLIT distance="175" swimtime="00:02:16.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="466" reactiontime="+75" swimtime="00:02:12.75" resultid="5366" lane="4" heatid="7065" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.25" />
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                    <SPLIT distance="75" swimtime="00:00:47.80" />
                    <SPLIT distance="100" swimtime="00:01:04.96" />
                    <SPLIT distance="125" swimtime="00:01:21.81" />
                    <SPLIT distance="150" swimtime="00:01:39.20" />
                    <SPLIT distance="175" swimtime="00:01:56.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="443" reactiontime="+72" swimtime="00:01:07.07" resultid="5363" heatid="6744" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.91" />
                    <SPLIT distance="50" swimtime="00:00:32.03" />
                    <SPLIT distance="75" swimtime="00:00:51.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="545" reactiontime="+72" swimtime="00:00:57.57" resultid="5364" lane="7" heatid="6845" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.44" />
                    <SPLIT distance="50" swimtime="00:00:28.05" />
                    <SPLIT distance="75" swimtime="00:00:42.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-01" firstname="Sabina" gender="F" lastname="Rogala-Łukaszewicz" nation="POL" athleteid="5370">
              <RESULTS>
                <RESULT eventid="1747" points="430" reactiontime="+69" swimtime="00:00:31.74" resultid="5376" lane="1" heatid="7334" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="413" reactiontime="+84" swimtime="00:01:10.96" resultid="5372" lane="4" heatid="6827" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.09" />
                    <SPLIT distance="50" swimtime="00:00:33.60" />
                    <SPLIT distance="75" swimtime="00:00:52.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1679" points="333" reactiontime="+83" swimtime="00:01:33.83" resultid="5375" lane="1" heatid="7299" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.62" />
                    <SPLIT distance="50" swimtime="00:00:43.17" />
                    <SPLIT distance="75" swimtime="00:01:08.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="241" reactiontime="+89" swimtime="00:06:27.67" resultid="5373" lane="1" heatid="6896" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.88" />
                    <SPLIT distance="50" swimtime="00:00:42.27" />
                    <SPLIT distance="75" swimtime="00:01:05.61" />
                    <SPLIT distance="100" swimtime="00:01:29.28" />
                    <SPLIT distance="125" swimtime="00:01:53.52" />
                    <SPLIT distance="150" swimtime="00:02:17.64" />
                    <SPLIT distance="175" swimtime="00:02:42.55" />
                    <SPLIT distance="200" swimtime="00:03:07.14" />
                    <SPLIT distance="225" swimtime="00:03:31.61" />
                    <SPLIT distance="250" swimtime="00:03:56.56" />
                    <SPLIT distance="275" swimtime="00:04:21.82" />
                    <SPLIT distance="300" swimtime="00:04:47.27" />
                    <SPLIT distance="325" swimtime="00:05:13.48" />
                    <SPLIT distance="350" swimtime="00:05:38.88" />
                    <SPLIT distance="375" swimtime="00:06:04.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="313" reactiontime="+75" swimtime="00:01:26.53" resultid="5371" lane="8" heatid="6727" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.56" />
                    <SPLIT distance="50" swimtime="00:00:41.28" />
                    <SPLIT distance="75" swimtime="00:01:07.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1547" status="DNS" swimtime="00:00:00.00" resultid="5374" lane="5" heatid="7051" entrytime="00:02:52.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1955-01-01" firstname="Paweł" gender="M" lastname="Łukaszewicz" nation="POL" athleteid="5377">
              <RESULTS>
                <RESULT eventid="1462" points="225" reactiontime="+93" swimtime="00:01:22.79" resultid="5381" lane="5" heatid="7018" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.63" />
                    <SPLIT distance="50" swimtime="00:00:36.07" />
                    <SPLIT distance="75" swimtime="00:00:58.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="252" reactiontime="+101" swimtime="00:01:23.08" resultid="5383" lane="6" heatid="7322" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.11" />
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                    <SPLIT distance="75" swimtime="00:01:01.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="255" reactiontime="+112" swimtime="00:02:59.64" resultid="5380" lane="1" heatid="6884" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.76" />
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                    <SPLIT distance="75" swimtime="00:01:03.86" />
                    <SPLIT distance="100" swimtime="00:01:26.89" />
                    <SPLIT distance="125" swimtime="00:01:50.59" />
                    <SPLIT distance="150" swimtime="00:02:14.32" />
                    <SPLIT distance="175" swimtime="00:02:37.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="230" swimtime="00:12:28.28" resultid="5378" lane="5" heatid="6718" entrytime="00:13:10.00" />
                <RESULT eventid="1205" points="305" reactiontime="+91" swimtime="00:01:09.84" resultid="5379" lane="2" heatid="6836" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.60" />
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                    <SPLIT distance="75" swimtime="00:00:51.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="5382" lane="1" heatid="7059" entrytime="00:02:41.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1967-01-01" firstname="Marek" gender="M" lastname="Nowak" nation="POL" athleteid="5384">
              <RESULTS>
                <RESULT eventid="1239" points="424" reactiontime="+74" swimtime="00:00:36.17" resultid="5385" lane="8" heatid="6864" entrytime="00:00:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" points="383" reactiontime="+74" swimtime="00:01:21.10" resultid="5387" lane="2" heatid="7309" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.29" />
                    <SPLIT distance="50" swimtime="00:00:37.63" />
                    <SPLIT distance="75" swimtime="00:00:58.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="355" reactiontime="+74" swimtime="00:02:59.92" resultid="5386" lane="7" heatid="7010" entrytime="00:03:01.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.49" />
                    <SPLIT distance="50" swimtime="00:00:40.68" />
                    <SPLIT distance="75" swimtime="00:01:03.54" />
                    <SPLIT distance="100" swimtime="00:01:26.75" />
                    <SPLIT distance="125" swimtime="00:01:50.05" />
                    <SPLIT distance="150" swimtime="00:02:13.87" />
                    <SPLIT distance="175" swimtime="00:02:37.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="5388" lane="5" heatid="7345" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-01" firstname="Paulina" gender="F" lastname="Dratwa" nation="POL" athleteid="5389">
              <RESULTS>
                <RESULT eventid="1222" status="DNS" swimtime="00:00:00.00" resultid="5390" lane="2" heatid="6853" entrytime="00:00:38.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1961-01-01" firstname="Wojciech" gender="M" lastname="Dmytrów" nation="POL" athleteid="5391">
              <RESULTS>
                <RESULT eventid="1696" points="396" reactiontime="+78" swimtime="00:01:20.21" resultid="5395" lane="5" heatid="7307" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.84" />
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                    <SPLIT distance="75" swimtime="00:00:58.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1411" points="356" reactiontime="+72" swimtime="00:02:59.82" resultid="5393" lane="2" heatid="7008" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.62" />
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                    <SPLIT distance="75" swimtime="00:01:01.26" />
                    <SPLIT distance="100" swimtime="00:01:24.14" />
                    <SPLIT distance="125" swimtime="00:01:47.37" />
                    <SPLIT distance="150" swimtime="00:02:11.49" />
                    <SPLIT distance="175" swimtime="00:02:35.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="429" reactiontime="+73" swimtime="00:00:36.02" resultid="5392" lane="3" heatid="6861" entrytime="00:00:37.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1598" points="240" reactiontime="+82" swimtime="00:03:03.80" resultid="5394" lane="8" heatid="7074" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.32" />
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                    <SPLIT distance="75" swimtime="00:01:05.58" />
                    <SPLIT distance="100" swimtime="00:01:31.12" />
                    <SPLIT distance="125" swimtime="00:01:54.52" />
                    <SPLIT distance="150" swimtime="00:02:19.22" />
                    <SPLIT distance="175" swimtime="00:02:42.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1960-01-01" firstname="Maciej" gender="M" lastname="Beszterda" nation="POL" athleteid="5396">
              <RESULTS>
                <RESULT eventid="1564" points="157" reactiontime="+109" swimtime="00:03:10.74" resultid="5399" lane="4" heatid="7056" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.65" />
                    <SPLIT distance="50" swimtime="00:00:41.86" />
                    <SPLIT distance="75" swimtime="00:01:05.28" />
                    <SPLIT distance="100" swimtime="00:01:29.62" />
                    <SPLIT distance="125" swimtime="00:01:54.58" />
                    <SPLIT distance="150" swimtime="00:02:20.79" />
                    <SPLIT distance="175" swimtime="00:02:46.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1307" points="126" reactiontime="+96" swimtime="00:03:46.71" resultid="5398" lane="1" heatid="6882" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.32" />
                    <SPLIT distance="50" swimtime="00:00:55.24" />
                    <SPLIT distance="75" swimtime="00:01:23.81" />
                    <SPLIT distance="100" swimtime="00:01:52.60" />
                    <SPLIT distance="125" swimtime="00:02:21.90" />
                    <SPLIT distance="150" swimtime="00:02:50.37" />
                    <SPLIT distance="175" swimtime="00:03:19.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" points="118" reactiontime="+127" swimtime="00:01:46.94" resultid="5400" lane="8" heatid="7320" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.74" />
                    <SPLIT distance="50" swimtime="00:00:53.33" />
                    <SPLIT distance="75" swimtime="00:01:21.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="5397" lane="6" heatid="6833" entrytime="00:01:20.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-01" firstname="Marek" gender="M" lastname="Libuda" nation="POL" athleteid="5401">
              <RESULTS>
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="5402" lane="5" heatid="7058" entrytime="00:02:45.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1965-01-01" firstname="Cezary" gender="M" lastname="Bąk" nation="POL" athleteid="5403">
              <RESULTS>
                <RESULT eventid="1496" points="151" reactiontime="+101" swimtime="00:00:45.88" resultid="5404" lane="8" heatid="7035" entrytime="00:00:48.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1730" status="DNS" swimtime="00:00:00.00" resultid="5405" lane="6" heatid="7320" entrytime="00:01:47.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariusz" gender="M" lastname="Rogowski" nation="POL" athleteid="5406">
              <RESULTS>
                <RESULT eventid="1530" points="30" swimtime="00:01:07.85" resultid="5407" lane="6" heatid="7046">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:31.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eugeniusz" gender="M" lastname="Gładyszak" nation="POL" athleteid="5408">
              <RESULTS>
                <RESULT eventid="1530" points="24" swimtime="00:01:13.50" resultid="5409" lane="8" heatid="7047">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:33.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edward" gender="M" lastname="Tomaszewski" nation="POL" athleteid="5410">
              <RESULTS>
                <RESULT eventid="1530" status="DNS" swimtime="00:00:00.00" resultid="5411" lane="1" heatid="7047" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Korneliusz" gender="M" lastname="Toliński" nation="POL" athleteid="5412">
              <RESULTS>
                <RESULT eventid="1530" status="DNS" swimtime="00:00:00.00" resultid="5413" lane="7" heatid="7046" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcin" gender="M" lastname="Straburzyński" nation="POL" athleteid="5414">
              <RESULTS>
                <RESULT eventid="1530" status="DNS" swimtime="00:00:00.00" resultid="5415" lane="7" heatid="7047" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateusz" gender="M" lastname="Suwriło" nation="POL" athleteid="5416">
              <RESULTS>
                <RESULT eventid="1530" status="DNS" swimtime="00:00:00.00" resultid="5417" lane="3" heatid="7046" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krzysztof" gender="M" lastname="Kołaczkowski" nation="POL" athleteid="5418">
              <RESULTS>
                <RESULT eventid="1530" points="125" swimtime="00:00:42.56" resultid="5419" lane="5" heatid="7046">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariola" gender="F" lastname="Dehr-Kołaczkowska" nation="POL" athleteid="5420">
              <RESULTS>
                <RESULT eventid="1513" points="72" swimtime="00:00:57.45" resultid="5421" lane="1" heatid="7044">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Małgorzata" gender="F" lastname="Kozłowska" nation="POL" athleteid="5422">
              <RESULTS>
                <RESULT eventid="1513" points="108" swimtime="00:00:50.18" resultid="5423" lane="6" heatid="7044">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="199" agemin="160" agetotalmax="-1" agetotalmin="-1" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1615" status="DNS" swimtime="00:00:00.00" resultid="5424" lane="4" heatid="7442" entrytime="00:02:08.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5384" number="1" />
                    <RELAYPOSITION athleteid="5389" number="2" />
                    <RELAYPOSITION athleteid="5370" number="3" />
                    <RELAYPOSITION athleteid="5362" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1815" status="DNS" swimtime="00:00:00.00" resultid="5425" lane="5" heatid="7503" entrytime="00:02:26.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="5384" number="1" />
                    <RELAYPOSITION athleteid="5389" number="2" />
                    <RELAYPOSITION athleteid="5362" number="3" />
                    <RELAYPOSITION athleteid="5370" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="UAPOZ" name="UAM Poznań">
          <ATHLETES>
            <ATHLETE birthdate="1987-01-01" firstname="Wojciech" gender="M" lastname="Górny" nation="POL" athleteid="5433">
              <RESULTS>
                <RESULT eventid="1696" status="DNS" swimtime="00:00:00.00" resultid="5442" lane="4" heatid="7301" />
                <RESULT eventid="1530" status="DNS" swimtime="00:00:00.00" resultid="5441" lane="3" heatid="7045" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Angelika" gender="F" lastname="Siemieniewska" athleteid="5435">
              <RESULTS>
                <RESULT eventid="1513" status="DNS" swimtime="00:00:00.00" resultid="5443" lane="8" heatid="7044" />
                <RESULT eventid="1222" status="DNS" swimtime="00:00:00.00" resultid="5444" lane="6" heatid="6847" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-01" firstname="Natalia" gender="F" lastname="Łukomska" athleteid="5436">
              <RESULTS>
                <RESULT eventid="1222" status="DNS" swimtime="00:00:00.00" resultid="5446" lane="2" heatid="6847" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Tymoteusz" gender="M" lastname="Leśniak" athleteid="5437">
              <RESULTS>
                <RESULT eventid="1530" points="185" reactiontime="+83" swimtime="00:00:37.33" resultid="5448" heatid="7047">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1696" status="DNS" swimtime="00:00:00.00" resultid="5447" lane="5" heatid="7301" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Norbert" gender="M" lastname="Kowalski" athleteid="5438">
              <RESULTS>
                <RESULT eventid="1239" status="DNS" swimtime="00:00:00.00" resultid="5450" heatid="6854" />
                <RESULT eventid="1530" points="184" reactiontime="+118" swimtime="00:00:37.38" resultid="5449" lane="1" heatid="7046">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1987-01-01" firstname="Adrian" gender="M" lastname="Gorczyca" athleteid="5439">
              <RESULTS>
                <RESULT eventid="1530" status="DNS" swimtime="00:00:00.00" resultid="5451" lane="4" heatid="7046" />
                <RESULT eventid="1496" status="DNS" swimtime="00:00:00.00" resultid="5452" lane="2" heatid="7032" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Michał" gender="M" lastname="Jurek" athleteid="5440">
              <RESULTS>
                <RESULT eventid="1530" points="160" reactiontime="+81" swimtime="00:00:39.16" resultid="5453" lane="5" heatid="7045">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1496" status="DNS" swimtime="00:00:00.00" resultid="5454" lane="6" heatid="7032" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ZIELO" name="Zielona Góra">
          <ATHLETES>
            <ATHLETE birthdate="1971-01-01" firstname="Sławomir" gender="M" lastname="Mąkowski" nation="POL" athleteid="5455">
              <RESULTS>
                <RESULT eventid="1496" points="318" reactiontime="+71" swimtime="00:00:35.84" resultid="5457" lane="5" heatid="7037" entrytime="00:00:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="370" reactiontime="+81" swimtime="00:00:29.62" resultid="5458" lane="4" heatid="7341" entrytime="00:00:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="RZESZO" name="Rzeszów">
          <ATHLETES>
            <ATHLETE birthdate="1957-01-01" firstname="Wiesław" gender="M" lastname="Ciekliński" nation="POL" athleteid="3893">
              <RESULTS>
                <RESULT eventid="1205" points="289" reactiontime="+80" swimtime="00:01:11.11" resultid="3895" lane="4" heatid="6837" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.49" />
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                    <SPLIT distance="75" swimtime="00:00:52.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1764" points="316" reactiontime="+86" swimtime="00:00:31.23" resultid="3899" lane="3" heatid="7343" entrytime="00:00:30.30">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="182" reactiontime="+86" swimtime="00:01:30.10" resultid="3894" lane="8" heatid="6734" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.18" />
                    <SPLIT distance="50" swimtime="00:00:40.71" />
                    <SPLIT distance="75" swimtime="00:01:10.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1375" status="DNS" swimtime="00:00:00.00" resultid="3896" lane="2" heatid="6903" entrytime="00:05:58.00" />
                <RESULT eventid="1564" status="DNS" swimtime="00:00:00.00" resultid="3897" lane="7" heatid="7059" entrytime="00:02:41.30" />
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="3898" heatid="7284" entrytime="00:00:37.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="GOWIE" name="Gorzów Wlkp.">
          <ATHLETES>
            <ATHLETE birthdate="1955-07-15" firstname="Marian" gender="M" lastname="Lasowy" nation="POL" athleteid="3341">
              <RESULTS>
                <RESULT eventid="1075" points="160" swimtime="00:14:03.72" resultid="3342" lane="1" heatid="6718" entrytime="00:13:59.00" entrycourse="SCM" />
                <RESULT eventid="1205" points="189" reactiontime="+113" swimtime="00:01:21.93" resultid="3343" heatid="6831" entrytime="00:01:43.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.25" />
                    <SPLIT distance="50" swimtime="00:00:37.52" />
                    <SPLIT distance="75" swimtime="00:00:59.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1530" status="DNS" swimtime="00:00:00.00" resultid="3344" lane="2" heatid="7047" entrytime="00:00:37.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="STSZC" name="Stargard Szczeciński">
          <ATHLETES>
            <ATHLETE birthdate="1983-01-01" firstname="Karol" gender="M" lastname="Grzywacz" nation="POL" athleteid="4755">
              <RESULTS>
                <RESULT eventid="1375" points="275" reactiontime="+79" swimtime="00:05:38.18" resultid="4758" lane="8" heatid="6906" entrytime="00:05:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.77" />
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                    <SPLIT distance="75" swimtime="00:00:53.13" />
                    <SPLIT distance="100" swimtime="00:01:13.64" />
                    <SPLIT distance="125" swimtime="00:01:34.87" />
                    <SPLIT distance="150" swimtime="00:01:56.47" />
                    <SPLIT distance="175" swimtime="00:02:18.55" />
                    <SPLIT distance="200" swimtime="00:02:40.70" />
                    <SPLIT distance="225" swimtime="00:03:02.82" />
                    <SPLIT distance="250" swimtime="00:03:25.02" />
                    <SPLIT distance="275" swimtime="00:03:47.19" />
                    <SPLIT distance="300" swimtime="00:04:09.32" />
                    <SPLIT distance="325" swimtime="00:04:31.63" />
                    <SPLIT distance="350" swimtime="00:04:53.70" />
                    <SPLIT distance="375" swimtime="00:05:16.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1564" points="276" reactiontime="+70" swimtime="00:02:37.97" resultid="4759" lane="8" heatid="7061" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.45" />
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                    <SPLIT distance="75" swimtime="00:00:52.10" />
                    <SPLIT distance="100" swimtime="00:01:12.09" />
                    <SPLIT distance="125" swimtime="00:01:33.90" />
                    <SPLIT distance="150" swimtime="00:01:55.25" />
                    <SPLIT distance="175" swimtime="00:02:17.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="315" reactiontime="+75" swimtime="00:01:09.09" resultid="4757" lane="8" heatid="6839" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.64" />
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                    <SPLIT distance="75" swimtime="00:00:49.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="252" reactiontime="+72" swimtime="00:01:20.88" resultid="4756" lane="4" heatid="6737" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.29" />
                    <SPLIT distance="50" swimtime="00:00:38.00" />
                    <SPLIT distance="75" swimtime="00:01:02.09" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="G 8" eventid="1598" status="DSQ" swimtime="00:00:00.00" resultid="4760" lane="6" heatid="7077" entrytime="00:02:55.00" />
                <RESULT eventid="1645" status="DNS" swimtime="00:00:00.00" resultid="4761" lane="5" heatid="7285" entrytime="00:00:35.00" />
                <RESULT eventid="1764" status="DNS" swimtime="00:00:00.00" resultid="4762" lane="2" heatid="7344" entrytime="00:00:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
